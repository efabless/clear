magic
tech sky130A
magscale 1 2
timestamp 1681041472
<< viali >>
rect 26433 24361 26467 24395
rect 27261 24361 27295 24395
rect 29745 24361 29779 24395
rect 41061 24361 41095 24395
rect 47869 24361 47903 24395
rect 25789 24293 25823 24327
rect 31217 24293 31251 24327
rect 38209 24293 38243 24327
rect 48513 24293 48547 24327
rect 2973 24225 3007 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10701 24225 10735 24259
rect 13277 24225 13311 24259
rect 15853 24225 15887 24259
rect 18429 24225 18463 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25145 24225 25179 24259
rect 29193 24225 29227 24259
rect 34253 24225 34287 24259
rect 35081 24225 35115 24259
rect 36553 24225 36587 24259
rect 36737 24225 36771 24259
rect 37565 24225 37599 24259
rect 40601 24225 40635 24259
rect 41429 24225 41463 24259
rect 45845 24225 45879 24259
rect 3433 24157 3467 24191
rect 3985 24157 4019 24191
rect 4629 24157 4663 24191
rect 6561 24157 6595 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 11161 24157 11195 24191
rect 11897 24157 11931 24191
rect 13737 24157 13771 24191
rect 14473 24157 14507 24191
rect 16313 24157 16347 24191
rect 18889 24157 18923 24191
rect 19625 24157 19659 24191
rect 21373 24157 21407 24191
rect 22017 24157 22051 24191
rect 23857 24157 23891 24191
rect 25973 24157 26007 24191
rect 27905 24157 27939 24191
rect 28549 24157 28583 24191
rect 29929 24157 29963 24191
rect 30389 24157 30423 24191
rect 31033 24157 31067 24191
rect 32505 24157 32539 24191
rect 33149 24157 33183 24191
rect 34069 24157 34103 24191
rect 38853 24157 38887 24191
rect 39497 24157 39531 24191
rect 42073 24157 42107 24191
rect 42625 24157 42659 24191
rect 43269 24157 43303 24191
rect 43913 24157 43947 24191
rect 44557 24157 44591 24191
rect 45201 24157 45235 24191
rect 47225 24157 47259 24191
rect 48697 24157 48731 24191
rect 49341 24157 49375 24191
rect 24961 24089 24995 24123
rect 26617 24089 26651 24123
rect 26801 24089 26835 24123
rect 27353 24089 27387 24123
rect 29009 24089 29043 24123
rect 33977 24089 34011 24123
rect 36461 24089 36495 24123
rect 37841 24089 37875 24123
rect 40417 24089 40451 24123
rect 47961 24089 47995 24123
rect 4169 24021 4203 24055
rect 6745 24021 6779 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 14289 24021 14323 24055
rect 17049 24021 17083 24055
rect 19441 24021 19475 24055
rect 24041 24021 24075 24055
rect 24593 24021 24627 24055
rect 25053 24021 25087 24055
rect 28089 24021 28123 24055
rect 28733 24021 28767 24055
rect 30573 24021 30607 24055
rect 31493 24021 31527 24055
rect 31677 24021 31711 24055
rect 31861 24021 31895 24055
rect 32321 24021 32355 24055
rect 32965 24021 32999 24055
rect 33609 24021 33643 24055
rect 35173 24021 35207 24055
rect 35265 24021 35299 24055
rect 35633 24021 35667 24055
rect 36093 24021 36127 24055
rect 37749 24021 37783 24055
rect 38669 24021 38703 24055
rect 39313 24021 39347 24055
rect 40049 24021 40083 24055
rect 40509 24021 40543 24055
rect 43729 24021 43763 24055
rect 44373 24021 44407 24055
rect 46121 24021 46155 24055
rect 46581 24021 46615 24055
rect 49157 24021 49191 24055
rect 2329 23817 2363 23851
rect 23305 23817 23339 23851
rect 28457 23817 28491 23851
rect 32321 23817 32355 23851
rect 32781 23817 32815 23851
rect 37473 23817 37507 23851
rect 37841 23817 37875 23851
rect 42165 23817 42199 23851
rect 47133 23817 47167 23851
rect 47685 23817 47719 23851
rect 49341 23817 49375 23851
rect 14289 23749 14323 23783
rect 20269 23749 20303 23783
rect 23673 23749 23707 23783
rect 26341 23749 26375 23783
rect 31493 23749 31527 23783
rect 37933 23749 37967 23783
rect 42625 23749 42659 23783
rect 49433 23749 49467 23783
rect 2145 23681 2179 23715
rect 4077 23681 4111 23715
rect 4721 23681 4755 23715
rect 6837 23681 6871 23715
rect 7297 23681 7331 23715
rect 9321 23681 9355 23715
rect 11161 23681 11195 23715
rect 12357 23681 12391 23715
rect 13093 23681 13127 23715
rect 16313 23681 16347 23715
rect 18245 23681 18279 23715
rect 21281 23705 21315 23739
rect 23765 23681 23799 23715
rect 27353 23681 27387 23715
rect 27813 23681 27847 23715
rect 28641 23681 28675 23715
rect 29101 23681 29135 23715
rect 29561 23681 29595 23715
rect 32689 23681 32723 23715
rect 36277 23681 36311 23715
rect 39221 23681 39255 23715
rect 40233 23681 40267 23715
rect 44833 23681 44867 23715
rect 45937 23681 45971 23715
rect 46673 23681 46707 23715
rect 48789 23681 48823 23715
rect 3709 23613 3743 23647
rect 5457 23613 5491 23647
rect 8861 23613 8895 23647
rect 10609 23613 10643 23647
rect 12633 23613 12667 23647
rect 15853 23613 15887 23647
rect 17877 23613 17911 23647
rect 20545 23613 20579 23647
rect 22569 23613 22603 23647
rect 22845 23613 22879 23647
rect 23857 23613 23891 23647
rect 26617 23613 26651 23647
rect 31769 23613 31803 23647
rect 32965 23613 32999 23647
rect 33609 23613 33643 23647
rect 35081 23613 35115 23647
rect 35357 23613 35391 23647
rect 36369 23613 36403 23647
rect 36461 23613 36495 23647
rect 38025 23613 38059 23647
rect 39313 23613 39347 23647
rect 39405 23613 39439 23647
rect 40693 23613 40727 23647
rect 40969 23613 41003 23647
rect 43085 23613 43119 23647
rect 47317 23613 47351 23647
rect 49065 23613 49099 23647
rect 7481 23545 7515 23579
rect 24501 23545 24535 23579
rect 27169 23545 27203 23579
rect 38853 23545 38887 23579
rect 40049 23545 40083 23579
rect 41797 23545 41831 23579
rect 46949 23545 46983 23579
rect 48145 23545 48179 23579
rect 6653 23477 6687 23511
rect 18797 23477 18831 23511
rect 21005 23477 21039 23511
rect 21465 23477 21499 23511
rect 24409 23477 24443 23511
rect 24869 23477 24903 23511
rect 27997 23477 28031 23511
rect 29285 23477 29319 23511
rect 30021 23477 30055 23511
rect 35909 23477 35943 23511
rect 36921 23477 36955 23511
rect 38577 23477 38611 23511
rect 41981 23477 42015 23511
rect 42441 23477 42475 23511
rect 45293 23477 45327 23511
rect 46489 23477 46523 23511
rect 47777 23477 47811 23511
rect 4721 23273 4755 23307
rect 14197 23273 14231 23307
rect 27905 23273 27939 23307
rect 29745 23273 29779 23307
rect 34161 23273 34195 23307
rect 38779 23273 38813 23307
rect 41061 23273 41095 23307
rect 44005 23273 44039 23307
rect 48881 23273 48915 23307
rect 49249 23273 49283 23307
rect 19625 23205 19659 23239
rect 24593 23205 24627 23239
rect 25237 23205 25271 23239
rect 29009 23205 29043 23239
rect 29377 23205 29411 23239
rect 33149 23205 33183 23239
rect 34437 23205 34471 23239
rect 46765 23205 46799 23239
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 10057 23137 10091 23171
rect 11253 23137 11287 23171
rect 13277 23137 13311 23171
rect 15761 23137 15795 23171
rect 21833 23137 21867 23171
rect 23949 23137 23983 23171
rect 25973 23137 26007 23171
rect 28457 23137 28491 23171
rect 29193 23137 29227 23171
rect 30205 23137 30239 23171
rect 30297 23137 30331 23171
rect 31033 23137 31067 23171
rect 35081 23137 35115 23171
rect 37289 23137 37323 23171
rect 39037 23137 39071 23171
rect 39497 23137 39531 23171
rect 40693 23137 40727 23171
rect 43545 23137 43579 23171
rect 45201 23137 45235 23171
rect 2973 23069 3007 23103
rect 4261 23069 4295 23103
rect 4905 23069 4939 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9321 23069 9355 23103
rect 11897 23069 11931 23103
rect 13737 23069 13771 23103
rect 14841 23069 14875 23103
rect 16681 23069 16715 23103
rect 18889 23069 18923 23103
rect 22109 23069 22143 23103
rect 23765 23069 23799 23103
rect 24777 23069 24811 23103
rect 25697 23069 25731 23103
rect 28365 23069 28399 23103
rect 31401 23069 31435 23103
rect 33885 23069 33919 23103
rect 34713 23069 34747 23103
rect 40417 23069 40451 23103
rect 44649 23069 44683 23103
rect 46949 23069 46983 23103
rect 47777 23069 47811 23103
rect 48237 23069 48271 23103
rect 1777 23001 1811 23035
rect 18613 23001 18647 23035
rect 19809 23001 19843 23035
rect 22569 23001 22603 23035
rect 22753 23001 22787 23035
rect 31677 23001 31711 23035
rect 35357 23001 35391 23035
rect 41521 23001 41555 23035
rect 43269 23001 43303 23035
rect 45385 23001 45419 23035
rect 46029 23001 46063 23035
rect 46213 23001 46247 23035
rect 4077 22933 4111 22967
rect 9229 22933 9263 22967
rect 14289 22933 14323 22967
rect 14657 22933 14691 22967
rect 17141 22933 17175 22967
rect 19257 22933 19291 22967
rect 20361 22933 20395 22967
rect 23305 22933 23339 22967
rect 23673 22933 23707 22967
rect 25329 22933 25363 22967
rect 27445 22933 27479 22967
rect 28273 22933 28307 22967
rect 30113 22933 30147 22967
rect 30757 22933 30791 22967
rect 33701 22933 33735 22967
rect 36829 22933 36863 22967
rect 39405 22933 39439 22967
rect 40049 22933 40083 22967
rect 40509 22933 40543 22967
rect 47593 22933 47627 22967
rect 49433 22933 49467 22967
rect 18613 22729 18647 22763
rect 19165 22729 19199 22763
rect 21189 22729 21223 22763
rect 32321 22729 32355 22763
rect 32689 22729 32723 22763
rect 35449 22729 35483 22763
rect 36093 22729 36127 22763
rect 37473 22729 37507 22763
rect 39497 22729 39531 22763
rect 39773 22729 39807 22763
rect 46213 22729 46247 22763
rect 47041 22729 47075 22763
rect 47685 22729 47719 22763
rect 48053 22729 48087 22763
rect 4813 22661 4847 22695
rect 7113 22661 7147 22695
rect 9965 22661 9999 22695
rect 12817 22661 12851 22695
rect 15117 22661 15151 22695
rect 24133 22661 24167 22695
rect 26341 22661 26375 22695
rect 38945 22661 38979 22695
rect 40417 22661 40451 22695
rect 43729 22661 43763 22695
rect 44373 22661 44407 22695
rect 2973 22593 3007 22627
rect 3985 22593 4019 22627
rect 6009 22593 6043 22627
rect 6653 22593 6687 22627
rect 7481 22593 7515 22627
rect 11161 22593 11195 22627
rect 11897 22593 11931 22627
rect 14013 22593 14047 22627
rect 16313 22593 16347 22627
rect 16865 22593 16899 22627
rect 19441 22593 19475 22627
rect 21649 22593 21683 22627
rect 22017 22593 22051 22627
rect 24409 22593 24443 22627
rect 26617 22593 26651 22627
rect 27169 22593 27203 22627
rect 29837 22593 29871 22627
rect 30665 22593 30699 22627
rect 30757 22593 30791 22627
rect 31677 22593 31711 22627
rect 32781 22593 32815 22627
rect 33701 22593 33735 22627
rect 36461 22593 36495 22627
rect 39221 22593 39255 22627
rect 40509 22593 40543 22627
rect 41429 22593 41463 22627
rect 42073 22593 42107 22627
rect 42625 22593 42659 22627
rect 45109 22593 45143 22627
rect 45753 22593 45787 22627
rect 46397 22593 46431 22627
rect 47225 22593 47259 22627
rect 47777 22593 47811 22627
rect 48605 22593 48639 22627
rect 49341 22593 49375 22627
rect 2513 22525 2547 22559
rect 7941 22525 7975 22559
rect 9321 22525 9355 22559
rect 17141 22525 17175 22559
rect 18889 22525 18923 22559
rect 19717 22525 19751 22559
rect 22293 22525 22327 22559
rect 28089 22525 28123 22559
rect 29561 22525 29595 22559
rect 30849 22525 30883 22559
rect 32873 22525 32907 22559
rect 33977 22525 34011 22559
rect 36553 22525 36587 22559
rect 36737 22525 36771 22559
rect 40601 22525 40635 22559
rect 42901 22525 42935 22559
rect 4169 22457 4203 22491
rect 6837 22457 6871 22491
rect 11713 22457 11747 22491
rect 24501 22457 24535 22491
rect 27353 22457 27387 22491
rect 44925 22457 44959 22491
rect 45569 22457 45603 22491
rect 9505 22389 9539 22423
rect 12357 22389 12391 22423
rect 14381 22389 14415 22423
rect 14565 22389 14599 22423
rect 23765 22389 23799 22423
rect 24869 22389 24903 22423
rect 27721 22389 27755 22423
rect 30297 22389 30331 22423
rect 31493 22389 31527 22423
rect 33425 22389 33459 22423
rect 35817 22389 35851 22423
rect 40049 22389 40083 22423
rect 41245 22389 41279 22423
rect 41889 22389 41923 22423
rect 44281 22389 44315 22423
rect 48421 22389 48455 22423
rect 49157 22389 49191 22423
rect 12357 22185 12391 22219
rect 15209 22185 15243 22219
rect 24593 22185 24627 22219
rect 27169 22185 27203 22219
rect 30297 22185 30331 22219
rect 40233 22185 40267 22219
rect 41429 22185 41463 22219
rect 43177 22185 43211 22219
rect 45201 22185 45235 22219
rect 45385 22185 45419 22219
rect 45661 22185 45695 22219
rect 47041 22185 47075 22219
rect 47593 22185 47627 22219
rect 25973 22117 26007 22151
rect 28365 22117 28399 22151
rect 39405 22117 39439 22151
rect 6009 22049 6043 22083
rect 9781 22049 9815 22083
rect 11897 22049 11931 22083
rect 13645 22049 13679 22083
rect 14473 22049 14507 22083
rect 17601 22049 17635 22083
rect 22017 22049 22051 22083
rect 23213 22049 23247 22083
rect 25053 22049 25087 22083
rect 25145 22049 25179 22083
rect 26617 22049 26651 22083
rect 27721 22049 27755 22083
rect 28917 22049 28951 22083
rect 33701 22049 33735 22083
rect 34437 22049 34471 22083
rect 35081 22049 35115 22083
rect 36185 22049 36219 22083
rect 38853 22049 38887 22083
rect 39129 22049 39163 22083
rect 40693 22049 40727 22083
rect 40877 22049 40911 22083
rect 41981 22049 42015 22083
rect 45017 22049 45051 22083
rect 48053 22049 48087 22083
rect 2973 21981 3007 22015
rect 5365 21981 5399 22015
rect 7205 21981 7239 22015
rect 7849 21981 7883 22015
rect 8585 21981 8619 22015
rect 9137 21981 9171 22015
rect 11621 21981 11655 22015
rect 12541 21981 12575 22015
rect 16957 21981 16991 22015
rect 18797 21981 18831 22015
rect 19441 21981 19475 22015
rect 21189 21981 21223 22015
rect 24041 21981 24075 22015
rect 26433 21981 26467 22015
rect 27629 21981 27663 22015
rect 28733 21981 28767 22015
rect 29929 21981 29963 22015
rect 30849 21981 30883 22015
rect 34069 21981 34103 22015
rect 36461 21981 36495 22015
rect 42809 21981 42843 22015
rect 43821 21981 43855 22015
rect 44097 21981 44131 22015
rect 46029 21981 46063 22015
rect 46581 21981 46615 22015
rect 47225 21981 47259 22015
rect 47685 21981 47719 22015
rect 1777 21913 1811 21947
rect 4169 21913 4203 21947
rect 7665 21913 7699 21947
rect 14657 21913 14691 21947
rect 16681 21913 16715 21947
rect 20361 21913 20395 21947
rect 21833 21913 21867 21947
rect 21925 21913 21959 21947
rect 23029 21913 23063 21947
rect 25697 21913 25731 21947
rect 27537 21913 27571 21947
rect 28825 21913 28859 21947
rect 31125 21913 31159 21947
rect 33517 21913 33551 21947
rect 35173 21913 35207 21947
rect 41797 21913 41831 21947
rect 48237 21913 48271 21947
rect 49249 21913 49283 21947
rect 8401 21845 8435 21879
rect 13001 21845 13035 21879
rect 13369 21845 13403 21879
rect 13461 21845 13495 21879
rect 14105 21845 14139 21879
rect 21465 21845 21499 21879
rect 22661 21845 22695 21879
rect 23121 21845 23155 21879
rect 23857 21845 23891 21879
rect 24961 21845 24995 21879
rect 26341 21845 26375 21879
rect 29745 21845 29779 21879
rect 30389 21845 30423 21879
rect 32597 21845 32631 21879
rect 33057 21845 33091 21879
rect 33425 21845 33459 21879
rect 34345 21845 34379 21879
rect 35265 21845 35299 21879
rect 35633 21845 35667 21879
rect 36369 21845 36403 21879
rect 36829 21845 36863 21879
rect 37381 21845 37415 21879
rect 39589 21845 39623 21879
rect 39865 21845 39899 21879
rect 40601 21845 40635 21879
rect 41889 21845 41923 21879
rect 42625 21845 42659 21879
rect 43361 21845 43395 21879
rect 43545 21845 43579 21879
rect 46397 21845 46431 21879
rect 48789 21845 48823 21879
rect 49157 21845 49191 21879
rect 10517 21641 10551 21675
rect 13921 21641 13955 21675
rect 16865 21641 16899 21675
rect 17417 21641 17451 21675
rect 17877 21641 17911 21675
rect 24777 21641 24811 21675
rect 25973 21641 26007 21675
rect 27169 21641 27203 21675
rect 27629 21641 27663 21675
rect 28365 21641 28399 21675
rect 28825 21641 28859 21675
rect 32781 21641 32815 21675
rect 33609 21641 33643 21675
rect 34713 21641 34747 21675
rect 34805 21641 34839 21675
rect 36921 21641 36955 21675
rect 40049 21641 40083 21675
rect 40233 21641 40267 21675
rect 40417 21641 40451 21675
rect 40693 21641 40727 21675
rect 42533 21641 42567 21675
rect 43729 21641 43763 21675
rect 44281 21641 44315 21675
rect 44465 21641 44499 21675
rect 47041 21641 47075 21675
rect 47869 21641 47903 21675
rect 3617 21573 3651 21607
rect 11713 21573 11747 21607
rect 13093 21573 13127 21607
rect 14841 21573 14875 21607
rect 21189 21573 21223 21607
rect 27537 21573 27571 21607
rect 31217 21573 31251 21607
rect 36093 21573 36127 21607
rect 40969 21573 41003 21607
rect 46765 21573 46799 21607
rect 2973 21505 3007 21539
rect 4629 21505 4663 21539
rect 5733 21505 5767 21539
rect 6653 21505 6687 21539
rect 8493 21505 8527 21539
rect 10701 21505 10735 21539
rect 12357 21505 12391 21539
rect 13277 21505 13311 21539
rect 14105 21505 14139 21539
rect 17785 21505 17819 21539
rect 21373 21505 21407 21539
rect 25145 21505 25179 21539
rect 25789 21505 25823 21539
rect 26617 21505 26651 21539
rect 28733 21505 28767 21539
rect 29929 21505 29963 21539
rect 30021 21505 30055 21539
rect 31125 21505 31159 21539
rect 33517 21505 33551 21539
rect 36737 21505 36771 21539
rect 37289 21505 37323 21539
rect 43453 21505 43487 21539
rect 43913 21505 43947 21539
rect 47225 21505 47259 21539
rect 47777 21505 47811 21539
rect 48605 21505 48639 21539
rect 49341 21505 49375 21539
rect 1777 21437 1811 21471
rect 7021 21437 7055 21471
rect 8861 21437 8895 21471
rect 12817 21437 12851 21471
rect 14565 21437 14599 21471
rect 18061 21437 18095 21471
rect 18613 21437 18647 21471
rect 18889 21437 18923 21471
rect 22477 21437 22511 21471
rect 22753 21437 22787 21471
rect 25237 21437 25271 21471
rect 25421 21437 25455 21471
rect 27721 21437 27755 21471
rect 28917 21437 28951 21471
rect 30113 21437 30147 21471
rect 31401 21437 31435 21471
rect 33333 21437 33367 21471
rect 34621 21437 34655 21471
rect 36185 21437 36219 21471
rect 36277 21437 36311 21471
rect 38025 21437 38059 21471
rect 38301 21437 38335 21471
rect 41245 21437 41279 21471
rect 41521 21437 41555 21471
rect 44097 21437 44131 21471
rect 5917 21369 5951 21403
rect 11161 21369 11195 21403
rect 11897 21369 11931 21403
rect 16773 21369 16807 21403
rect 17141 21369 17175 21403
rect 20361 21369 20395 21403
rect 26433 21369 26467 21403
rect 42717 21369 42751 21403
rect 48421 21369 48455 21403
rect 11345 21301 11379 21335
rect 12265 21301 12299 21335
rect 16313 21301 16347 21335
rect 20729 21301 20763 21335
rect 20913 21301 20947 21335
rect 21925 21301 21959 21335
rect 22109 21301 22143 21335
rect 24225 21301 24259 21335
rect 29561 21301 29595 21335
rect 30757 21301 30791 21335
rect 31769 21301 31803 21335
rect 33977 21301 34011 21335
rect 35173 21301 35207 21335
rect 35725 21301 35759 21335
rect 37565 21301 37599 21335
rect 37657 21301 37691 21335
rect 39773 21301 39807 21335
rect 42809 21301 42843 21335
rect 43269 21301 43303 21335
rect 49157 21301 49191 21335
rect 7481 21097 7515 21131
rect 9229 21097 9263 21131
rect 12449 21097 12483 21131
rect 14289 21097 14323 21131
rect 17141 21097 17175 21131
rect 24041 21097 24075 21131
rect 26893 21097 26927 21131
rect 29745 21097 29779 21131
rect 30205 21097 30239 21131
rect 40049 21097 40083 21131
rect 42533 21097 42567 21131
rect 42901 21097 42935 21131
rect 47317 21097 47351 21131
rect 49157 21097 49191 21131
rect 12725 21029 12759 21063
rect 13553 21029 13587 21063
rect 19349 21029 19383 21063
rect 19993 21029 20027 21063
rect 21189 21029 21223 21063
rect 23397 21029 23431 21063
rect 25697 21029 25731 21063
rect 30389 21029 30423 21063
rect 34253 21029 34287 21063
rect 42625 21029 42659 21063
rect 48421 21029 48455 21063
rect 2513 20961 2547 20995
rect 4169 20961 4203 20995
rect 6009 20961 6043 20995
rect 10057 20961 10091 20995
rect 10701 20961 10735 20995
rect 20545 20961 20579 20995
rect 22661 20961 22695 20995
rect 24225 20961 24259 20995
rect 25145 20961 25179 20995
rect 25329 20961 25363 20995
rect 26249 20961 26283 20995
rect 27905 20961 27939 20995
rect 28549 20961 28583 20995
rect 31309 20961 31343 20995
rect 31493 20961 31527 20995
rect 32781 20961 32815 20995
rect 37105 20961 37139 20995
rect 39405 20961 39439 20995
rect 40509 20961 40543 20995
rect 40601 20961 40635 20995
rect 41797 20961 41831 20995
rect 2973 20893 3007 20927
rect 5365 20893 5399 20927
rect 7205 20893 7239 20927
rect 8033 20893 8067 20927
rect 8401 20893 8435 20927
rect 9413 20893 9447 20927
rect 11345 20893 11379 20927
rect 11989 20893 12023 20927
rect 13737 20893 13771 20927
rect 16037 20893 16071 20927
rect 18889 20893 18923 20927
rect 20361 20893 20395 20927
rect 22937 20893 22971 20927
rect 24593 20893 24627 20927
rect 27445 20893 27479 20927
rect 29929 20893 29963 20927
rect 32505 20893 32539 20927
rect 36645 20893 36679 20927
rect 47961 20893 47995 20927
rect 48605 20893 48639 20927
rect 49341 20893 49375 20927
rect 12909 20825 12943 20859
rect 15761 20825 15795 20859
rect 16681 20825 16715 20859
rect 18613 20825 18647 20859
rect 23581 20825 23615 20859
rect 36369 20825 36403 20859
rect 37289 20825 37323 20859
rect 39129 20825 39163 20859
rect 40417 20825 40451 20859
rect 41705 20825 41739 20859
rect 42349 20825 42383 20859
rect 47501 20825 47535 20859
rect 7849 20757 7883 20791
rect 11161 20757 11195 20791
rect 11897 20757 11931 20791
rect 19533 20757 19567 20791
rect 19625 20757 19659 20791
rect 20453 20757 20487 20791
rect 24777 20757 24811 20791
rect 26065 20757 26099 20791
rect 26157 20757 26191 20791
rect 26709 20757 26743 20791
rect 28641 20757 28675 20791
rect 28733 20757 28767 20791
rect 29101 20757 29135 20791
rect 30849 20757 30883 20791
rect 31217 20757 31251 20791
rect 31953 20757 31987 20791
rect 34897 20757 34931 20791
rect 36921 20757 36955 20791
rect 37657 20757 37691 20791
rect 41245 20757 41279 20791
rect 41613 20757 41647 20791
rect 47777 20757 47811 20791
rect 5457 20553 5491 20587
rect 9689 20553 9723 20587
rect 10333 20553 10367 20587
rect 13737 20553 13771 20587
rect 14105 20553 14139 20587
rect 14933 20553 14967 20587
rect 15577 20553 15611 20587
rect 15945 20553 15979 20587
rect 16037 20553 16071 20587
rect 18797 20553 18831 20587
rect 19717 20553 19751 20587
rect 35265 20553 35299 20587
rect 41153 20553 41187 20587
rect 48053 20553 48087 20587
rect 3617 20485 3651 20519
rect 12633 20485 12667 20519
rect 19073 20485 19107 20519
rect 21189 20485 21223 20519
rect 22385 20485 22419 20519
rect 29837 20485 29871 20519
rect 31033 20485 31067 20519
rect 31125 20485 31159 20519
rect 31769 20485 31803 20519
rect 33793 20485 33827 20519
rect 40233 20485 40267 20519
rect 41797 20485 41831 20519
rect 2973 20417 3007 20451
rect 4813 20417 4847 20451
rect 5273 20417 5307 20451
rect 6561 20417 6595 20451
rect 9229 20417 9263 20451
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 11713 20417 11747 20451
rect 11897 20417 11931 20451
rect 12449 20417 12483 20451
rect 14197 20417 14231 20451
rect 15117 20417 15151 20451
rect 17049 20417 17083 20451
rect 21465 20417 21499 20451
rect 23397 20417 23431 20451
rect 23857 20417 23891 20451
rect 26065 20417 26099 20451
rect 27261 20417 27295 20451
rect 29745 20417 29779 20451
rect 34897 20417 34931 20451
rect 35725 20417 35759 20451
rect 36461 20417 36495 20451
rect 36553 20417 36587 20451
rect 39497 20417 39531 20451
rect 40325 20417 40359 20451
rect 48605 20417 48639 20451
rect 49341 20417 49375 20451
rect 2513 20349 2547 20383
rect 7021 20349 7055 20383
rect 11161 20349 11195 20383
rect 14289 20349 14323 20383
rect 16221 20349 16255 20383
rect 17325 20349 17359 20383
rect 22477 20349 22511 20383
rect 22569 20349 22603 20383
rect 24133 20349 24167 20383
rect 27537 20349 27571 20383
rect 29009 20349 29043 20383
rect 29561 20349 29595 20383
rect 31217 20349 31251 20383
rect 32321 20349 32355 20383
rect 34069 20349 34103 20383
rect 34713 20349 34747 20383
rect 34805 20349 34839 20383
rect 36737 20349 36771 20383
rect 39221 20349 39255 20383
rect 40141 20349 40175 20383
rect 47961 20349 47995 20383
rect 23213 20281 23247 20315
rect 26617 20281 26651 20315
rect 31953 20281 31987 20315
rect 35541 20281 35575 20315
rect 36093 20281 36127 20315
rect 41705 20281 41739 20315
rect 49157 20281 49191 20315
rect 9045 20213 9079 20247
rect 13001 20213 13035 20247
rect 13185 20213 13219 20247
rect 13461 20213 13495 20247
rect 16773 20213 16807 20247
rect 19349 20213 19383 20247
rect 22017 20213 22051 20247
rect 25605 20213 25639 20247
rect 26249 20213 26283 20247
rect 30205 20213 30239 20247
rect 30665 20213 30699 20247
rect 37381 20213 37415 20247
rect 37749 20213 37783 20247
rect 40693 20213 40727 20247
rect 48421 20213 48455 20247
rect 11345 20009 11379 20043
rect 14473 20009 14507 20043
rect 16865 20009 16899 20043
rect 18153 20009 18187 20043
rect 25605 20009 25639 20043
rect 26801 20009 26835 20043
rect 29009 20009 29043 20043
rect 31677 20009 31711 20043
rect 39037 20009 39071 20043
rect 41245 20009 41279 20043
rect 48789 20009 48823 20043
rect 9965 19941 9999 19975
rect 14933 19941 14967 19975
rect 15669 19941 15703 19975
rect 19625 19941 19659 19975
rect 24041 19941 24075 19975
rect 29285 19941 29319 19975
rect 34161 19941 34195 19975
rect 4261 19873 4295 19907
rect 6009 19873 6043 19907
rect 11989 19873 12023 19907
rect 16313 19873 16347 19907
rect 17509 19873 17543 19907
rect 18797 19873 18831 19907
rect 19349 19873 19383 19907
rect 22293 19873 22327 19907
rect 23397 19873 23431 19907
rect 23581 19873 23615 19907
rect 24593 19873 24627 19907
rect 26249 19873 26283 19907
rect 27353 19873 27387 19907
rect 28549 19873 28583 19907
rect 30205 19873 30239 19907
rect 30297 19873 30331 19907
rect 31125 19873 31159 19907
rect 32689 19873 32723 19907
rect 33609 19873 33643 19907
rect 33701 19873 33735 19907
rect 35081 19873 35115 19907
rect 36737 19873 36771 19907
rect 38025 19873 38059 19907
rect 40141 19873 40175 19907
rect 40325 19873 40359 19907
rect 2973 19805 3007 19839
rect 5365 19805 5399 19839
rect 7205 19805 7239 19839
rect 7941 19805 7975 19839
rect 10149 19805 10183 19839
rect 10793 19805 10827 19839
rect 14289 19805 14323 19839
rect 15117 19805 15151 19839
rect 18521 19805 18555 19839
rect 20269 19805 20303 19839
rect 22753 19805 22787 19839
rect 23029 19805 23063 19839
rect 23673 19805 23707 19839
rect 32505 19805 32539 19839
rect 33793 19805 33827 19839
rect 35265 19805 35299 19839
rect 38117 19805 38151 19839
rect 38209 19805 38243 19839
rect 38853 19805 38887 19839
rect 40417 19805 40451 19839
rect 41061 19805 41095 19839
rect 1777 19737 1811 19771
rect 11437 19737 11471 19771
rect 12265 19737 12299 19771
rect 16037 19737 16071 19771
rect 19809 19737 19843 19771
rect 22017 19737 22051 19771
rect 25145 19737 25179 19771
rect 25973 19737 26007 19771
rect 28457 19737 28491 19771
rect 31217 19737 31251 19771
rect 32597 19737 32631 19771
rect 36461 19737 36495 19771
rect 48605 19737 48639 19771
rect 49249 19737 49283 19771
rect 7757 19669 7791 19703
rect 10609 19669 10643 19703
rect 13737 19669 13771 19703
rect 16129 19669 16163 19703
rect 17233 19669 17267 19703
rect 17325 19669 17359 19703
rect 18613 19669 18647 19703
rect 20545 19669 20579 19703
rect 22661 19669 22695 19703
rect 25329 19669 25363 19703
rect 26065 19669 26099 19703
rect 27169 19669 27203 19703
rect 27261 19669 27295 19703
rect 27997 19669 28031 19703
rect 28365 19669 28399 19703
rect 29745 19669 29779 19703
rect 30113 19669 30147 19703
rect 31309 19669 31343 19703
rect 32137 19669 32171 19703
rect 34437 19669 34471 19703
rect 35173 19669 35207 19703
rect 35633 19669 35667 19703
rect 36093 19669 36127 19703
rect 36553 19669 36587 19703
rect 37381 19669 37415 19703
rect 37565 19669 37599 19703
rect 38577 19669 38611 19703
rect 39589 19669 39623 19703
rect 40785 19669 40819 19703
rect 49157 19669 49191 19703
rect 10977 19465 11011 19499
rect 15393 19465 15427 19499
rect 16865 19465 16899 19499
rect 21189 19465 21223 19499
rect 26157 19465 26191 19499
rect 28457 19465 28491 19499
rect 32689 19465 32723 19499
rect 33057 19465 33091 19499
rect 33793 19465 33827 19499
rect 35081 19465 35115 19499
rect 35449 19465 35483 19499
rect 37289 19465 37323 19499
rect 37473 19465 37507 19499
rect 40141 19465 40175 19499
rect 40601 19465 40635 19499
rect 41337 19465 41371 19499
rect 3617 19397 3651 19431
rect 10517 19397 10551 19431
rect 26249 19397 26283 19431
rect 31493 19397 31527 19431
rect 36185 19397 36219 19431
rect 40509 19397 40543 19431
rect 1777 19329 1811 19363
rect 2973 19329 3007 19363
rect 4813 19329 4847 19363
rect 5457 19329 5491 19363
rect 11161 19329 11195 19363
rect 11713 19329 11747 19363
rect 12173 19329 12207 19363
rect 14473 19329 14507 19363
rect 15485 19329 15519 19363
rect 16221 19329 16255 19363
rect 17233 19329 17267 19363
rect 17325 19329 17359 19363
rect 18061 19329 18095 19363
rect 21097 19329 21131 19363
rect 22937 19329 22971 19363
rect 25237 19329 25271 19363
rect 27629 19329 27663 19363
rect 28825 19329 28859 19363
rect 29745 19329 29779 19363
rect 30757 19329 30791 19363
rect 32597 19329 32631 19363
rect 33885 19329 33919 19363
rect 36277 19329 36311 19363
rect 39681 19329 39715 19363
rect 48605 19329 48639 19363
rect 49249 19329 49283 19363
rect 5273 19261 5307 19295
rect 9873 19261 9907 19295
rect 11989 19261 12023 19295
rect 14197 19261 14231 19295
rect 15025 19261 15059 19295
rect 16037 19261 16071 19295
rect 17417 19261 17451 19295
rect 19809 19261 19843 19295
rect 20085 19261 20119 19295
rect 20453 19261 20487 19295
rect 21373 19261 21407 19295
rect 22201 19261 22235 19295
rect 24961 19261 24995 19295
rect 26433 19261 26467 19295
rect 27721 19261 27755 19295
rect 27905 19261 27939 19295
rect 28917 19261 28951 19295
rect 29009 19261 29043 19295
rect 32505 19261 32539 19295
rect 33701 19261 33735 19295
rect 34897 19261 34931 19295
rect 34989 19261 35023 19295
rect 36001 19261 36035 19295
rect 39405 19261 39439 19295
rect 40693 19261 40727 19295
rect 34253 19193 34287 19227
rect 49065 19193 49099 19227
rect 5825 19125 5859 19159
rect 12725 19125 12759 19159
rect 14841 19125 14875 19159
rect 20729 19125 20763 19159
rect 23489 19125 23523 19159
rect 25789 19125 25823 19159
rect 27261 19125 27295 19159
rect 30205 19125 30239 19159
rect 30389 19125 30423 19159
rect 36645 19125 36679 19159
rect 36921 19125 36955 19159
rect 37933 19125 37967 19159
rect 41153 19125 41187 19159
rect 48789 19125 48823 19159
rect 9229 18921 9263 18955
rect 11897 18921 11931 18955
rect 16037 18921 16071 18955
rect 16405 18921 16439 18955
rect 16957 18921 16991 18955
rect 18153 18921 18187 18955
rect 19901 18921 19935 18955
rect 21097 18921 21131 18955
rect 27537 18921 27571 18955
rect 31493 18921 31527 18955
rect 37381 18921 37415 18955
rect 42073 18921 42107 18955
rect 13645 18853 13679 18887
rect 28181 18853 28215 18887
rect 29009 18853 29043 18887
rect 30941 18853 30975 18887
rect 33425 18853 33459 18887
rect 34161 18853 34195 18887
rect 34529 18853 34563 18887
rect 38025 18853 38059 18887
rect 49157 18853 49191 18887
rect 4169 18785 4203 18819
rect 10977 18785 11011 18819
rect 13093 18785 13127 18819
rect 14289 18785 14323 18819
rect 17509 18785 17543 18819
rect 18613 18785 18647 18819
rect 18797 18785 18831 18819
rect 20453 18785 20487 18819
rect 21649 18785 21683 18819
rect 22293 18785 22327 18819
rect 25053 18785 25087 18819
rect 25237 18785 25271 18819
rect 25789 18785 25823 18819
rect 28089 18785 28123 18819
rect 29837 18785 29871 18819
rect 30021 18785 30055 18819
rect 32137 18785 32171 18819
rect 32781 18785 32815 18819
rect 32965 18785 32999 18819
rect 33885 18785 33919 18819
rect 35633 18785 35667 18819
rect 38577 18785 38611 18819
rect 41797 18785 41831 18819
rect 2973 18717 3007 18751
rect 5365 18717 5399 18751
rect 8309 18717 8343 18751
rect 12081 18717 12115 18751
rect 24041 18717 24075 18751
rect 27905 18717 27939 18751
rect 29193 18717 29227 18751
rect 30113 18717 30147 18751
rect 38393 18717 38427 18751
rect 48605 18717 48639 18751
rect 49341 18717 49375 18751
rect 1777 18649 1811 18683
rect 8125 18649 8159 18683
rect 10701 18649 10735 18683
rect 12909 18649 12943 18683
rect 13001 18649 13035 18683
rect 14565 18649 14599 18683
rect 17417 18649 17451 18683
rect 19349 18649 19383 18683
rect 20269 18649 20303 18683
rect 23765 18649 23799 18683
rect 26065 18649 26099 18683
rect 35909 18649 35943 18683
rect 39589 18649 39623 18683
rect 41521 18649 41555 18683
rect 11345 18581 11379 18615
rect 11621 18581 11655 18615
rect 12541 18581 12575 18615
rect 13921 18581 13955 18615
rect 16681 18581 16715 18615
rect 17325 18581 17359 18615
rect 18521 18581 18555 18615
rect 19625 18581 19659 18615
rect 20361 18581 20395 18615
rect 21465 18581 21499 18615
rect 21557 18581 21591 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 28365 18581 28399 18615
rect 28549 18581 28583 18615
rect 30481 18581 30515 18615
rect 30849 18581 30883 18615
rect 31217 18581 31251 18615
rect 31861 18581 31895 18615
rect 31953 18581 31987 18615
rect 33057 18581 33091 18615
rect 33701 18581 33735 18615
rect 34253 18581 34287 18615
rect 35173 18581 35207 18615
rect 37657 18581 37691 18615
rect 38485 18581 38519 18615
rect 40049 18581 40083 18615
rect 48421 18581 48455 18615
rect 3617 18377 3651 18411
rect 9781 18377 9815 18411
rect 10793 18377 10827 18411
rect 14289 18377 14323 18411
rect 17969 18377 18003 18411
rect 19073 18377 19107 18411
rect 26249 18377 26283 18411
rect 27537 18377 27571 18411
rect 27629 18377 27663 18411
rect 28733 18377 28767 18411
rect 30389 18377 30423 18411
rect 30849 18377 30883 18411
rect 32689 18377 32723 18411
rect 33057 18377 33091 18411
rect 35357 18377 35391 18411
rect 35909 18377 35943 18411
rect 36921 18377 36955 18411
rect 37289 18377 37323 18411
rect 40417 18377 40451 18411
rect 40877 18377 40911 18411
rect 48789 18377 48823 18411
rect 7665 18309 7699 18343
rect 13185 18309 13219 18343
rect 17233 18309 17267 18343
rect 17417 18309 17451 18343
rect 19901 18309 19935 18343
rect 22477 18309 22511 18343
rect 24133 18309 24167 18343
rect 28825 18309 28859 18343
rect 40785 18309 40819 18343
rect 2973 18241 3007 18275
rect 3433 18241 3467 18275
rect 4445 18241 4479 18275
rect 7849 18241 7883 18275
rect 9965 18241 9999 18275
rect 10885 18241 10919 18275
rect 13461 18241 13495 18275
rect 15209 18241 15243 18275
rect 16313 18241 16347 18275
rect 18337 18241 18371 18275
rect 22569 18241 22603 18275
rect 23305 18241 23339 18275
rect 25053 18241 25087 18275
rect 25145 18241 25179 18275
rect 26341 18241 26375 18275
rect 30481 18241 30515 18275
rect 31309 18241 31343 18275
rect 36277 18241 36311 18275
rect 36369 18241 36403 18275
rect 39773 18241 39807 18275
rect 48605 18241 48639 18275
rect 49341 18241 49375 18275
rect 1777 18173 1811 18207
rect 4169 18173 4203 18207
rect 10977 18173 11011 18207
rect 14381 18173 14415 18207
rect 14565 18173 14599 18207
rect 15669 18173 15703 18207
rect 16681 18173 16715 18207
rect 18429 18173 18463 18207
rect 18613 18173 18647 18207
rect 19349 18173 19383 18207
rect 19625 18173 19659 18207
rect 22661 18173 22695 18207
rect 25237 18173 25271 18207
rect 26433 18173 26467 18207
rect 27721 18173 27755 18207
rect 28917 18173 28951 18207
rect 30297 18173 30331 18207
rect 32413 18173 32447 18207
rect 32597 18173 32631 18207
rect 33609 18173 33643 18207
rect 33885 18173 33919 18207
rect 36553 18173 36587 18207
rect 39497 18173 39531 18207
rect 40969 18173 41003 18207
rect 13921 18105 13955 18139
rect 16129 18105 16163 18139
rect 16865 18105 16899 18139
rect 22109 18105 22143 18139
rect 24685 18105 24719 18139
rect 28365 18105 28399 18139
rect 37565 18105 37599 18139
rect 38025 18105 38059 18139
rect 10425 18037 10459 18071
rect 11713 18037 11747 18071
rect 15025 18037 15059 18071
rect 21373 18037 21407 18071
rect 25881 18037 25915 18071
rect 27169 18037 27203 18071
rect 29745 18037 29779 18071
rect 37657 18037 37691 18071
rect 40049 18037 40083 18071
rect 49157 18037 49191 18071
rect 10149 17833 10183 17867
rect 10609 17833 10643 17867
rect 12909 17833 12943 17867
rect 14289 17833 14323 17867
rect 17509 17833 17543 17867
rect 19441 17833 19475 17867
rect 23305 17833 23339 17867
rect 25789 17833 25823 17867
rect 26249 17833 26283 17867
rect 29101 17833 29135 17867
rect 29653 17833 29687 17867
rect 33885 17833 33919 17867
rect 40509 17833 40543 17867
rect 24593 17765 24627 17799
rect 34069 17765 34103 17799
rect 34345 17765 34379 17799
rect 38761 17765 38795 17799
rect 10333 17697 10367 17731
rect 12357 17697 12391 17731
rect 15761 17697 15795 17731
rect 16037 17697 16071 17731
rect 16865 17697 16899 17731
rect 18705 17697 18739 17731
rect 21741 17697 21775 17731
rect 22017 17697 22051 17731
rect 23949 17697 23983 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 28549 17697 28583 17731
rect 31493 17697 31527 17731
rect 31585 17697 31619 17731
rect 32965 17697 32999 17731
rect 33057 17697 33091 17731
rect 35817 17697 35851 17731
rect 38117 17697 38151 17731
rect 39221 17697 39255 17731
rect 40969 17697 41003 17731
rect 41061 17697 41095 17731
rect 2973 17629 3007 17663
rect 13093 17629 13127 17663
rect 13737 17629 13771 17663
rect 17141 17629 17175 17663
rect 17969 17629 18003 17663
rect 19625 17629 19659 17663
rect 25973 17629 26007 17663
rect 28825 17629 28859 17663
rect 31677 17629 31711 17663
rect 34437 17629 34471 17663
rect 37565 17629 37599 17663
rect 48605 17629 48639 17663
rect 49341 17629 49375 17663
rect 1777 17561 1811 17595
rect 12081 17561 12115 17595
rect 22293 17561 22327 17595
rect 22845 17561 22879 17595
rect 23673 17561 23707 17595
rect 26433 17561 26467 17595
rect 29377 17561 29411 17595
rect 29929 17561 29963 17595
rect 30757 17561 30791 17595
rect 37289 17561 37323 17595
rect 38393 17561 38427 17595
rect 40877 17561 40911 17595
rect 48789 17561 48823 17595
rect 13553 17493 13587 17527
rect 16497 17493 16531 17527
rect 17049 17493 17083 17527
rect 20269 17493 20303 17527
rect 23765 17493 23799 17527
rect 24961 17493 24995 17527
rect 27077 17493 27111 17527
rect 32045 17493 32079 17527
rect 32321 17493 32355 17527
rect 33149 17493 33183 17527
rect 33517 17493 33551 17527
rect 35081 17493 35115 17527
rect 35449 17493 35483 17527
rect 38301 17493 38335 17527
rect 39037 17493 39071 17527
rect 49157 17493 49191 17527
rect 11805 17289 11839 17323
rect 13093 17289 13127 17323
rect 14933 17289 14967 17323
rect 15577 17289 15611 17323
rect 19165 17289 19199 17323
rect 22661 17289 22695 17323
rect 24869 17289 24903 17323
rect 25329 17289 25363 17323
rect 27353 17289 27387 17323
rect 27721 17289 27755 17323
rect 29009 17289 29043 17323
rect 30113 17289 30147 17323
rect 30573 17289 30607 17323
rect 31309 17289 31343 17323
rect 31401 17289 31435 17323
rect 34069 17289 34103 17323
rect 37841 17289 37875 17323
rect 48421 17289 48455 17323
rect 11897 17221 11931 17255
rect 13001 17221 13035 17255
rect 14289 17221 14323 17255
rect 15945 17221 15979 17255
rect 17969 17221 18003 17255
rect 20637 17221 20671 17255
rect 22109 17221 22143 17255
rect 25973 17221 26007 17255
rect 28917 17221 28951 17255
rect 35541 17221 35575 17255
rect 37013 17221 37047 17255
rect 38577 17221 38611 17255
rect 40417 17221 40451 17255
rect 2973 17153 3007 17187
rect 10701 17153 10735 17187
rect 10793 17153 10827 17187
rect 15117 17153 15151 17187
rect 17049 17153 17083 17187
rect 18705 17153 18739 17187
rect 20913 17153 20947 17187
rect 24409 17153 24443 17187
rect 25237 17153 25271 17187
rect 30205 17153 30239 17187
rect 32321 17153 32355 17187
rect 36277 17153 36311 17187
rect 36369 17153 36403 17187
rect 37933 17153 37967 17187
rect 48605 17153 48639 17187
rect 49249 17153 49283 17187
rect 1777 17085 1811 17119
rect 9873 17085 9907 17119
rect 10609 17085 10643 17119
rect 12817 17085 12851 17119
rect 14105 17085 14139 17119
rect 16037 17085 16071 17119
rect 16129 17085 16163 17119
rect 22017 17085 22051 17119
rect 24133 17085 24167 17119
rect 25513 17085 25547 17119
rect 27813 17085 27847 17119
rect 27905 17085 27939 17119
rect 28733 17085 28767 17119
rect 29929 17085 29963 17119
rect 31125 17085 31159 17119
rect 32597 17085 32631 17119
rect 34805 17085 34839 17119
rect 36185 17085 36219 17119
rect 38025 17085 38059 17119
rect 40693 17085 40727 17119
rect 49065 17085 49099 17119
rect 9781 17017 9815 17051
rect 10149 17017 10183 17051
rect 11161 17017 11195 17051
rect 29377 17017 29411 17051
rect 37473 17017 37507 17051
rect 9505 16949 9539 16983
rect 12449 16949 12483 16983
rect 13461 16949 13495 16983
rect 13829 16949 13863 16983
rect 16957 16949 16991 16983
rect 17417 16949 17451 16983
rect 21189 16949 21223 16983
rect 21557 16949 21591 16983
rect 31769 16949 31803 16983
rect 36737 16949 36771 16983
rect 38945 16949 38979 16983
rect 40969 16949 41003 16983
rect 10425 16745 10459 16779
rect 21005 16745 21039 16779
rect 24777 16745 24811 16779
rect 29193 16745 29227 16779
rect 36277 16745 36311 16779
rect 41061 16745 41095 16779
rect 41245 16745 41279 16779
rect 48789 16745 48823 16779
rect 14197 16677 14231 16711
rect 28733 16677 28767 16711
rect 34437 16677 34471 16711
rect 41521 16677 41555 16711
rect 7941 16609 7975 16643
rect 11161 16609 11195 16643
rect 13185 16609 13219 16643
rect 13277 16609 13311 16643
rect 14565 16609 14599 16643
rect 16129 16609 16163 16643
rect 16221 16609 16255 16643
rect 18889 16609 18923 16643
rect 22477 16609 22511 16643
rect 22753 16609 22787 16643
rect 23765 16609 23799 16643
rect 23949 16609 23983 16643
rect 27077 16609 27111 16643
rect 27997 16609 28031 16643
rect 28273 16609 28307 16643
rect 28365 16609 28399 16643
rect 28641 16609 28675 16643
rect 29285 16609 29319 16643
rect 29837 16609 29871 16643
rect 30021 16609 30055 16643
rect 31125 16609 31159 16643
rect 31217 16609 31251 16643
rect 32229 16609 32263 16643
rect 35081 16609 35115 16643
rect 36737 16609 36771 16643
rect 36829 16609 36863 16643
rect 37289 16609 37323 16643
rect 39221 16609 39255 16643
rect 40233 16609 40267 16643
rect 2973 16541 3007 16575
rect 8125 16541 8159 16575
rect 12357 16541 12391 16575
rect 13369 16541 13403 16575
rect 14749 16541 14783 16575
rect 16037 16541 16071 16575
rect 20269 16541 20303 16575
rect 27353 16541 27387 16575
rect 35817 16541 35851 16575
rect 39497 16541 39531 16575
rect 48605 16541 48639 16575
rect 49341 16541 49375 16575
rect 1777 16473 1811 16507
rect 8033 16473 8067 16507
rect 10057 16473 10091 16507
rect 10517 16473 10551 16507
rect 11437 16473 11471 16507
rect 16681 16473 16715 16507
rect 18613 16473 18647 16507
rect 24593 16473 24627 16507
rect 30113 16473 30147 16507
rect 32505 16473 32539 16507
rect 40325 16473 40359 16507
rect 40417 16473 40451 16507
rect 8493 16405 8527 16439
rect 9045 16405 9079 16439
rect 11345 16405 11379 16439
rect 11805 16405 11839 16439
rect 12541 16405 12575 16439
rect 13737 16405 13771 16439
rect 14841 16405 14875 16439
rect 15209 16405 15243 16439
rect 15669 16405 15703 16439
rect 17141 16405 17175 16439
rect 19441 16405 19475 16439
rect 20085 16405 20119 16439
rect 20637 16405 20671 16439
rect 23305 16405 23339 16439
rect 23673 16405 23707 16439
rect 25605 16405 25639 16439
rect 27629 16405 27663 16439
rect 30481 16405 30515 16439
rect 31309 16405 31343 16439
rect 31677 16405 31711 16439
rect 33977 16405 34011 16439
rect 34345 16405 34379 16439
rect 36645 16405 36679 16439
rect 37749 16405 37783 16439
rect 40785 16405 40819 16439
rect 49157 16405 49191 16439
rect 8309 16201 8343 16235
rect 9229 16201 9263 16235
rect 11989 16201 12023 16235
rect 12449 16201 12483 16235
rect 13185 16201 13219 16235
rect 15945 16201 15979 16235
rect 17417 16201 17451 16235
rect 17785 16201 17819 16235
rect 30941 16201 30975 16235
rect 33793 16201 33827 16235
rect 40509 16201 40543 16235
rect 40969 16201 41003 16235
rect 13553 16133 13587 16167
rect 14841 16133 14875 16167
rect 17049 16133 17083 16167
rect 19441 16133 19475 16167
rect 34529 16133 34563 16167
rect 38485 16133 38519 16167
rect 2973 16065 3007 16099
rect 8217 16065 8251 16099
rect 9321 16065 9355 16099
rect 10425 16065 10459 16099
rect 11069 16065 11103 16099
rect 12357 16065 12391 16099
rect 14749 16065 14783 16099
rect 19165 16065 19199 16099
rect 23489 16065 23523 16099
rect 26341 16065 26375 16099
rect 26709 16065 26743 16099
rect 27537 16065 27571 16099
rect 27629 16065 27663 16099
rect 28365 16065 28399 16099
rect 30849 16065 30883 16099
rect 32597 16065 32631 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 36921 16065 36955 16099
rect 38209 16065 38243 16099
rect 40877 16065 40911 16099
rect 48789 16065 48823 16099
rect 49341 16065 49375 16099
rect 1777 15997 1811 16031
rect 8125 15997 8159 16031
rect 12633 15997 12667 16031
rect 13645 15997 13679 16031
rect 13737 15997 13771 16031
rect 14933 15997 14967 16031
rect 15669 15997 15703 16031
rect 15853 15997 15887 16031
rect 16773 15997 16807 16031
rect 17877 15997 17911 16031
rect 17969 15997 18003 16031
rect 23305 15997 23339 16031
rect 23397 15997 23431 16031
rect 24593 15997 24627 16031
rect 26065 15997 26099 16031
rect 27721 15997 27755 16031
rect 28641 15997 28675 16031
rect 30665 15997 30699 16031
rect 32505 15997 32539 16031
rect 33609 15997 33643 16031
rect 36645 15997 36679 16031
rect 37473 15997 37507 16031
rect 41061 15997 41095 16031
rect 8677 15929 8711 15963
rect 16313 15929 16347 15963
rect 20913 15929 20947 15963
rect 22753 15929 22787 15963
rect 23857 15929 23891 15963
rect 34713 15929 34747 15963
rect 49157 15929 49191 15963
rect 10517 15861 10551 15895
rect 10977 15861 11011 15895
rect 11621 15861 11655 15895
rect 14381 15861 14415 15895
rect 16957 15861 16991 15895
rect 18889 15861 18923 15895
rect 21281 15861 21315 15895
rect 27169 15861 27203 15895
rect 30113 15861 30147 15895
rect 31309 15861 31343 15895
rect 31677 15861 31711 15895
rect 31861 15861 31895 15895
rect 33057 15861 33091 15895
rect 34253 15861 34287 15895
rect 35173 15861 35207 15895
rect 39957 15861 39991 15895
rect 41613 15861 41647 15895
rect 10793 15657 10827 15691
rect 14289 15657 14323 15691
rect 16773 15657 16807 15691
rect 17877 15657 17911 15691
rect 18061 15657 18095 15691
rect 18981 15657 19015 15691
rect 19349 15657 19383 15691
rect 19901 15657 19935 15691
rect 21189 15657 21223 15691
rect 27077 15657 27111 15691
rect 34345 15657 34379 15691
rect 36645 15657 36679 15691
rect 37749 15657 37783 15691
rect 41797 15657 41831 15691
rect 42073 15657 42107 15691
rect 49157 15657 49191 15691
rect 18429 15589 18463 15623
rect 22477 15589 22511 15623
rect 32229 15589 32263 15623
rect 33425 15589 33459 15623
rect 12265 15521 12299 15555
rect 12541 15521 12575 15555
rect 13185 15521 13219 15555
rect 14933 15521 14967 15555
rect 16129 15521 16163 15555
rect 17325 15521 17359 15555
rect 20361 15521 20395 15555
rect 20545 15521 20579 15555
rect 21741 15521 21775 15555
rect 23765 15521 23799 15555
rect 25237 15521 25271 15555
rect 26433 15521 26467 15555
rect 27997 15521 28031 15555
rect 30481 15521 30515 15555
rect 32873 15521 32907 15555
rect 32965 15521 32999 15555
rect 34897 15521 34931 15555
rect 35173 15521 35207 15555
rect 39497 15521 39531 15555
rect 40049 15521 40083 15555
rect 40325 15521 40359 15555
rect 2973 15453 3007 15487
rect 13277 15453 13311 15487
rect 13369 15453 13403 15487
rect 14749 15453 14783 15487
rect 18613 15453 18647 15487
rect 23581 15453 23615 15487
rect 27813 15453 27847 15487
rect 28457 15453 28491 15487
rect 29009 15453 29043 15487
rect 48881 15453 48915 15487
rect 49341 15453 49375 15487
rect 1777 15385 1811 15419
rect 6377 15385 6411 15419
rect 6561 15385 6595 15419
rect 10517 15385 10551 15419
rect 15945 15385 15979 15419
rect 17141 15385 17175 15419
rect 17233 15385 17267 15419
rect 21557 15385 21591 15419
rect 23489 15385 23523 15419
rect 25053 15385 25087 15419
rect 26341 15385 26375 15419
rect 27905 15385 27939 15419
rect 28641 15385 28675 15419
rect 29193 15385 29227 15419
rect 30757 15385 30791 15419
rect 39221 15385 39255 15419
rect 9045 15317 9079 15351
rect 13737 15317 13771 15351
rect 14657 15317 14691 15351
rect 15577 15317 15611 15351
rect 16037 15317 16071 15351
rect 19533 15317 19567 15351
rect 20269 15317 20303 15351
rect 21649 15317 21683 15351
rect 22201 15317 22235 15351
rect 23121 15317 23155 15351
rect 24685 15317 24719 15351
rect 25145 15317 25179 15351
rect 25881 15317 25915 15351
rect 26249 15317 26283 15351
rect 26985 15317 27019 15351
rect 27445 15317 27479 15351
rect 29377 15317 29411 15351
rect 30021 15317 30055 15351
rect 33057 15317 33091 15351
rect 33885 15317 33919 15351
rect 37105 15317 37139 15351
rect 9689 15113 9723 15147
rect 9781 15113 9815 15147
rect 11897 15113 11931 15147
rect 13369 15113 13403 15147
rect 15577 15113 15611 15147
rect 15945 15113 15979 15147
rect 18337 15113 18371 15147
rect 18705 15113 18739 15147
rect 19533 15113 19567 15147
rect 22017 15113 22051 15147
rect 24133 15113 24167 15147
rect 27077 15113 27111 15147
rect 27537 15113 27571 15147
rect 29745 15113 29779 15147
rect 30573 15113 30607 15147
rect 31401 15113 31435 15147
rect 33885 15113 33919 15147
rect 35081 15113 35115 15147
rect 36277 15113 36311 15147
rect 40141 15113 40175 15147
rect 10885 15045 10919 15079
rect 11069 15045 11103 15079
rect 19901 15045 19935 15079
rect 21097 15045 21131 15079
rect 21833 15045 21867 15079
rect 23397 15045 23431 15079
rect 36185 15045 36219 15079
rect 37749 15045 37783 15079
rect 40049 15045 40083 15079
rect 1777 14977 1811 15011
rect 2973 14977 3007 15011
rect 12265 14977 12299 15011
rect 12357 14977 12391 15011
rect 15117 14977 15151 15011
rect 17233 14977 17267 15011
rect 19993 14977 20027 15011
rect 23305 14977 23339 15011
rect 24501 14977 24535 15011
rect 25329 14977 25363 15011
rect 25605 14977 25639 15011
rect 26249 14977 26283 15011
rect 27261 14977 27295 15011
rect 27997 14977 28031 15011
rect 32689 14977 32723 15011
rect 37473 14977 37507 15011
rect 40877 14977 40911 15011
rect 48789 14977 48823 15011
rect 49341 14977 49375 15011
rect 9597 14909 9631 14943
rect 11621 14909 11655 14943
rect 12449 14909 12483 14943
rect 14841 14909 14875 14943
rect 16037 14909 16071 14943
rect 16129 14909 16163 14943
rect 17325 14909 17359 14943
rect 17417 14909 17451 14943
rect 18061 14909 18095 14943
rect 18797 14909 18831 14943
rect 18889 14909 18923 14943
rect 20177 14909 20211 14943
rect 21189 14909 21223 14943
rect 21281 14909 21315 14943
rect 23581 14909 23615 14943
rect 24593 14909 24627 14943
rect 24685 14909 24719 14943
rect 26341 14909 26375 14943
rect 26433 14909 26467 14943
rect 28273 14909 28307 14943
rect 30665 14909 30699 14943
rect 30757 14909 30791 14943
rect 32781 14909 32815 14943
rect 32873 14909 32907 14943
rect 33701 14909 33735 14943
rect 33793 14909 33827 14943
rect 34897 14909 34931 14943
rect 34989 14909 35023 14943
rect 36001 14909 36035 14943
rect 37013 14909 37047 14943
rect 39221 14909 39255 14943
rect 40233 14909 40267 14943
rect 10149 14841 10183 14875
rect 20729 14841 20763 14875
rect 22937 14841 22971 14875
rect 25881 14841 25915 14875
rect 27445 14841 27479 14875
rect 32321 14841 32355 14875
rect 39681 14841 39715 14875
rect 49157 14841 49191 14875
rect 10609 14773 10643 14807
rect 13001 14773 13035 14807
rect 16865 14773 16899 14807
rect 25145 14773 25179 14807
rect 30205 14773 30239 14807
rect 31861 14773 31895 14807
rect 34253 14773 34287 14807
rect 35449 14773 35483 14807
rect 36645 14773 36679 14807
rect 41061 14773 41095 14807
rect 11805 14569 11839 14603
rect 13001 14569 13035 14603
rect 14197 14569 14231 14603
rect 14473 14569 14507 14603
rect 18153 14569 18187 14603
rect 24593 14569 24627 14603
rect 25605 14569 25639 14603
rect 30481 14569 30515 14603
rect 36645 14569 36679 14603
rect 39957 14569 39991 14603
rect 40049 14569 40083 14603
rect 10241 14501 10275 14535
rect 22845 14501 22879 14535
rect 31677 14501 31711 14535
rect 34069 14501 34103 14535
rect 49065 14501 49099 14535
rect 1777 14433 1811 14467
rect 12449 14433 12483 14467
rect 13553 14433 13587 14467
rect 15117 14433 15151 14467
rect 16957 14433 16991 14467
rect 17509 14433 17543 14467
rect 18705 14433 18739 14467
rect 20085 14433 20119 14467
rect 21097 14433 21131 14467
rect 21373 14433 21407 14467
rect 27997 14433 28031 14467
rect 29929 14433 29963 14467
rect 31033 14433 31067 14467
rect 32321 14433 32355 14467
rect 33425 14433 33459 14467
rect 34345 14433 34379 14467
rect 34897 14433 34931 14467
rect 38853 14433 38887 14467
rect 2973 14365 3007 14399
rect 9505 14365 9539 14399
rect 9689 14365 9723 14399
rect 14933 14365 14967 14399
rect 18613 14365 18647 14399
rect 19901 14365 19935 14399
rect 27353 14365 27387 14399
rect 30113 14365 30147 14399
rect 31309 14365 31343 14399
rect 33609 14365 33643 14399
rect 33701 14365 33735 14399
rect 39313 14365 39347 14399
rect 48605 14365 48639 14399
rect 49249 14365 49283 14399
rect 10425 14297 10459 14331
rect 11253 14297 11287 14331
rect 12173 14297 12207 14331
rect 13369 14297 13403 14331
rect 15945 14297 15979 14331
rect 16773 14297 16807 14331
rect 17877 14297 17911 14331
rect 19993 14297 20027 14331
rect 27077 14297 27111 14331
rect 28181 14297 28215 14331
rect 31217 14297 31251 14331
rect 32505 14297 32539 14331
rect 35173 14297 35207 14331
rect 38577 14297 38611 14331
rect 11161 14229 11195 14263
rect 12265 14229 12299 14263
rect 13461 14229 13495 14263
rect 14841 14229 14875 14263
rect 16405 14229 16439 14263
rect 16865 14229 16899 14263
rect 17601 14229 17635 14263
rect 18521 14229 18555 14263
rect 19533 14229 19567 14263
rect 20545 14229 20579 14263
rect 20729 14229 20763 14263
rect 23213 14229 23247 14263
rect 23489 14229 23523 14263
rect 23857 14229 23891 14263
rect 24409 14229 24443 14263
rect 25145 14229 25179 14263
rect 28089 14229 28123 14263
rect 28549 14229 28583 14263
rect 29009 14229 29043 14263
rect 30021 14229 30055 14263
rect 32413 14229 32447 14263
rect 32873 14229 32907 14263
rect 37105 14229 37139 14263
rect 39497 14229 39531 14263
rect 48697 14229 48731 14263
rect 9965 14025 9999 14059
rect 10425 14025 10459 14059
rect 11989 14025 12023 14059
rect 15025 14025 15059 14059
rect 15577 14025 15611 14059
rect 17141 14025 17175 14059
rect 17509 14025 17543 14059
rect 17601 14025 17635 14059
rect 18337 14025 18371 14059
rect 18705 14025 18739 14059
rect 19441 14025 19475 14059
rect 21465 14025 21499 14059
rect 24869 14025 24903 14059
rect 27629 14025 27663 14059
rect 31769 14025 31803 14059
rect 34897 14025 34931 14059
rect 35265 14025 35299 14059
rect 36461 14025 36495 14059
rect 37841 14025 37875 14059
rect 38209 14025 38243 14059
rect 45845 14025 45879 14059
rect 48421 14025 48455 14059
rect 49157 14025 49191 14059
rect 1777 13957 1811 13991
rect 10701 13957 10735 13991
rect 13277 13957 13311 13991
rect 16037 13957 16071 13991
rect 23489 13957 23523 13991
rect 26341 13957 26375 13991
rect 36093 13957 36127 13991
rect 37749 13957 37783 13991
rect 38577 13957 38611 13991
rect 38945 13957 38979 13991
rect 45017 13957 45051 13991
rect 48145 13957 48179 13991
rect 49249 13957 49283 13991
rect 2973 13889 3007 13923
rect 3525 13889 3559 13923
rect 3985 13889 4019 13923
rect 11161 13889 11195 13923
rect 12081 13889 12115 13923
rect 15945 13889 15979 13923
rect 16865 13889 16899 13923
rect 18797 13889 18831 13923
rect 26617 13889 26651 13923
rect 28917 13889 28951 13923
rect 31125 13889 31159 13923
rect 34805 13889 34839 13923
rect 36921 13889 36955 13923
rect 45661 13889 45695 13923
rect 48605 13889 48639 13923
rect 3709 13821 3743 13855
rect 11897 13821 11931 13855
rect 13001 13821 13035 13855
rect 14749 13821 14783 13855
rect 16129 13821 16163 13855
rect 17785 13821 17819 13855
rect 18889 13821 18923 13855
rect 19717 13821 19751 13855
rect 19993 13821 20027 13855
rect 22017 13821 22051 13855
rect 23765 13821 23799 13855
rect 24225 13821 24259 13855
rect 29377 13821 29411 13855
rect 30849 13821 30883 13855
rect 32321 13821 32355 13855
rect 34069 13821 34103 13855
rect 34621 13821 34655 13855
rect 35909 13821 35943 13855
rect 36001 13821 36035 13855
rect 36737 13821 36771 13855
rect 37657 13821 37691 13855
rect 45201 13821 45235 13855
rect 12449 13685 12483 13719
rect 15301 13685 15335 13719
rect 33811 13685 33845 13719
rect 13737 13481 13771 13515
rect 13921 13481 13955 13515
rect 18153 13481 18187 13515
rect 19441 13481 19475 13515
rect 20453 13481 20487 13515
rect 20913 13481 20947 13515
rect 22109 13481 22143 13515
rect 24041 13481 24075 13515
rect 25605 13481 25639 13515
rect 26709 13481 26743 13515
rect 27445 13481 27479 13515
rect 27721 13481 27755 13515
rect 27813 13481 27847 13515
rect 28181 13481 28215 13515
rect 29193 13481 29227 13515
rect 35633 13481 35667 13515
rect 36001 13481 36035 13515
rect 38209 13481 38243 13515
rect 38577 13481 38611 13515
rect 39589 13481 39623 13515
rect 14289 13413 14323 13447
rect 14841 13413 14875 13447
rect 31125 13413 31159 13447
rect 33333 13413 33367 13447
rect 36093 13413 36127 13447
rect 1777 13345 1811 13379
rect 10793 13345 10827 13379
rect 12541 13345 12575 13379
rect 13093 13345 13127 13379
rect 15393 13345 15427 13379
rect 15485 13345 15519 13379
rect 16405 13345 16439 13379
rect 16681 13345 16715 13379
rect 19901 13345 19935 13379
rect 21465 13345 21499 13379
rect 22753 13345 22787 13379
rect 23489 13345 23523 13379
rect 23581 13345 23615 13379
rect 25053 13345 25087 13379
rect 28641 13345 28675 13379
rect 29837 13345 29871 13379
rect 30021 13345 30055 13379
rect 33885 13345 33919 13379
rect 34345 13345 34379 13379
rect 35081 13345 35115 13379
rect 36737 13345 36771 13379
rect 2973 13277 3007 13311
rect 14473 13277 14507 13311
rect 15577 13277 15611 13311
rect 25237 13277 25271 13311
rect 28825 13277 28859 13311
rect 30113 13277 30147 13311
rect 32873 13277 32907 13311
rect 36461 13277 36495 13311
rect 41337 13277 41371 13311
rect 47961 13277 47995 13311
rect 49157 13277 49191 13311
rect 11069 13209 11103 13243
rect 18889 13209 18923 13243
rect 20085 13209 20119 13243
rect 21373 13209 21407 13243
rect 22477 13209 22511 13243
rect 23673 13209 23707 13243
rect 26065 13209 26099 13243
rect 32597 13209 32631 13243
rect 35173 13209 35207 13243
rect 35265 13209 35299 13243
rect 10517 13141 10551 13175
rect 15945 13141 15979 13175
rect 19993 13141 20027 13175
rect 21281 13141 21315 13175
rect 22569 13141 22603 13175
rect 24501 13141 24535 13175
rect 25145 13141 25179 13175
rect 28733 13141 28767 13175
rect 30481 13141 30515 13175
rect 33701 13141 33735 13175
rect 33793 13141 33827 13175
rect 41521 13141 41555 13175
rect 3065 12937 3099 12971
rect 10977 12937 11011 12971
rect 11161 12937 11195 12971
rect 11989 12937 12023 12971
rect 12081 12937 12115 12971
rect 12725 12937 12759 12971
rect 13093 12937 13127 12971
rect 15209 12937 15243 12971
rect 15853 12937 15887 12971
rect 20729 12937 20763 12971
rect 21189 12937 21223 12971
rect 22937 12937 22971 12971
rect 26065 12937 26099 12971
rect 26341 12937 26375 12971
rect 26709 12937 26743 12971
rect 31769 12937 31803 12971
rect 33425 12937 33459 12971
rect 36461 12937 36495 12971
rect 1685 12869 1719 12903
rect 2145 12869 2179 12903
rect 15945 12869 15979 12903
rect 18705 12869 18739 12903
rect 25329 12869 25363 12903
rect 29653 12869 29687 12903
rect 30297 12869 30331 12903
rect 32689 12869 32723 12903
rect 34805 12869 34839 12903
rect 35817 12869 35851 12903
rect 2881 12801 2915 12835
rect 3341 12801 3375 12835
rect 16957 12801 16991 12835
rect 17877 12801 17911 12835
rect 19625 12801 19659 12835
rect 21097 12801 21131 12835
rect 23029 12801 23063 12835
rect 25605 12801 25639 12835
rect 29193 12801 29227 12835
rect 30021 12801 30055 12835
rect 32597 12801 32631 12835
rect 34069 12801 34103 12835
rect 36645 12801 36679 12835
rect 37473 12801 37507 12835
rect 40049 12801 40083 12835
rect 40509 12801 40543 12835
rect 45937 12801 45971 12835
rect 47961 12801 47995 12835
rect 49157 12801 49191 12835
rect 1869 12733 1903 12767
rect 11805 12733 11839 12767
rect 14565 12733 14599 12767
rect 14841 12733 14875 12767
rect 15761 12733 15795 12767
rect 17417 12733 17451 12767
rect 19717 12733 19751 12767
rect 19901 12733 19935 12767
rect 21281 12733 21315 12767
rect 22017 12733 22051 12767
rect 22753 12733 22787 12767
rect 23857 12733 23891 12767
rect 25881 12733 25915 12767
rect 27169 12733 27203 12767
rect 28917 12733 28951 12767
rect 32413 12733 32447 12767
rect 35541 12733 35575 12767
rect 35725 12733 35759 12767
rect 37749 12733 37783 12767
rect 39497 12733 39531 12767
rect 16681 12665 16715 12699
rect 19257 12665 19291 12699
rect 23397 12665 23431 12699
rect 33057 12665 33091 12699
rect 36185 12665 36219 12699
rect 40233 12665 40267 12699
rect 11253 12597 11287 12631
rect 12449 12597 12483 12631
rect 16313 12597 16347 12631
rect 20361 12597 20395 12631
rect 26433 12597 26467 12631
rect 33609 12597 33643 12631
rect 33793 12597 33827 12631
rect 36829 12597 36863 12631
rect 37013 12597 37047 12631
rect 46121 12597 46155 12631
rect 11253 12393 11287 12427
rect 16405 12393 16439 12427
rect 19441 12393 19475 12427
rect 21649 12393 21683 12427
rect 23305 12393 23339 12427
rect 27721 12393 27755 12427
rect 31861 12393 31895 12427
rect 33885 12393 33919 12427
rect 39313 12393 39347 12427
rect 26341 12325 26375 12359
rect 34253 12325 34287 12359
rect 39037 12325 39071 12359
rect 39497 12325 39531 12359
rect 40325 12325 40359 12359
rect 2421 12257 2455 12291
rect 2697 12257 2731 12291
rect 9505 12257 9539 12291
rect 11713 12257 11747 12291
rect 13737 12257 13771 12291
rect 16129 12257 16163 12291
rect 17417 12257 17451 12291
rect 19993 12257 20027 12291
rect 20637 12257 20671 12291
rect 21097 12257 21131 12291
rect 22293 12257 22327 12291
rect 23765 12257 23799 12291
rect 23949 12257 23983 12291
rect 27077 12257 27111 12291
rect 28457 12257 28491 12291
rect 29745 12257 29779 12291
rect 32413 12257 32447 12291
rect 35173 12257 35207 12291
rect 37197 12257 37231 12291
rect 37381 12257 37415 12291
rect 38393 12257 38427 12291
rect 38577 12257 38611 12291
rect 49157 12257 49191 12291
rect 2145 12189 2179 12223
rect 17141 12189 17175 12223
rect 17233 12189 17267 12223
rect 19809 12189 19843 12223
rect 21189 12189 21223 12223
rect 21281 12189 21315 12223
rect 24593 12189 24627 12223
rect 26709 12189 26743 12223
rect 32137 12189 32171 12223
rect 34897 12189 34931 12223
rect 40785 12189 40819 12223
rect 41429 12189 41463 12223
rect 45937 12189 45971 12223
rect 47961 12189 47995 12223
rect 9781 12121 9815 12155
rect 11989 12121 12023 12155
rect 15853 12121 15887 12155
rect 18153 12121 18187 12155
rect 18889 12121 18923 12155
rect 22385 12121 22419 12155
rect 22477 12121 22511 12155
rect 23673 12121 23707 12155
rect 24869 12121 24903 12155
rect 29193 12121 29227 12155
rect 30021 12121 30055 12155
rect 40141 12121 40175 12155
rect 14381 12053 14415 12087
rect 16773 12053 16807 12087
rect 19901 12053 19935 12087
rect 22845 12053 22879 12087
rect 27261 12053 27295 12087
rect 27353 12053 27387 12087
rect 31493 12053 31527 12087
rect 34345 12053 34379 12087
rect 36645 12053 36679 12087
rect 37473 12053 37507 12087
rect 37841 12053 37875 12087
rect 38669 12053 38703 12087
rect 40969 12053 41003 12087
rect 41613 12053 41647 12087
rect 46121 12053 46155 12087
rect 2513 11849 2547 11883
rect 11621 11849 11655 11883
rect 12081 11849 12115 11883
rect 12725 11849 12759 11883
rect 13369 11849 13403 11883
rect 14197 11849 14231 11883
rect 14289 11849 14323 11883
rect 15485 11849 15519 11883
rect 16497 11849 16531 11883
rect 26617 11849 26651 11883
rect 27905 11849 27939 11883
rect 31493 11849 31527 11883
rect 31861 11849 31895 11883
rect 32597 11849 32631 11883
rect 32689 11849 32723 11883
rect 34805 11849 34839 11883
rect 37749 11849 37783 11883
rect 38669 11849 38703 11883
rect 39129 11849 39163 11883
rect 21189 11781 21223 11815
rect 24225 11781 24259 11815
rect 26157 11781 26191 11815
rect 27537 11781 27571 11815
rect 30021 11781 30055 11815
rect 39957 11781 39991 11815
rect 40601 11781 40635 11815
rect 45109 11781 45143 11815
rect 49157 11781 49191 11815
rect 1593 11713 1627 11747
rect 2329 11713 2363 11747
rect 13553 11713 13587 11747
rect 19257 11713 19291 11747
rect 19901 11713 19935 11747
rect 21097 11713 21131 11747
rect 22293 11713 22327 11747
rect 22569 11713 22603 11747
rect 31125 11713 31159 11747
rect 33793 11713 33827 11747
rect 33885 11713 33919 11747
rect 37841 11713 37875 11747
rect 39037 11713 39071 11747
rect 40417 11713 40451 11747
rect 47961 11713 47995 11747
rect 2789 11645 2823 11679
rect 12817 11645 12851 11679
rect 12909 11645 12943 11679
rect 14013 11645 14047 11679
rect 15577 11645 15611 11679
rect 15761 11645 15795 11679
rect 16865 11645 16899 11679
rect 18337 11645 18371 11679
rect 18613 11645 18647 11679
rect 19717 11645 19751 11679
rect 19809 11645 19843 11679
rect 21373 11645 21407 11679
rect 22109 11645 22143 11679
rect 23397 11645 23431 11679
rect 23949 11645 23983 11679
rect 25697 11645 25731 11679
rect 27261 11645 27295 11679
rect 27445 11645 27479 11679
rect 28549 11645 28583 11679
rect 30297 11645 30331 11679
rect 30849 11645 30883 11679
rect 31033 11645 31067 11679
rect 32505 11645 32539 11679
rect 33609 11645 33643 11679
rect 34529 11645 34563 11679
rect 35173 11645 35207 11679
rect 35449 11645 35483 11679
rect 37565 11645 37599 11679
rect 39221 11645 39255 11679
rect 1777 11577 1811 11611
rect 14657 11577 14691 11611
rect 19073 11577 19107 11611
rect 20269 11577 20303 11611
rect 20729 11577 20763 11611
rect 34253 11577 34287 11611
rect 36921 11577 36955 11611
rect 40141 11577 40175 11611
rect 45293 11577 45327 11611
rect 12357 11509 12391 11543
rect 15117 11509 15151 11543
rect 16313 11509 16347 11543
rect 21925 11509 21959 11543
rect 33057 11509 33091 11543
rect 38209 11509 38243 11543
rect 2145 11305 2179 11339
rect 14381 11305 14415 11339
rect 16313 11305 16347 11339
rect 19073 11305 19107 11339
rect 19257 11305 19291 11339
rect 19533 11305 19567 11339
rect 20453 11305 20487 11339
rect 21943 11305 21977 11339
rect 23305 11305 23339 11339
rect 26341 11305 26375 11339
rect 29009 11305 29043 11339
rect 34713 11305 34747 11339
rect 38393 11305 38427 11339
rect 1777 11237 1811 11271
rect 16773 11237 16807 11271
rect 17969 11237 18003 11271
rect 28641 11237 28675 11271
rect 30481 11237 30515 11271
rect 32873 11237 32907 11271
rect 38761 11237 38795 11271
rect 39589 11237 39623 11271
rect 40969 11237 41003 11271
rect 10977 11169 11011 11203
rect 12449 11169 12483 11203
rect 14841 11169 14875 11203
rect 15025 11169 15059 11203
rect 15761 11169 15795 11203
rect 15853 11169 15887 11203
rect 17417 11169 17451 11203
rect 18521 11169 18555 11203
rect 19993 11169 20027 11203
rect 23949 11169 23983 11203
rect 24869 11169 24903 11203
rect 29193 11169 29227 11203
rect 29285 11169 29319 11203
rect 29929 11169 29963 11203
rect 34069 11169 34103 11203
rect 37749 11169 37783 11203
rect 49157 11169 49191 11203
rect 1593 11101 1627 11135
rect 2329 11101 2363 11135
rect 12725 11101 12759 11135
rect 13737 11101 13771 11135
rect 17233 11101 17267 11135
rect 22201 11101 22235 11135
rect 24593 11101 24627 11135
rect 26893 11101 26927 11135
rect 31125 11101 31159 11135
rect 33333 11101 33367 11135
rect 38209 11101 38243 11135
rect 40141 11101 40175 11135
rect 40785 11101 40819 11135
rect 45661 11101 45695 11135
rect 47961 11101 47995 11135
rect 13001 11033 13035 11067
rect 15945 11033 15979 11067
rect 17141 11033 17175 11067
rect 23673 11033 23707 11067
rect 27169 11033 27203 11067
rect 30021 11033 30055 11067
rect 31401 11033 31435 11067
rect 35725 11033 35759 11067
rect 37473 11033 37507 11067
rect 40325 11033 40359 11067
rect 45845 11033 45879 11067
rect 13277 10965 13311 10999
rect 14749 10965 14783 10999
rect 18337 10965 18371 10999
rect 18429 10965 18463 10999
rect 22661 10965 22695 10999
rect 23765 10965 23799 10999
rect 30113 10965 30147 10999
rect 30757 10965 30791 10999
rect 1777 10761 1811 10795
rect 12541 10761 12575 10795
rect 13185 10761 13219 10795
rect 14381 10761 14415 10795
rect 15945 10761 15979 10795
rect 17141 10761 17175 10795
rect 19533 10761 19567 10795
rect 21097 10761 21131 10795
rect 24225 10761 24259 10795
rect 25881 10761 25915 10795
rect 26433 10761 26467 10795
rect 31401 10761 31435 10795
rect 33885 10761 33919 10795
rect 36829 10761 36863 10795
rect 14841 10693 14875 10727
rect 17509 10693 17543 10727
rect 19993 10693 20027 10727
rect 21189 10693 21223 10727
rect 28549 10693 28583 10727
rect 28825 10693 28859 10727
rect 33425 10693 33459 10727
rect 39773 10693 39807 10727
rect 40233 10693 40267 10727
rect 49157 10693 49191 10727
rect 1593 10625 1627 10659
rect 2329 10625 2363 10659
rect 2881 10625 2915 10659
rect 13553 10625 13587 10659
rect 14749 10625 14783 10659
rect 16865 10625 16899 10659
rect 18705 10625 18739 10659
rect 18797 10625 18831 10659
rect 19901 10625 19935 10659
rect 24593 10625 24627 10659
rect 25421 10625 25455 10659
rect 26341 10625 26375 10659
rect 26801 10625 26835 10659
rect 27537 10625 27571 10659
rect 30573 10625 30607 10659
rect 32689 10625 32723 10659
rect 35633 10625 35667 10659
rect 36461 10625 36495 10659
rect 47961 10625 47995 10659
rect 3065 10557 3099 10591
rect 12725 10557 12759 10591
rect 13645 10557 13679 10591
rect 13829 10557 13863 10591
rect 14933 10557 14967 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 17601 10557 17635 10591
rect 17693 10557 17727 10591
rect 18889 10557 18923 10591
rect 20177 10557 20211 10591
rect 21373 10557 21407 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24685 10557 24719 10591
rect 24869 10557 24903 10591
rect 27261 10557 27295 10591
rect 27445 10557 27479 10591
rect 29561 10557 29595 10591
rect 30389 10557 30423 10591
rect 30481 10557 30515 10591
rect 32413 10557 32447 10591
rect 32597 10557 32631 10591
rect 35357 10557 35391 10591
rect 36185 10557 36219 10591
rect 36369 10557 36403 10591
rect 37289 10557 37323 10591
rect 37473 10557 37507 10591
rect 2513 10489 2547 10523
rect 26065 10489 26099 10523
rect 27905 10489 27939 10523
rect 33057 10489 33091 10523
rect 39957 10489 39991 10523
rect 12265 10421 12299 10455
rect 12909 10421 12943 10455
rect 15577 10421 15611 10455
rect 18337 10421 18371 10455
rect 20729 10421 20763 10455
rect 23765 10421 23799 10455
rect 30941 10421 30975 10455
rect 31953 10421 31987 10455
rect 13461 10217 13495 10251
rect 16497 10217 16531 10251
rect 18153 10217 18187 10251
rect 20269 10217 20303 10251
rect 24593 10217 24627 10251
rect 28733 10217 28767 10251
rect 30389 10217 30423 10251
rect 36645 10217 36679 10251
rect 36921 10217 36955 10251
rect 13921 10149 13955 10183
rect 26709 10149 26743 10183
rect 29285 10149 29319 10183
rect 2145 10081 2179 10115
rect 12909 10081 12943 10115
rect 13001 10081 13035 10115
rect 17417 10081 17451 10115
rect 17601 10081 17635 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 19717 10081 19751 10115
rect 21741 10081 21775 10115
rect 23765 10081 23799 10115
rect 26065 10081 26099 10115
rect 26341 10081 26375 10115
rect 26985 10081 27019 10115
rect 29929 10081 29963 10115
rect 32137 10081 32171 10115
rect 32689 10081 32723 10115
rect 32873 10081 32907 10115
rect 35173 10081 35207 10115
rect 40601 10081 40635 10115
rect 49157 10081 49191 10115
rect 2421 10013 2455 10047
rect 13093 10013 13127 10047
rect 16037 10013 16071 10047
rect 18521 10013 18555 10047
rect 22017 10013 22051 10047
rect 23213 10013 23247 10047
rect 33793 10013 33827 10047
rect 34897 10013 34931 10047
rect 38301 10013 38335 10047
rect 38761 10013 38795 10047
rect 40141 10013 40175 10047
rect 40325 10013 40359 10047
rect 46121 10013 46155 10047
rect 47961 10013 47995 10047
rect 15761 9945 15795 9979
rect 22477 9945 22511 9979
rect 23857 9945 23891 9979
rect 27261 9945 27295 9979
rect 31861 9945 31895 9979
rect 32965 9945 32999 9979
rect 44373 9945 44407 9979
rect 44557 9945 44591 9979
rect 47317 9945 47351 9979
rect 12449 9877 12483 9911
rect 14289 9877 14323 9911
rect 16589 9877 16623 9911
rect 16957 9877 16991 9911
rect 17325 9877 17359 9911
rect 24041 9877 24075 9911
rect 29009 9877 29043 9911
rect 33333 9877 33367 9911
rect 38393 9877 38427 9911
rect 2145 9673 2179 9707
rect 21097 9673 21131 9707
rect 22293 9673 22327 9707
rect 31769 9673 31803 9707
rect 32873 9673 32907 9707
rect 35633 9673 35667 9707
rect 36185 9673 36219 9707
rect 12449 9605 12483 9639
rect 13369 9605 13403 9639
rect 16129 9605 16163 9639
rect 16313 9605 16347 9639
rect 16865 9605 16899 9639
rect 19625 9605 19659 9639
rect 21373 9605 21407 9639
rect 29009 9605 29043 9639
rect 49157 9605 49191 9639
rect 1593 9537 1627 9571
rect 2329 9537 2363 9571
rect 12541 9537 12575 9571
rect 15393 9537 15427 9571
rect 15853 9537 15887 9571
rect 22661 9537 22695 9571
rect 22753 9537 22787 9571
rect 25237 9537 25271 9571
rect 26065 9537 26099 9571
rect 32965 9537 32999 9571
rect 33885 9537 33919 9571
rect 47961 9537 47995 9571
rect 12265 9469 12299 9503
rect 15117 9469 15151 9503
rect 18613 9469 18647 9503
rect 18889 9469 18923 9503
rect 19349 9469 19383 9503
rect 22937 9469 22971 9503
rect 24961 9469 24995 9503
rect 25881 9469 25915 9503
rect 25973 9469 26007 9503
rect 27537 9469 27571 9503
rect 29285 9469 29319 9503
rect 29745 9469 29779 9503
rect 30021 9469 30055 9503
rect 31493 9469 31527 9503
rect 32689 9469 32723 9503
rect 34161 9469 34195 9503
rect 35909 9469 35943 9503
rect 1777 9401 1811 9435
rect 26433 9401 26467 9435
rect 12909 9333 12943 9367
rect 15669 9333 15703 9367
rect 16405 9333 16439 9367
rect 21557 9333 21591 9367
rect 21833 9333 21867 9367
rect 23489 9333 23523 9367
rect 32137 9333 32171 9367
rect 33333 9333 33367 9367
rect 1777 9129 1811 9163
rect 16405 9129 16439 9163
rect 17889 9129 17923 9163
rect 19441 9129 19475 9163
rect 22293 9129 22327 9163
rect 24501 9129 24535 9163
rect 25605 9129 25639 9163
rect 32873 9129 32907 9163
rect 33057 9129 33091 9163
rect 34069 9129 34103 9163
rect 30757 9061 30791 9095
rect 36737 9061 36771 9095
rect 2881 8993 2915 9027
rect 15301 8993 15335 9027
rect 15485 8993 15519 9027
rect 18153 8993 18187 9027
rect 20913 8993 20947 9027
rect 23765 8993 23799 9027
rect 24041 8993 24075 9027
rect 24685 8993 24719 9027
rect 24869 8993 24903 9027
rect 25421 8993 25455 9027
rect 28365 8993 28399 9027
rect 32505 8993 32539 9027
rect 33517 8993 33551 9027
rect 33609 8993 33643 9027
rect 34989 8993 35023 9027
rect 49157 8993 49191 9027
rect 2329 8925 2363 8959
rect 3065 8925 3099 8959
rect 14289 8925 14323 8959
rect 15577 8925 15611 8959
rect 18705 8925 18739 8959
rect 21189 8925 21223 8959
rect 36553 8925 36587 8959
rect 37657 8925 37691 8959
rect 39865 8925 39899 8959
rect 47961 8925 47995 8959
rect 1685 8857 1719 8891
rect 28549 8857 28583 8891
rect 29745 8857 29779 8891
rect 32229 8857 32263 8891
rect 35265 8857 35299 8891
rect 39313 8857 39347 8891
rect 39497 8857 39531 8891
rect 2513 8789 2547 8823
rect 14473 8789 14507 8823
rect 14933 8789 14967 8823
rect 15945 8789 15979 8823
rect 21833 8789 21867 8823
rect 25697 8789 25731 8823
rect 27813 8789 27847 8823
rect 28457 8789 28491 8823
rect 28917 8789 28951 8823
rect 30297 8789 30331 8823
rect 33701 8789 33735 8823
rect 34345 8789 34379 8823
rect 35173 8789 35207 8823
rect 35633 8789 35667 8823
rect 37841 8789 37875 8823
rect 15761 8585 15795 8619
rect 16221 8585 16255 8619
rect 18613 8585 18647 8619
rect 19717 8585 19751 8619
rect 22017 8585 22051 8619
rect 24133 8585 24167 8619
rect 31401 8585 31435 8619
rect 31769 8585 31803 8619
rect 34069 8585 34103 8619
rect 34345 8585 34379 8619
rect 37657 8585 37691 8619
rect 13921 8517 13955 8551
rect 17141 8517 17175 8551
rect 21189 8517 21223 8551
rect 29101 8517 29135 8551
rect 34713 8517 34747 8551
rect 44189 8517 44223 8551
rect 44373 8517 44407 8551
rect 49157 8517 49191 8551
rect 2145 8449 2179 8483
rect 13645 8449 13679 8483
rect 16865 8449 16899 8483
rect 23765 8449 23799 8483
rect 32321 8449 32355 8483
rect 37473 8449 37507 8483
rect 38945 8449 38979 8483
rect 40325 8449 40359 8483
rect 40785 8449 40819 8483
rect 45845 8449 45879 8483
rect 47961 8449 47995 8483
rect 2421 8381 2455 8415
rect 15393 8381 15427 8415
rect 19073 8381 19107 8415
rect 21465 8381 21499 8415
rect 23489 8381 23523 8415
rect 28825 8381 28859 8415
rect 31217 8381 31251 8415
rect 31309 8381 31343 8415
rect 32597 8381 32631 8415
rect 40509 8381 40543 8415
rect 46857 8381 46891 8415
rect 30573 8313 30607 8347
rect 34529 8313 34563 8347
rect 39129 8313 39163 8347
rect 2145 8041 2179 8075
rect 18981 8041 19015 8075
rect 19441 8041 19475 8075
rect 22017 8041 22051 8075
rect 30389 8041 30423 8075
rect 31769 8041 31803 8075
rect 15761 7973 15795 8007
rect 33057 7973 33091 8007
rect 16773 7905 16807 7939
rect 16957 7905 16991 7939
rect 18061 7905 18095 7939
rect 20913 7905 20947 7939
rect 22661 7905 22695 7939
rect 29929 7905 29963 7939
rect 31217 7905 31251 7939
rect 32505 7905 32539 7939
rect 33425 7905 33459 7939
rect 49157 7905 49191 7939
rect 1593 7837 1627 7871
rect 2329 7837 2363 7871
rect 15577 7837 15611 7871
rect 17049 7837 17083 7871
rect 18153 7837 18187 7871
rect 21189 7837 21223 7871
rect 22385 7837 22419 7871
rect 31309 7837 31343 7871
rect 32689 7837 32723 7871
rect 38761 7837 38795 7871
rect 39221 7837 39255 7871
rect 47961 7837 47995 7871
rect 18245 7769 18279 7803
rect 30481 7769 30515 7803
rect 37565 7769 37599 7803
rect 38025 7769 38059 7803
rect 38945 7769 38979 7803
rect 1777 7701 1811 7735
rect 17417 7701 17451 7735
rect 18613 7701 18647 7735
rect 21465 7701 21499 7735
rect 21649 7701 21683 7735
rect 22477 7701 22511 7735
rect 23029 7701 23063 7735
rect 30665 7701 30699 7735
rect 31401 7701 31435 7735
rect 32597 7701 32631 7735
rect 38117 7701 38151 7735
rect 18337 7497 18371 7531
rect 18797 7497 18831 7531
rect 19073 7497 19107 7531
rect 22017 7497 22051 7531
rect 22477 7497 22511 7531
rect 23029 7497 23063 7531
rect 31125 7497 31159 7531
rect 32321 7497 32355 7531
rect 31953 7429 31987 7463
rect 37381 7429 37415 7463
rect 37841 7429 37875 7463
rect 44925 7429 44959 7463
rect 49157 7429 49191 7463
rect 1593 7361 1627 7395
rect 2145 7361 2179 7395
rect 22385 7361 22419 7395
rect 38577 7361 38611 7395
rect 39037 7361 39071 7395
rect 47961 7361 47995 7395
rect 22569 7293 22603 7327
rect 1777 7225 1811 7259
rect 32781 7225 32815 7259
rect 38761 7225 38795 7259
rect 45109 7225 45143 7259
rect 21189 7157 21223 7191
rect 21373 7157 21407 7191
rect 21557 7157 21591 7191
rect 37933 7157 37967 7191
rect 21833 6817 21867 6851
rect 49157 6817 49191 6851
rect 2329 6749 2363 6783
rect 2789 6749 2823 6783
rect 17693 6749 17727 6783
rect 19625 6749 19659 6783
rect 46121 6749 46155 6783
rect 47961 6749 47995 6783
rect 1685 6681 1719 6715
rect 47317 6681 47351 6715
rect 1777 6613 1811 6647
rect 2513 6613 2547 6647
rect 17877 6613 17911 6647
rect 19809 6613 19843 6647
rect 2145 6409 2179 6443
rect 44005 6341 44039 6375
rect 49157 6341 49191 6375
rect 1593 6273 1627 6307
rect 37565 6273 37599 6307
rect 38025 6273 38059 6307
rect 47961 6273 47995 6307
rect 2329 6205 2363 6239
rect 18061 6205 18095 6239
rect 18245 6205 18279 6239
rect 1777 6137 1811 6171
rect 44189 6137 44223 6171
rect 18705 6069 18739 6103
rect 37657 6069 37691 6103
rect 2513 5865 2547 5899
rect 3065 5729 3099 5763
rect 49157 5729 49191 5763
rect 1593 5661 1627 5695
rect 2329 5661 2363 5695
rect 2881 5661 2915 5695
rect 43729 5661 43763 5695
rect 47961 5661 47995 5695
rect 43913 5593 43947 5627
rect 1777 5525 1811 5559
rect 37289 5321 37323 5355
rect 37749 5253 37783 5287
rect 38485 5253 38519 5287
rect 38945 5253 38979 5287
rect 49157 5253 49191 5287
rect 2145 5185 2179 5219
rect 18889 5185 18923 5219
rect 45845 5185 45879 5219
rect 47961 5185 47995 5219
rect 2421 5117 2455 5151
rect 19073 5117 19107 5151
rect 46857 5117 46891 5151
rect 38669 5049 38703 5083
rect 19533 4981 19567 5015
rect 37841 4981 37875 5015
rect 2145 4777 2179 4811
rect 36829 4777 36863 4811
rect 1777 4709 1811 4743
rect 22569 4709 22603 4743
rect 46489 4709 46523 4743
rect 20453 4641 20487 4675
rect 21925 4641 21959 4675
rect 26801 4641 26835 4675
rect 47225 4641 47259 4675
rect 49157 4641 49191 4675
rect 1593 4573 1627 4607
rect 2329 4573 2363 4607
rect 20637 4573 20671 4607
rect 22109 4573 22143 4607
rect 23096 4573 23130 4607
rect 26985 4573 27019 4607
rect 37289 4573 37323 4607
rect 38025 4573 38059 4607
rect 38485 4573 38519 4607
rect 47961 4573 47995 4607
rect 25145 4505 25179 4539
rect 38209 4505 38243 4539
rect 46673 4505 46707 4539
rect 47409 4505 47443 4539
rect 21097 4437 21131 4471
rect 23167 4437 23201 4471
rect 37381 4437 37415 4471
rect 46213 4437 46247 4471
rect 1685 4165 1719 4199
rect 25881 4165 25915 4199
rect 2329 4097 2363 4131
rect 3065 4097 3099 4131
rect 22360 4096 22394 4130
rect 22972 4097 23006 4131
rect 23075 4097 23109 4131
rect 23616 4097 23650 4131
rect 26065 4097 26099 4131
rect 45845 4097 45879 4131
rect 47961 4097 47995 4131
rect 49157 4097 49191 4131
rect 2881 4029 2915 4063
rect 24869 4029 24903 4063
rect 27169 4029 27203 4063
rect 28825 4029 28859 4063
rect 29009 4029 29043 4063
rect 46673 4029 46707 4063
rect 2513 3961 2547 3995
rect 23719 3961 23753 3995
rect 1777 3893 1811 3927
rect 22431 3893 22465 3927
rect 47685 3893 47719 3927
rect 23029 3689 23063 3723
rect 23581 3689 23615 3723
rect 23949 3689 23983 3723
rect 45385 3621 45419 3655
rect 2145 3553 2179 3587
rect 26249 3553 26283 3587
rect 36645 3553 36679 3587
rect 49157 3553 49191 3587
rect 2421 3485 2455 3519
rect 9689 3485 9723 3519
rect 16589 3485 16623 3519
rect 21005 3485 21039 3519
rect 23305 3485 23339 3519
rect 24041 3485 24075 3519
rect 24593 3485 24627 3519
rect 26433 3485 26467 3519
rect 46121 3485 46155 3519
rect 47961 3485 47995 3519
rect 16405 3417 16439 3451
rect 21281 3417 21315 3451
rect 36461 3417 36495 3451
rect 36921 3417 36955 3451
rect 45109 3417 45143 3451
rect 45569 3417 45603 3451
rect 47317 3417 47351 3451
rect 10333 3349 10367 3383
rect 22753 3349 22787 3383
rect 2145 3145 2179 3179
rect 10333 3145 10367 3179
rect 16313 3145 16347 3179
rect 19993 3145 20027 3179
rect 21465 3145 21499 3179
rect 28365 3145 28399 3179
rect 16773 3077 16807 3111
rect 49157 3077 49191 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 9413 3009 9447 3043
rect 9689 3009 9723 3043
rect 12357 3009 12391 3043
rect 14565 3009 14599 3043
rect 17601 3009 17635 3043
rect 19533 3009 19567 3043
rect 20177 3009 20211 3043
rect 20637 3009 20671 3043
rect 21281 3009 21315 3043
rect 22661 3009 22695 3043
rect 23029 3009 23063 3043
rect 23765 3009 23799 3043
rect 26433 3009 26467 3043
rect 27997 3009 28031 3043
rect 28917 3009 28951 3043
rect 44005 3009 44039 3043
rect 45845 3009 45879 3043
rect 47961 3009 47995 3043
rect 13001 2941 13035 2975
rect 14841 2941 14875 2975
rect 18337 2941 18371 2975
rect 24225 2941 24259 2975
rect 24501 2941 24535 2975
rect 25973 2941 26007 2975
rect 29193 2941 29227 2975
rect 31033 2941 31067 2975
rect 45201 2941 45235 2975
rect 46857 2941 46891 2975
rect 1777 2873 1811 2907
rect 20821 2873 20855 2907
rect 22201 2873 22235 2907
rect 27537 2873 27571 2907
rect 2329 2805 2363 2839
rect 2789 2805 2823 2839
rect 17417 2805 17451 2839
rect 22385 2805 22419 2839
rect 23305 2805 23339 2839
rect 23489 2805 23523 2839
rect 26617 2805 26651 2839
rect 27905 2805 27939 2839
rect 30665 2805 30699 2839
rect 2513 2601 2547 2635
rect 24041 2601 24075 2635
rect 26341 2601 26375 2635
rect 29009 2601 29043 2635
rect 35081 2601 35115 2635
rect 1777 2533 1811 2567
rect 3249 2533 3283 2567
rect 9597 2533 9631 2567
rect 30849 2533 30883 2567
rect 32965 2533 32999 2567
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 25053 2465 25087 2499
rect 27629 2465 27663 2499
rect 37749 2465 37783 2499
rect 41429 2465 41463 2499
rect 43821 2465 43855 2499
rect 49157 2465 49191 2499
rect 1593 2397 1627 2431
rect 3065 2397 3099 2431
rect 3525 2397 3559 2431
rect 9413 2397 9447 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 13185 2397 13219 2431
rect 15669 2397 15703 2431
rect 18245 2397 18279 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 22385 2397 22419 2431
rect 24593 2397 24627 2431
rect 27169 2397 27203 2431
rect 29193 2397 29227 2431
rect 29561 2397 29595 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33149 2397 33183 2431
rect 33425 2397 33459 2431
rect 35265 2397 35299 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 40693 2397 40727 2431
rect 43545 2397 43579 2431
rect 45845 2397 45879 2431
rect 47961 2397 47995 2431
rect 2421 2329 2455 2363
rect 11989 2329 12023 2363
rect 14473 2329 14507 2363
rect 17049 2329 17083 2363
rect 47041 2329 47075 2363
rect 18705 2261 18739 2295
rect 19625 2261 19659 2295
rect 37105 2261 37139 2295
rect 43269 2261 43303 2295
<< metal1 >>
rect 3142 25440 3148 25492
rect 3200 25480 3206 25492
rect 9766 25480 9772 25492
rect 3200 25452 9772 25480
rect 3200 25440 3206 25452
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 39574 24964 39580 25016
rect 39632 25004 39638 25016
rect 45738 25004 45744 25016
rect 39632 24976 45744 25004
rect 39632 24964 39638 24976
rect 45738 24964 45744 24976
rect 45796 24964 45802 25016
rect 21542 24896 21548 24948
rect 21600 24936 21606 24948
rect 25958 24936 25964 24948
rect 21600 24908 25964 24936
rect 21600 24896 21606 24908
rect 25958 24896 25964 24908
rect 26016 24896 26022 24948
rect 26050 24896 26056 24948
rect 26108 24936 26114 24948
rect 40954 24936 40960 24948
rect 26108 24908 40960 24936
rect 26108 24896 26114 24908
rect 40954 24896 40960 24908
rect 41012 24896 41018 24948
rect 25866 24828 25872 24880
rect 25924 24868 25930 24880
rect 40402 24868 40408 24880
rect 25924 24840 40408 24868
rect 25924 24828 25930 24840
rect 40402 24828 40408 24840
rect 40460 24828 40466 24880
rect 3878 24760 3884 24812
rect 3936 24800 3942 24812
rect 5902 24800 5908 24812
rect 3936 24772 5908 24800
rect 3936 24760 3942 24772
rect 5902 24760 5908 24772
rect 5960 24760 5966 24812
rect 16022 24760 16028 24812
rect 16080 24800 16086 24812
rect 21726 24800 21732 24812
rect 16080 24772 21732 24800
rect 16080 24760 16086 24772
rect 21726 24760 21732 24772
rect 21784 24760 21790 24812
rect 29914 24760 29920 24812
rect 29972 24800 29978 24812
rect 32858 24800 32864 24812
rect 29972 24772 32864 24800
rect 29972 24760 29978 24772
rect 32858 24760 32864 24772
rect 32916 24760 32922 24812
rect 34882 24760 34888 24812
rect 34940 24800 34946 24812
rect 44358 24800 44364 24812
rect 34940 24772 44364 24800
rect 34940 24760 34946 24772
rect 44358 24760 44364 24772
rect 44416 24760 44422 24812
rect 18874 24692 18880 24744
rect 18932 24732 18938 24744
rect 27246 24732 27252 24744
rect 18932 24704 27252 24732
rect 18932 24692 18938 24704
rect 27246 24692 27252 24704
rect 27304 24692 27310 24744
rect 29546 24692 29552 24744
rect 29604 24732 29610 24744
rect 30650 24732 30656 24744
rect 29604 24704 30656 24732
rect 29604 24692 29610 24704
rect 30650 24692 30656 24704
rect 30708 24692 30714 24744
rect 33962 24692 33968 24744
rect 34020 24732 34026 24744
rect 35158 24732 35164 24744
rect 34020 24704 35164 24732
rect 34020 24692 34026 24704
rect 35158 24692 35164 24704
rect 35216 24732 35222 24744
rect 40586 24732 40592 24744
rect 35216 24704 40592 24732
rect 35216 24692 35222 24704
rect 40586 24692 40592 24704
rect 40644 24692 40650 24744
rect 16206 24624 16212 24676
rect 16264 24664 16270 24676
rect 24026 24664 24032 24676
rect 16264 24636 24032 24664
rect 16264 24624 16270 24636
rect 24026 24624 24032 24636
rect 24084 24624 24090 24676
rect 26418 24624 26424 24676
rect 26476 24664 26482 24676
rect 34974 24664 34980 24676
rect 26476 24636 34980 24664
rect 26476 24624 26482 24636
rect 34974 24624 34980 24636
rect 35032 24664 35038 24676
rect 37550 24664 37556 24676
rect 35032 24636 37556 24664
rect 35032 24624 35038 24636
rect 37550 24624 37556 24636
rect 37608 24624 37614 24676
rect 37642 24624 37648 24676
rect 37700 24664 37706 24676
rect 41046 24664 41052 24676
rect 37700 24636 41052 24664
rect 37700 24624 37706 24636
rect 41046 24624 41052 24636
rect 41104 24624 41110 24676
rect 46290 24624 46296 24676
rect 46348 24664 46354 24676
rect 47762 24664 47768 24676
rect 46348 24636 47768 24664
rect 46348 24624 46354 24636
rect 47762 24624 47768 24636
rect 47820 24624 47826 24676
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 21634 24596 21640 24608
rect 17920 24568 21640 24596
rect 17920 24556 17926 24568
rect 21634 24556 21640 24568
rect 21692 24556 21698 24608
rect 21726 24556 21732 24608
rect 21784 24596 21790 24608
rect 24486 24596 24492 24608
rect 21784 24568 24492 24596
rect 21784 24556 21790 24568
rect 24486 24556 24492 24568
rect 24544 24556 24550 24608
rect 24762 24556 24768 24608
rect 24820 24596 24826 24608
rect 30374 24596 30380 24608
rect 24820 24568 30380 24596
rect 24820 24556 24826 24568
rect 30374 24556 30380 24568
rect 30432 24556 30438 24608
rect 30650 24556 30656 24608
rect 30708 24596 30714 24608
rect 31018 24596 31024 24608
rect 30708 24568 31024 24596
rect 30708 24556 30714 24568
rect 31018 24556 31024 24568
rect 31076 24596 31082 24608
rect 32490 24596 32496 24608
rect 31076 24568 32496 24596
rect 31076 24556 31082 24568
rect 32490 24556 32496 24568
rect 32548 24556 32554 24608
rect 33134 24556 33140 24608
rect 33192 24596 33198 24608
rect 39850 24596 39856 24608
rect 33192 24568 39856 24596
rect 33192 24556 33198 24568
rect 39850 24556 39856 24568
rect 39908 24556 39914 24608
rect 40034 24556 40040 24608
rect 40092 24596 40098 24608
rect 44542 24596 44548 24608
rect 40092 24568 44548 24596
rect 40092 24556 40098 24568
rect 44542 24556 44548 24568
rect 44600 24556 44606 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 10042 24392 10048 24404
rect 3988 24364 10048 24392
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 3510 24256 3516 24268
rect 3007 24228 3516 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 3421 24191 3479 24197
rect 3421 24157 3433 24191
rect 3467 24188 3479 24191
rect 3878 24188 3884 24200
rect 3467 24160 3884 24188
rect 3467 24157 3479 24160
rect 3421 24151 3479 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 3988 24197 4016 24364
rect 10042 24352 10048 24364
rect 10100 24352 10106 24404
rect 20714 24392 20720 24404
rect 18340 24364 20720 24392
rect 15562 24324 15568 24336
rect 9324 24296 15568 24324
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6730 24256 6736 24268
rect 5859 24228 6736 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6730 24216 6736 24228
rect 6788 24216 6794 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8662 24256 8668 24268
rect 8251 24228 8668 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 4614 24148 4620 24200
rect 4672 24148 4678 24200
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24157 6607 24191
rect 6549 24151 6607 24157
rect 6564 24120 6592 24151
rect 7098 24148 7104 24200
rect 7156 24188 7162 24200
rect 7377 24191 7435 24197
rect 7377 24188 7389 24191
rect 7156 24160 7389 24188
rect 7156 24148 7162 24160
rect 7377 24157 7389 24160
rect 7423 24188 7435 24191
rect 7466 24188 7472 24200
rect 7423 24160 7472 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 7466 24148 7472 24160
rect 7524 24148 7530 24200
rect 9324 24197 9352 24296
rect 15562 24284 15568 24296
rect 15620 24284 15626 24336
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24256 10747 24259
rect 11790 24256 11796 24268
rect 10735 24228 11796 24256
rect 10735 24225 10747 24228
rect 10689 24219 10747 24225
rect 11790 24216 11796 24228
rect 11848 24216 11854 24268
rect 13265 24259 13323 24265
rect 13265 24225 13277 24259
rect 13311 24256 13323 24259
rect 13814 24256 13820 24268
rect 13311 24228 13820 24256
rect 13311 24225 13323 24228
rect 13265 24219 13323 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 15841 24259 15899 24265
rect 15841 24225 15853 24259
rect 15887 24256 15899 24259
rect 17678 24256 17684 24268
rect 15887 24228 17684 24256
rect 15887 24225 15899 24228
rect 15841 24219 15899 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24157 11207 24191
rect 11149 24151 11207 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 13725 24191 13783 24197
rect 11931 24160 13676 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 9490 24120 9496 24132
rect 6564 24092 9496 24120
rect 9490 24080 9496 24092
rect 9548 24080 9554 24132
rect 11164 24120 11192 24151
rect 12618 24120 12624 24132
rect 11164 24092 12624 24120
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 13648 24120 13676 24160
rect 13725 24157 13737 24191
rect 13771 24188 13783 24191
rect 14274 24188 14280 24200
rect 13771 24160 14280 24188
rect 13771 24157 13783 24160
rect 13725 24151 13783 24157
rect 14274 24148 14280 24160
rect 14332 24148 14338 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24188 16359 24191
rect 18340 24188 18368 24364
rect 20714 24352 20720 24364
rect 20772 24352 20778 24404
rect 22554 24352 22560 24404
rect 22612 24392 22618 24404
rect 26326 24392 26332 24404
rect 22612 24364 26332 24392
rect 22612 24352 22618 24364
rect 26326 24352 26332 24364
rect 26384 24352 26390 24404
rect 26418 24352 26424 24404
rect 26476 24352 26482 24404
rect 27246 24352 27252 24404
rect 27304 24352 27310 24404
rect 29733 24395 29791 24401
rect 29733 24392 29745 24395
rect 27356 24364 29745 24392
rect 19628 24296 25728 24324
rect 18417 24259 18475 24265
rect 18417 24225 18429 24259
rect 18463 24256 18475 24259
rect 19518 24256 19524 24268
rect 18463 24228 19524 24256
rect 18463 24225 18475 24228
rect 18417 24219 18475 24225
rect 19518 24216 19524 24228
rect 19576 24216 19582 24268
rect 16347 24160 18368 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 18874 24148 18880 24200
rect 18932 24148 18938 24200
rect 19628 24197 19656 24296
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 20990 24216 20996 24268
rect 21048 24256 21054 24268
rect 22186 24256 22192 24268
rect 21048 24228 22192 24256
rect 21048 24216 21054 24228
rect 22186 24216 22192 24228
rect 22244 24216 22250 24268
rect 22462 24216 22468 24268
rect 22520 24216 22526 24268
rect 25133 24259 25191 24265
rect 25133 24256 25145 24259
rect 23584 24228 25145 24256
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 14918 24120 14924 24132
rect 13648 24092 14924 24120
rect 14918 24080 14924 24092
rect 14976 24080 14982 24132
rect 18690 24080 18696 24132
rect 18748 24120 18754 24132
rect 21376 24120 21404 24151
rect 21450 24148 21456 24200
rect 21508 24188 21514 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21508 24160 22017 24188
rect 21508 24148 21514 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 22646 24120 22652 24132
rect 18748 24092 19656 24120
rect 21376 24092 22652 24120
rect 18748 24080 18754 24092
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24052 4215 24055
rect 6638 24052 6644 24064
rect 4203 24024 6644 24052
rect 4203 24021 4215 24024
rect 4157 24015 4215 24021
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 6733 24055 6791 24061
rect 6733 24021 6745 24055
rect 6779 24052 6791 24055
rect 7466 24052 7472 24064
rect 6779 24024 7472 24052
rect 6779 24021 6791 24024
rect 6733 24015 6791 24021
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 11146 24012 11152 24064
rect 11204 24052 11210 24064
rect 11701 24055 11759 24061
rect 11701 24052 11713 24055
rect 11204 24024 11713 24052
rect 11204 24012 11210 24024
rect 11701 24021 11713 24024
rect 11747 24021 11759 24055
rect 11701 24015 11759 24021
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 11848 24024 14289 24052
rect 11848 24012 11854 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 17037 24055 17095 24061
rect 17037 24021 17049 24055
rect 17083 24052 17095 24055
rect 18598 24052 18604 24064
rect 17083 24024 18604 24052
rect 17083 24021 17095 24024
rect 17037 24015 17095 24021
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 19628 24052 19656 24092
rect 22646 24080 22652 24092
rect 22704 24080 22710 24132
rect 23584 24052 23612 24228
rect 25133 24225 25145 24228
rect 25179 24225 25191 24259
rect 25700 24256 25728 24296
rect 25774 24284 25780 24336
rect 25832 24284 25838 24336
rect 27356 24324 27384 24364
rect 29733 24361 29745 24364
rect 29779 24361 29791 24395
rect 29733 24355 29791 24361
rect 33042 24352 33048 24404
rect 33100 24392 33106 24404
rect 33100 24364 33272 24392
rect 33100 24352 33106 24364
rect 25884 24296 27384 24324
rect 25884 24256 25912 24296
rect 28626 24284 28632 24336
rect 28684 24324 28690 24336
rect 31205 24327 31263 24333
rect 28684 24296 30972 24324
rect 28684 24284 28690 24296
rect 26418 24256 26424 24268
rect 25700 24228 25912 24256
rect 25976 24228 26424 24256
rect 25133 24219 25191 24225
rect 23845 24191 23903 24197
rect 23845 24157 23857 24191
rect 23891 24188 23903 24191
rect 25222 24188 25228 24200
rect 23891 24160 25228 24188
rect 23891 24157 23903 24160
rect 23845 24151 23903 24157
rect 25222 24148 25228 24160
rect 25280 24148 25286 24200
rect 25976 24197 26004 24228
rect 26418 24216 26424 24228
rect 26476 24216 26482 24268
rect 27338 24216 27344 24268
rect 27396 24256 27402 24268
rect 29181 24259 29239 24265
rect 29181 24256 29193 24259
rect 27396 24228 29193 24256
rect 27396 24216 27402 24228
rect 25961 24191 26019 24197
rect 25961 24157 25973 24191
rect 26007 24157 26019 24191
rect 25961 24151 26019 24157
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 28552 24197 28580 24228
rect 29181 24225 29193 24228
rect 29227 24225 29239 24259
rect 29181 24219 29239 24225
rect 30944 24256 30972 24296
rect 31205 24293 31217 24327
rect 31251 24324 31263 24327
rect 31570 24324 31576 24336
rect 31251 24296 31576 24324
rect 31251 24293 31263 24296
rect 31205 24287 31263 24293
rect 31570 24284 31576 24296
rect 31628 24284 31634 24336
rect 33244 24324 33272 24364
rect 34606 24352 34612 24404
rect 34664 24392 34670 24404
rect 39482 24392 39488 24404
rect 34664 24364 39488 24392
rect 34664 24352 34670 24364
rect 39482 24352 39488 24364
rect 39540 24352 39546 24404
rect 41046 24352 41052 24404
rect 41104 24352 41110 24404
rect 42518 24352 42524 24404
rect 42576 24392 42582 24404
rect 47857 24395 47915 24401
rect 47857 24392 47869 24395
rect 42576 24364 47869 24392
rect 42576 24352 42582 24364
rect 47857 24361 47869 24364
rect 47903 24361 47915 24395
rect 47857 24355 47915 24361
rect 36446 24324 36452 24336
rect 33244 24296 36452 24324
rect 36446 24284 36452 24296
rect 36504 24284 36510 24336
rect 38197 24327 38255 24333
rect 36556 24296 38148 24324
rect 30944 24228 31616 24256
rect 27893 24191 27951 24197
rect 27893 24188 27905 24191
rect 26292 24160 27905 24188
rect 26292 24148 26298 24160
rect 27893 24157 27905 24160
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 24486 24080 24492 24132
rect 24544 24120 24550 24132
rect 24949 24123 25007 24129
rect 24544 24092 24624 24120
rect 24544 24080 24550 24092
rect 19628 24024 23612 24052
rect 24029 24055 24087 24061
rect 24029 24021 24041 24055
rect 24075 24052 24087 24055
rect 24394 24052 24400 24064
rect 24075 24024 24400 24052
rect 24075 24021 24087 24024
rect 24029 24015 24087 24021
rect 24394 24012 24400 24024
rect 24452 24012 24458 24064
rect 24596 24061 24624 24092
rect 24949 24089 24961 24123
rect 24995 24120 25007 24123
rect 25314 24120 25320 24132
rect 24995 24092 25320 24120
rect 24995 24089 25007 24092
rect 24949 24083 25007 24089
rect 25314 24080 25320 24092
rect 25372 24080 25378 24132
rect 26602 24120 26608 24132
rect 26252 24092 26608 24120
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 26252 24052 26280 24092
rect 26602 24080 26608 24092
rect 26660 24080 26666 24132
rect 26789 24123 26847 24129
rect 26789 24089 26801 24123
rect 26835 24120 26847 24123
rect 27246 24120 27252 24132
rect 26835 24092 27252 24120
rect 26835 24089 26847 24092
rect 26789 24083 26847 24089
rect 27246 24080 27252 24092
rect 27304 24080 27310 24132
rect 27338 24080 27344 24132
rect 27396 24080 27402 24132
rect 27908 24120 27936 24151
rect 29914 24148 29920 24200
rect 29972 24148 29978 24200
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 30944 24188 30972 24228
rect 31021 24191 31079 24197
rect 31021 24188 31033 24191
rect 30432 24160 30696 24188
rect 30944 24160 31033 24188
rect 30432 24148 30438 24160
rect 28997 24123 29055 24129
rect 28997 24120 29009 24123
rect 27908 24092 29009 24120
rect 28997 24089 29009 24092
rect 29043 24089 29055 24123
rect 28997 24083 29055 24089
rect 25087 24024 26280 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 26970 24012 26976 24064
rect 27028 24052 27034 24064
rect 27798 24052 27804 24064
rect 27028 24024 27804 24052
rect 27028 24012 27034 24024
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 28077 24055 28135 24061
rect 28077 24021 28089 24055
rect 28123 24052 28135 24055
rect 28534 24052 28540 24064
rect 28123 24024 28540 24052
rect 28123 24021 28135 24024
rect 28077 24015 28135 24021
rect 28534 24012 28540 24024
rect 28592 24012 28598 24064
rect 28626 24012 28632 24064
rect 28684 24052 28690 24064
rect 28721 24055 28779 24061
rect 28721 24052 28733 24055
rect 28684 24024 28733 24052
rect 28684 24012 28690 24024
rect 28721 24021 28733 24024
rect 28767 24021 28779 24055
rect 28721 24015 28779 24021
rect 30558 24012 30564 24064
rect 30616 24012 30622 24064
rect 30668 24052 30696 24160
rect 31021 24157 31033 24160
rect 31067 24157 31079 24191
rect 31021 24151 31079 24157
rect 31481 24055 31539 24061
rect 31481 24052 31493 24055
rect 30668 24024 31493 24052
rect 31481 24021 31493 24024
rect 31527 24021 31539 24055
rect 31588 24052 31616 24228
rect 34238 24216 34244 24268
rect 34296 24216 34302 24268
rect 35069 24259 35127 24265
rect 35069 24225 35081 24259
rect 35115 24256 35127 24259
rect 35158 24256 35164 24268
rect 35115 24228 35164 24256
rect 35115 24225 35127 24228
rect 35069 24219 35127 24225
rect 35158 24216 35164 24228
rect 35216 24216 35222 24268
rect 36556 24265 36584 24296
rect 36541 24259 36599 24265
rect 36541 24225 36553 24259
rect 36587 24225 36599 24259
rect 36541 24219 36599 24225
rect 36725 24259 36783 24265
rect 36725 24225 36737 24259
rect 36771 24256 36783 24259
rect 37182 24256 37188 24268
rect 36771 24228 37188 24256
rect 36771 24225 36783 24228
rect 36725 24219 36783 24225
rect 37182 24216 37188 24228
rect 37240 24216 37246 24268
rect 37366 24216 37372 24268
rect 37424 24256 37430 24268
rect 37553 24259 37611 24265
rect 37553 24256 37565 24259
rect 37424 24228 37565 24256
rect 37424 24216 37430 24228
rect 37553 24225 37565 24228
rect 37599 24225 37611 24259
rect 38120 24256 38148 24296
rect 38197 24293 38209 24327
rect 38243 24324 38255 24327
rect 39666 24324 39672 24336
rect 38243 24296 39672 24324
rect 38243 24293 38255 24296
rect 38197 24287 38255 24293
rect 39666 24284 39672 24296
rect 39724 24284 39730 24336
rect 43916 24296 45232 24324
rect 40310 24256 40316 24268
rect 38120 24228 40316 24256
rect 37553 24219 37611 24225
rect 40310 24216 40316 24228
rect 40368 24216 40374 24268
rect 40586 24216 40592 24268
rect 40644 24216 40650 24268
rect 41417 24259 41475 24265
rect 41417 24225 41429 24259
rect 41463 24256 41475 24259
rect 43916 24256 43944 24296
rect 41463 24228 43944 24256
rect 41463 24225 41475 24228
rect 41417 24219 41475 24225
rect 32490 24148 32496 24200
rect 32548 24148 32554 24200
rect 32858 24148 32864 24200
rect 32916 24188 32922 24200
rect 33137 24191 33195 24197
rect 33137 24188 33149 24191
rect 32916 24160 33149 24188
rect 32916 24148 32922 24160
rect 33137 24157 33149 24160
rect 33183 24188 33195 24191
rect 33870 24188 33876 24200
rect 33183 24160 33876 24188
rect 33183 24157 33195 24160
rect 33137 24151 33195 24157
rect 33870 24148 33876 24160
rect 33928 24148 33934 24200
rect 34057 24191 34115 24197
rect 34057 24157 34069 24191
rect 34103 24188 34115 24191
rect 34103 24160 38792 24188
rect 34103 24157 34115 24160
rect 34057 24151 34115 24157
rect 33965 24123 34023 24129
rect 33965 24089 33977 24123
rect 34011 24120 34023 24123
rect 35526 24120 35532 24132
rect 34011 24092 35532 24120
rect 34011 24089 34023 24092
rect 33965 24083 34023 24089
rect 35526 24080 35532 24092
rect 35584 24080 35590 24132
rect 36449 24123 36507 24129
rect 36449 24089 36461 24123
rect 36495 24120 36507 24123
rect 36814 24120 36820 24132
rect 36495 24092 36820 24120
rect 36495 24089 36507 24092
rect 36449 24083 36507 24089
rect 36814 24080 36820 24092
rect 36872 24080 36878 24132
rect 37642 24080 37648 24132
rect 37700 24120 37706 24132
rect 37829 24123 37887 24129
rect 37829 24120 37841 24123
rect 37700 24092 37841 24120
rect 37700 24080 37706 24092
rect 37829 24089 37841 24092
rect 37875 24089 37887 24123
rect 38764 24120 38792 24160
rect 38838 24148 38844 24200
rect 38896 24148 38902 24200
rect 39390 24148 39396 24200
rect 39448 24188 39454 24200
rect 39485 24191 39543 24197
rect 39485 24188 39497 24191
rect 39448 24160 39497 24188
rect 39448 24148 39454 24160
rect 39485 24157 39497 24160
rect 39531 24157 39543 24191
rect 39485 24151 39543 24157
rect 42061 24191 42119 24197
rect 42061 24157 42073 24191
rect 42107 24188 42119 24191
rect 42613 24191 42671 24197
rect 42613 24188 42625 24191
rect 42107 24160 42625 24188
rect 42107 24157 42119 24160
rect 42061 24151 42119 24157
rect 42613 24157 42625 24160
rect 42659 24157 42671 24191
rect 42613 24151 42671 24157
rect 42794 24148 42800 24200
rect 42852 24188 42858 24200
rect 43257 24191 43315 24197
rect 43257 24188 43269 24191
rect 42852 24160 43269 24188
rect 42852 24148 42858 24160
rect 43257 24157 43269 24160
rect 43303 24188 43315 24191
rect 43346 24188 43352 24200
rect 43303 24160 43352 24188
rect 43303 24157 43315 24160
rect 43257 24151 43315 24157
rect 43346 24148 43352 24160
rect 43404 24148 43410 24200
rect 43901 24191 43959 24197
rect 43901 24157 43913 24191
rect 43947 24157 43959 24191
rect 43901 24151 43959 24157
rect 40126 24120 40132 24132
rect 38764 24092 40132 24120
rect 37829 24083 37887 24089
rect 40126 24080 40132 24092
rect 40184 24080 40190 24132
rect 40405 24123 40463 24129
rect 40405 24089 40417 24123
rect 40451 24120 40463 24123
rect 40451 24092 41184 24120
rect 40451 24089 40463 24092
rect 40405 24083 40463 24089
rect 31665 24055 31723 24061
rect 31665 24052 31677 24055
rect 31588 24024 31677 24052
rect 31481 24015 31539 24021
rect 31665 24021 31677 24024
rect 31711 24021 31723 24055
rect 31665 24015 31723 24021
rect 31846 24012 31852 24064
rect 31904 24012 31910 24064
rect 32030 24012 32036 24064
rect 32088 24052 32094 24064
rect 32309 24055 32367 24061
rect 32309 24052 32321 24055
rect 32088 24024 32321 24052
rect 32088 24012 32094 24024
rect 32309 24021 32321 24024
rect 32355 24021 32367 24055
rect 32309 24015 32367 24021
rect 32950 24012 32956 24064
rect 33008 24012 33014 24064
rect 33594 24012 33600 24064
rect 33652 24012 33658 24064
rect 34974 24012 34980 24064
rect 35032 24052 35038 24064
rect 35161 24055 35219 24061
rect 35161 24052 35173 24055
rect 35032 24024 35173 24052
rect 35032 24012 35038 24024
rect 35161 24021 35173 24024
rect 35207 24021 35219 24055
rect 35161 24015 35219 24021
rect 35253 24055 35311 24061
rect 35253 24021 35265 24055
rect 35299 24052 35311 24055
rect 35434 24052 35440 24064
rect 35299 24024 35440 24052
rect 35299 24021 35311 24024
rect 35253 24015 35311 24021
rect 35434 24012 35440 24024
rect 35492 24012 35498 24064
rect 35618 24012 35624 24064
rect 35676 24012 35682 24064
rect 36078 24012 36084 24064
rect 36136 24012 36142 24064
rect 37550 24012 37556 24064
rect 37608 24052 37614 24064
rect 37737 24055 37795 24061
rect 37737 24052 37749 24055
rect 37608 24024 37749 24052
rect 37608 24012 37614 24024
rect 37737 24021 37749 24024
rect 37783 24052 37795 24055
rect 38562 24052 38568 24064
rect 37783 24024 38568 24052
rect 37783 24021 37795 24024
rect 37737 24015 37795 24021
rect 38562 24012 38568 24024
rect 38620 24012 38626 24064
rect 38657 24055 38715 24061
rect 38657 24021 38669 24055
rect 38703 24052 38715 24055
rect 38746 24052 38752 24064
rect 38703 24024 38752 24052
rect 38703 24021 38715 24024
rect 38657 24015 38715 24021
rect 38746 24012 38752 24024
rect 38804 24012 38810 24064
rect 39298 24012 39304 24064
rect 39356 24012 39362 24064
rect 40034 24012 40040 24064
rect 40092 24012 40098 24064
rect 40497 24055 40555 24061
rect 40497 24021 40509 24055
rect 40543 24052 40555 24055
rect 40770 24052 40776 24064
rect 40543 24024 40776 24052
rect 40543 24021 40555 24024
rect 40497 24015 40555 24021
rect 40770 24012 40776 24024
rect 40828 24012 40834 24064
rect 41156 24052 41184 24092
rect 41230 24080 41236 24132
rect 41288 24120 41294 24132
rect 43916 24120 43944 24151
rect 44542 24148 44548 24200
rect 44600 24148 44606 24200
rect 45204 24197 45232 24296
rect 46474 24284 46480 24336
rect 46532 24324 46538 24336
rect 48501 24327 48559 24333
rect 48501 24324 48513 24327
rect 46532 24296 48513 24324
rect 46532 24284 46538 24296
rect 48501 24293 48513 24296
rect 48547 24293 48559 24327
rect 48501 24287 48559 24293
rect 45833 24259 45891 24265
rect 45833 24225 45845 24259
rect 45879 24256 45891 24259
rect 45879 24228 48728 24256
rect 45879 24225 45891 24228
rect 45833 24219 45891 24225
rect 48700 24197 48728 24228
rect 45189 24191 45247 24197
rect 45189 24157 45201 24191
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 47213 24191 47271 24197
rect 47213 24157 47225 24191
rect 47259 24188 47271 24191
rect 48685 24191 48743 24197
rect 47259 24160 48636 24188
rect 47259 24157 47271 24160
rect 47213 24151 47271 24157
rect 47118 24120 47124 24132
rect 41288 24092 47124 24120
rect 41288 24080 41294 24092
rect 47118 24080 47124 24092
rect 47176 24080 47182 24132
rect 47762 24080 47768 24132
rect 47820 24120 47826 24132
rect 47949 24123 48007 24129
rect 47949 24120 47961 24123
rect 47820 24092 47961 24120
rect 47820 24080 47826 24092
rect 47949 24089 47961 24092
rect 47995 24089 48007 24123
rect 48608 24120 48636 24160
rect 48685 24157 48697 24191
rect 48731 24157 48743 24191
rect 48685 24151 48743 24157
rect 49050 24148 49056 24200
rect 49108 24188 49114 24200
rect 49329 24191 49387 24197
rect 49329 24188 49341 24191
rect 49108 24160 49341 24188
rect 49108 24148 49114 24160
rect 49329 24157 49341 24160
rect 49375 24157 49387 24191
rect 49329 24151 49387 24157
rect 48608 24092 49372 24120
rect 47949 24083 48007 24089
rect 49344 24064 49372 24092
rect 43622 24052 43628 24064
rect 41156 24024 43628 24052
rect 43622 24012 43628 24024
rect 43680 24012 43686 24064
rect 43714 24012 43720 24064
rect 43772 24012 43778 24064
rect 44358 24012 44364 24064
rect 44416 24012 44422 24064
rect 46014 24012 46020 24064
rect 46072 24052 46078 24064
rect 46109 24055 46167 24061
rect 46109 24052 46121 24055
rect 46072 24024 46121 24052
rect 46072 24012 46078 24024
rect 46109 24021 46121 24024
rect 46155 24021 46167 24055
rect 46109 24015 46167 24021
rect 46566 24012 46572 24064
rect 46624 24012 46630 24064
rect 49142 24012 49148 24064
rect 49200 24012 49206 24064
rect 49326 24012 49332 24064
rect 49384 24012 49390 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 4614 23848 4620 23860
rect 2363 23820 4620 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 10318 23848 10324 23860
rect 6564 23820 10324 23848
rect 6564 23780 6592 23820
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 16206 23848 16212 23860
rect 12360 23820 16212 23848
rect 11790 23780 11796 23792
rect 2148 23752 6592 23780
rect 9324 23752 11796 23780
rect 2148 23721 2176 23752
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 4062 23672 4068 23724
rect 4120 23672 4126 23724
rect 4706 23672 4712 23724
rect 4764 23672 4770 23724
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 7285 23715 7343 23721
rect 7285 23681 7297 23715
rect 7331 23712 7343 23715
rect 8294 23712 8300 23724
rect 7331 23684 8300 23712
rect 7331 23681 7343 23684
rect 7285 23675 7343 23681
rect 3697 23647 3755 23653
rect 3697 23613 3709 23647
rect 3743 23644 3755 23647
rect 4154 23644 4160 23656
rect 3743 23616 4160 23644
rect 3743 23613 3755 23616
rect 3697 23607 3755 23613
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6840 23644 6868 23675
rect 8294 23672 8300 23684
rect 8352 23672 8358 23724
rect 9324 23721 9352 23752
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 12360 23721 12388 23820
rect 16206 23808 16212 23820
rect 16264 23808 16270 23860
rect 19610 23848 19616 23860
rect 16316 23820 19616 23848
rect 14182 23780 14188 23792
rect 13004 23752 14188 23780
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 12345 23715 12403 23721
rect 12345 23681 12357 23715
rect 12391 23681 12403 23715
rect 12710 23712 12716 23724
rect 12345 23675 12403 23681
rect 12544 23684 12716 23712
rect 8386 23644 8392 23656
rect 6840 23616 8392 23644
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 8849 23647 8907 23653
rect 8849 23613 8861 23647
rect 8895 23644 8907 23647
rect 9214 23644 9220 23656
rect 8895 23616 9220 23644
rect 8895 23613 8907 23616
rect 8849 23607 8907 23613
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 10594 23604 10600 23656
rect 10652 23604 10658 23656
rect 11164 23644 11192 23675
rect 12544 23644 12572 23684
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 11164 23616 12572 23644
rect 12621 23647 12679 23653
rect 12621 23613 12633 23647
rect 12667 23644 12679 23647
rect 13004 23644 13032 23752
rect 14182 23740 14188 23752
rect 14240 23740 14246 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 14366 23780 14372 23792
rect 14323 23752 14372 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 14366 23740 14372 23752
rect 14424 23740 14430 23792
rect 16316 23721 16344 23820
rect 19610 23808 19616 23820
rect 19668 23808 19674 23860
rect 21542 23848 21548 23860
rect 20364 23820 21548 23848
rect 20364 23792 20392 23820
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 21634 23808 21640 23860
rect 21692 23848 21698 23860
rect 23293 23851 23351 23857
rect 23293 23848 23305 23851
rect 21692 23820 23305 23848
rect 21692 23808 21698 23820
rect 23293 23817 23305 23820
rect 23339 23817 23351 23851
rect 28445 23851 28503 23857
rect 28445 23848 28457 23851
rect 23293 23811 23351 23817
rect 23400 23820 28457 23848
rect 18874 23740 18880 23792
rect 18932 23780 18938 23792
rect 20257 23783 20315 23789
rect 18932 23752 19090 23780
rect 18932 23740 18938 23752
rect 20257 23749 20269 23783
rect 20303 23780 20315 23783
rect 20346 23780 20352 23792
rect 20303 23752 20352 23780
rect 20303 23749 20315 23752
rect 20257 23743 20315 23749
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 23400 23780 23428 23820
rect 28445 23817 28457 23820
rect 28491 23817 28503 23851
rect 32309 23851 32367 23857
rect 32309 23848 32321 23851
rect 28445 23811 28503 23817
rect 28644 23820 32321 23848
rect 21468 23752 23428 23780
rect 23661 23783 23719 23789
rect 21269 23739 21327 23745
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23681 16359 23715
rect 16301 23675 16359 23681
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 18279 23684 19104 23712
rect 21269 23705 21281 23739
rect 21315 23736 21327 23739
rect 21468 23736 21496 23752
rect 23661 23749 23673 23783
rect 23707 23780 23719 23783
rect 24302 23780 24308 23792
rect 23707 23752 24308 23780
rect 23707 23749 23719 23752
rect 23661 23743 23719 23749
rect 24302 23740 24308 23752
rect 24360 23740 24366 23792
rect 25774 23740 25780 23792
rect 25832 23740 25838 23792
rect 26329 23783 26387 23789
rect 26329 23749 26341 23783
rect 26375 23780 26387 23783
rect 27614 23780 27620 23792
rect 26375 23752 27620 23780
rect 26375 23749 26387 23752
rect 26329 23743 26387 23749
rect 27614 23740 27620 23752
rect 27672 23740 27678 23792
rect 21315 23708 21496 23736
rect 21315 23705 21327 23708
rect 21269 23699 21327 23705
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 12667 23616 13032 23644
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 3970 23536 3976 23588
rect 4028 23576 4034 23588
rect 5810 23576 5816 23588
rect 4028 23548 5816 23576
rect 4028 23536 4034 23548
rect 5810 23536 5816 23548
rect 5868 23536 5874 23588
rect 7469 23579 7527 23585
rect 7469 23545 7481 23579
rect 7515 23576 7527 23579
rect 13096 23576 13124 23675
rect 15841 23647 15899 23653
rect 15841 23613 15853 23647
rect 15887 23644 15899 23647
rect 16390 23644 16396 23656
rect 15887 23616 16396 23644
rect 15887 23613 15899 23616
rect 15841 23607 15899 23613
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18322 23644 18328 23656
rect 17911 23616 18328 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 7515 23548 13124 23576
rect 7515 23545 7527 23548
rect 7469 23539 7527 23545
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 5718 23508 5724 23520
rect 2832 23480 5724 23508
rect 2832 23468 2838 23480
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 5994 23468 6000 23520
rect 6052 23508 6058 23520
rect 6641 23511 6699 23517
rect 6641 23508 6653 23511
rect 6052 23480 6653 23508
rect 6052 23468 6058 23480
rect 6641 23477 6653 23480
rect 6687 23477 6699 23511
rect 6641 23471 6699 23477
rect 18782 23468 18788 23520
rect 18840 23468 18846 23520
rect 19076 23508 19104 23684
rect 21542 23672 21548 23724
rect 21600 23712 21606 23724
rect 23753 23715 23811 23721
rect 21600 23684 22968 23712
rect 21600 23672 21606 23684
rect 20533 23647 20591 23653
rect 20533 23613 20545 23647
rect 20579 23644 20591 23647
rect 22094 23644 22100 23656
rect 20579 23616 22100 23644
rect 20579 23613 20591 23616
rect 20533 23607 20591 23613
rect 22094 23604 22100 23616
rect 22152 23604 22158 23656
rect 22554 23604 22560 23656
rect 22612 23604 22618 23656
rect 22833 23647 22891 23653
rect 22833 23613 22845 23647
rect 22879 23613 22891 23647
rect 22940 23644 22968 23684
rect 23753 23681 23765 23715
rect 23799 23712 23811 23715
rect 25038 23712 25044 23724
rect 23799 23684 25044 23712
rect 23799 23681 23811 23684
rect 23753 23675 23811 23681
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 23845 23647 23903 23653
rect 23845 23644 23857 23647
rect 22940 23616 23857 23644
rect 22833 23607 22891 23613
rect 23845 23613 23857 23616
rect 23891 23613 23903 23647
rect 23845 23607 23903 23613
rect 22738 23576 22744 23588
rect 20456 23548 22744 23576
rect 20456 23508 20484 23548
rect 22738 23536 22744 23548
rect 22796 23536 22802 23588
rect 19076 23480 20484 23508
rect 20993 23511 21051 23517
rect 20993 23477 21005 23511
rect 21039 23508 21051 23511
rect 21082 23508 21088 23520
rect 21039 23480 21088 23508
rect 21039 23477 21051 23480
rect 20993 23471 21051 23477
rect 21082 23468 21088 23480
rect 21140 23468 21146 23520
rect 21450 23468 21456 23520
rect 21508 23468 21514 23520
rect 22848 23508 22876 23607
rect 24210 23604 24216 23656
rect 24268 23644 24274 23656
rect 24268 23616 26556 23644
rect 24268 23604 24274 23616
rect 24489 23579 24547 23585
rect 24489 23576 24501 23579
rect 24044 23548 24501 23576
rect 23474 23508 23480 23520
rect 22848 23480 23480 23508
rect 23474 23468 23480 23480
rect 23532 23508 23538 23520
rect 24044 23508 24072 23548
rect 24489 23545 24501 23548
rect 24535 23545 24547 23579
rect 26528 23576 26556 23616
rect 26602 23604 26608 23656
rect 26660 23604 26666 23656
rect 27157 23579 27215 23585
rect 27157 23576 27169 23579
rect 26528 23548 27169 23576
rect 24489 23539 24547 23545
rect 27157 23545 27169 23548
rect 27203 23545 27215 23579
rect 27356 23576 27384 23675
rect 27798 23672 27804 23724
rect 27856 23672 27862 23724
rect 28644 23721 28672 23820
rect 32309 23817 32321 23820
rect 32355 23817 32367 23851
rect 32309 23811 32367 23817
rect 32769 23851 32827 23857
rect 32769 23817 32781 23851
rect 32815 23848 32827 23851
rect 37461 23851 37519 23857
rect 37461 23848 37473 23851
rect 32815 23820 37473 23848
rect 32815 23817 32827 23820
rect 32769 23811 32827 23817
rect 37461 23817 37473 23820
rect 37507 23817 37519 23851
rect 37461 23811 37519 23817
rect 37829 23851 37887 23857
rect 37829 23817 37841 23851
rect 37875 23848 37887 23851
rect 40034 23848 40040 23860
rect 37875 23820 40040 23848
rect 37875 23817 37887 23820
rect 37829 23811 37887 23817
rect 40034 23808 40040 23820
rect 40092 23808 40098 23860
rect 41046 23808 41052 23860
rect 41104 23848 41110 23860
rect 42153 23851 42211 23857
rect 42153 23848 42165 23851
rect 41104 23820 42165 23848
rect 41104 23808 41110 23820
rect 42153 23817 42165 23820
rect 42199 23848 42211 23851
rect 46750 23848 46756 23860
rect 42199 23820 46756 23848
rect 42199 23817 42211 23820
rect 42153 23811 42211 23817
rect 46750 23808 46756 23820
rect 46808 23808 46814 23860
rect 47118 23808 47124 23860
rect 47176 23808 47182 23860
rect 47302 23808 47308 23860
rect 47360 23848 47366 23860
rect 47673 23851 47731 23857
rect 47673 23848 47685 23851
rect 47360 23820 47685 23848
rect 47360 23808 47366 23820
rect 47673 23817 47685 23820
rect 47719 23848 47731 23851
rect 48590 23848 48596 23860
rect 47719 23820 48596 23848
rect 47719 23817 47731 23820
rect 47673 23811 47731 23817
rect 48590 23808 48596 23820
rect 48648 23808 48654 23860
rect 49326 23808 49332 23860
rect 49384 23808 49390 23860
rect 31481 23783 31539 23789
rect 31481 23749 31493 23783
rect 31527 23780 31539 23783
rect 32582 23780 32588 23792
rect 31527 23752 32588 23780
rect 31527 23749 31539 23752
rect 31481 23743 31539 23749
rect 32582 23740 32588 23752
rect 32640 23780 32646 23792
rect 33042 23780 33048 23792
rect 32640 23752 33048 23780
rect 32640 23740 32646 23752
rect 33042 23740 33048 23752
rect 33100 23740 33106 23792
rect 35618 23740 35624 23792
rect 35676 23780 35682 23792
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 35676 23752 37933 23780
rect 35676 23740 35682 23752
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 38838 23740 38844 23792
rect 38896 23780 38902 23792
rect 39758 23780 39764 23792
rect 38896 23752 39764 23780
rect 38896 23740 38902 23752
rect 39758 23740 39764 23752
rect 39816 23740 39822 23792
rect 39850 23740 39856 23792
rect 39908 23780 39914 23792
rect 42613 23783 42671 23789
rect 42613 23780 42625 23783
rect 39908 23752 42625 23780
rect 39908 23740 39914 23752
rect 28629 23715 28687 23721
rect 28629 23681 28641 23715
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 29089 23715 29147 23721
rect 29089 23681 29101 23715
rect 29135 23712 29147 23715
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 29135 23684 29561 23712
rect 29135 23681 29147 23684
rect 29089 23675 29147 23681
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 28350 23604 28356 23656
rect 28408 23644 28414 23656
rect 29104 23644 29132 23675
rect 30374 23672 30380 23724
rect 30432 23672 30438 23724
rect 32674 23672 32680 23724
rect 32732 23672 32738 23724
rect 34054 23712 34060 23724
rect 32876 23684 34060 23712
rect 28408 23616 29132 23644
rect 28408 23604 28414 23616
rect 29178 23604 29184 23656
rect 29236 23644 29242 23656
rect 29236 23616 31708 23644
rect 29236 23604 29242 23616
rect 29730 23576 29736 23588
rect 27356 23548 29736 23576
rect 27157 23539 27215 23545
rect 29730 23536 29736 23548
rect 29788 23536 29794 23588
rect 30190 23536 30196 23588
rect 30248 23576 30254 23588
rect 31680 23576 31708 23616
rect 31754 23604 31760 23656
rect 31812 23604 31818 23656
rect 31846 23604 31852 23656
rect 31904 23644 31910 23656
rect 32876 23644 32904 23684
rect 34054 23672 34060 23684
rect 34112 23672 34118 23724
rect 35434 23672 35440 23724
rect 35492 23712 35498 23724
rect 36265 23715 36323 23721
rect 35492 23684 35664 23712
rect 35492 23672 35498 23684
rect 35636 23656 35664 23684
rect 36265 23681 36277 23715
rect 36311 23712 36323 23715
rect 39209 23715 39267 23721
rect 36311 23684 38148 23712
rect 36311 23681 36323 23684
rect 36265 23675 36323 23681
rect 31904 23616 32904 23644
rect 32953 23647 33011 23653
rect 31904 23604 31910 23616
rect 32953 23613 32965 23647
rect 32999 23644 33011 23647
rect 33597 23647 33655 23653
rect 33597 23644 33609 23647
rect 32999 23616 33609 23644
rect 32999 23613 33011 23616
rect 32953 23607 33011 23613
rect 33597 23613 33609 23616
rect 33643 23644 33655 23647
rect 34514 23644 34520 23656
rect 33643 23616 34520 23644
rect 33643 23613 33655 23616
rect 33597 23607 33655 23613
rect 34514 23604 34520 23616
rect 34572 23604 34578 23656
rect 35069 23647 35127 23653
rect 35069 23613 35081 23647
rect 35115 23644 35127 23647
rect 35115 23616 35296 23644
rect 35115 23613 35127 23616
rect 35069 23607 35127 23613
rect 32030 23576 32036 23588
rect 30248 23548 30420 23576
rect 31680 23548 32036 23576
rect 30248 23536 30254 23548
rect 23532 23480 24072 23508
rect 23532 23468 23538 23480
rect 24394 23468 24400 23520
rect 24452 23468 24458 23520
rect 24854 23468 24860 23520
rect 24912 23468 24918 23520
rect 27985 23511 28043 23517
rect 27985 23477 27997 23511
rect 28031 23508 28043 23511
rect 28350 23508 28356 23520
rect 28031 23480 28356 23508
rect 28031 23477 28043 23480
rect 27985 23471 28043 23477
rect 28350 23468 28356 23480
rect 28408 23468 28414 23520
rect 29273 23511 29331 23517
rect 29273 23477 29285 23511
rect 29319 23508 29331 23511
rect 29362 23508 29368 23520
rect 29319 23480 29368 23508
rect 29319 23477 29331 23480
rect 29273 23471 29331 23477
rect 29362 23468 29368 23480
rect 29420 23468 29426 23520
rect 30009 23511 30067 23517
rect 30009 23477 30021 23511
rect 30055 23508 30067 23511
rect 30282 23508 30288 23520
rect 30055 23480 30288 23508
rect 30055 23477 30067 23480
rect 30009 23471 30067 23477
rect 30282 23468 30288 23480
rect 30340 23468 30346 23520
rect 30392 23508 30420 23548
rect 32030 23536 32036 23548
rect 32088 23536 32094 23588
rect 35268 23576 35296 23616
rect 35342 23604 35348 23656
rect 35400 23604 35406 23656
rect 35618 23604 35624 23656
rect 35676 23604 35682 23656
rect 35986 23604 35992 23656
rect 36044 23644 36050 23656
rect 36357 23647 36415 23653
rect 36357 23644 36369 23647
rect 36044 23616 36369 23644
rect 36044 23604 36050 23616
rect 36357 23613 36369 23616
rect 36403 23613 36415 23647
rect 36357 23607 36415 23613
rect 36446 23604 36452 23656
rect 36504 23604 36510 23656
rect 38013 23647 38071 23653
rect 38013 23644 38025 23647
rect 36556 23616 38025 23644
rect 35434 23576 35440 23588
rect 32232 23548 33732 23576
rect 35268 23548 35440 23576
rect 32232 23508 32260 23548
rect 30392 23480 32260 23508
rect 33704 23508 33732 23548
rect 35434 23536 35440 23548
rect 35492 23576 35498 23588
rect 36556 23576 36584 23616
rect 38013 23613 38025 23616
rect 38059 23613 38071 23647
rect 38013 23607 38071 23613
rect 35492 23548 36584 23576
rect 38120 23576 38148 23684
rect 39209 23681 39221 23715
rect 39255 23712 39267 23715
rect 39574 23712 39580 23724
rect 39255 23684 39580 23712
rect 39255 23681 39267 23684
rect 39209 23675 39267 23681
rect 39574 23672 39580 23684
rect 39632 23672 39638 23724
rect 40236 23721 40264 23752
rect 42613 23749 42625 23752
rect 42659 23749 42671 23783
rect 42613 23743 42671 23749
rect 45554 23740 45560 23792
rect 45612 23780 45618 23792
rect 45612 23752 46704 23780
rect 45612 23740 45618 23752
rect 40221 23715 40279 23721
rect 40221 23681 40233 23715
rect 40267 23681 40279 23715
rect 40221 23675 40279 23681
rect 43990 23672 43996 23724
rect 44048 23712 44054 23724
rect 44821 23715 44879 23721
rect 44821 23712 44833 23715
rect 44048 23684 44833 23712
rect 44048 23672 44054 23684
rect 44821 23681 44833 23684
rect 44867 23681 44879 23715
rect 44821 23675 44879 23681
rect 45922 23672 45928 23724
rect 45980 23672 45986 23724
rect 46676 23721 46704 23752
rect 47762 23740 47768 23792
rect 47820 23780 47826 23792
rect 49421 23783 49479 23789
rect 49421 23780 49433 23783
rect 47820 23752 49433 23780
rect 47820 23740 47826 23752
rect 49421 23749 49433 23752
rect 49467 23749 49479 23783
rect 49421 23743 49479 23749
rect 46661 23715 46719 23721
rect 46661 23681 46673 23715
rect 46707 23712 46719 23715
rect 46707 23684 47440 23712
rect 46707 23681 46719 23684
rect 46661 23675 46719 23681
rect 39301 23647 39359 23653
rect 39301 23644 39313 23647
rect 39224 23616 39313 23644
rect 39224 23588 39252 23616
rect 39301 23613 39313 23616
rect 39347 23613 39359 23647
rect 39301 23607 39359 23613
rect 39393 23647 39451 23653
rect 39393 23613 39405 23647
rect 39439 23613 39451 23647
rect 39393 23607 39451 23613
rect 38841 23579 38899 23585
rect 38841 23576 38853 23579
rect 38120 23548 38853 23576
rect 35492 23536 35498 23548
rect 38841 23545 38853 23548
rect 38887 23545 38899 23579
rect 38841 23539 38899 23545
rect 39206 23536 39212 23588
rect 39264 23536 39270 23588
rect 39408 23576 39436 23607
rect 39758 23604 39764 23656
rect 39816 23644 39822 23656
rect 39816 23616 40172 23644
rect 39816 23604 39822 23616
rect 39316 23548 39436 23576
rect 35897 23511 35955 23517
rect 35897 23508 35909 23511
rect 33704 23480 35909 23508
rect 35897 23477 35909 23480
rect 35943 23477 35955 23511
rect 35897 23471 35955 23477
rect 36262 23468 36268 23520
rect 36320 23508 36326 23520
rect 36909 23511 36967 23517
rect 36909 23508 36921 23511
rect 36320 23480 36921 23508
rect 36320 23468 36326 23480
rect 36909 23477 36921 23480
rect 36955 23477 36967 23511
rect 36909 23471 36967 23477
rect 38562 23468 38568 23520
rect 38620 23468 38626 23520
rect 39114 23468 39120 23520
rect 39172 23508 39178 23520
rect 39316 23508 39344 23548
rect 39482 23536 39488 23588
rect 39540 23576 39546 23588
rect 40037 23579 40095 23585
rect 40037 23576 40049 23579
rect 39540 23548 40049 23576
rect 39540 23536 39546 23548
rect 40037 23545 40049 23548
rect 40083 23545 40095 23579
rect 40144 23576 40172 23616
rect 40678 23604 40684 23656
rect 40736 23604 40742 23656
rect 40954 23604 40960 23656
rect 41012 23604 41018 23656
rect 42794 23604 42800 23656
rect 42852 23644 42858 23656
rect 43073 23647 43131 23653
rect 43073 23644 43085 23647
rect 42852 23616 43085 23644
rect 42852 23604 42858 23616
rect 43073 23613 43085 23616
rect 43119 23613 43131 23647
rect 43073 23607 43131 23613
rect 44542 23604 44548 23656
rect 44600 23644 44606 23656
rect 47305 23647 47363 23653
rect 47305 23644 47317 23647
rect 44600 23616 47317 23644
rect 44600 23604 44606 23616
rect 47305 23613 47317 23616
rect 47351 23613 47363 23647
rect 47412 23644 47440 23684
rect 48774 23672 48780 23724
rect 48832 23672 48838 23724
rect 49053 23647 49111 23653
rect 49053 23644 49065 23647
rect 47412 23616 49065 23644
rect 47305 23607 47363 23613
rect 49053 23613 49065 23616
rect 49099 23613 49111 23647
rect 49053 23607 49111 23613
rect 41785 23579 41843 23585
rect 41785 23576 41797 23579
rect 40144 23548 41797 23576
rect 40037 23539 40095 23545
rect 41785 23545 41797 23548
rect 41831 23545 41843 23579
rect 41785 23539 41843 23545
rect 42058 23536 42064 23588
rect 42116 23576 42122 23588
rect 46937 23579 46995 23585
rect 46937 23576 46949 23579
rect 42116 23548 46949 23576
rect 42116 23536 42122 23548
rect 46937 23545 46949 23548
rect 46983 23545 46995 23579
rect 46937 23539 46995 23545
rect 47394 23536 47400 23588
rect 47452 23576 47458 23588
rect 48133 23579 48191 23585
rect 48133 23576 48145 23579
rect 47452 23548 48145 23576
rect 47452 23536 47458 23548
rect 48133 23545 48145 23548
rect 48179 23545 48191 23579
rect 48133 23539 48191 23545
rect 39172 23480 39344 23508
rect 39172 23468 39178 23480
rect 39390 23468 39396 23520
rect 39448 23508 39454 23520
rect 41969 23511 42027 23517
rect 41969 23508 41981 23511
rect 39448 23480 41981 23508
rect 39448 23468 39454 23480
rect 41969 23477 41981 23480
rect 42015 23477 42027 23511
rect 41969 23471 42027 23477
rect 42426 23468 42432 23520
rect 42484 23468 42490 23520
rect 43530 23468 43536 23520
rect 43588 23508 43594 23520
rect 45281 23511 45339 23517
rect 45281 23508 45293 23511
rect 43588 23480 45293 23508
rect 43588 23468 43594 23480
rect 45281 23477 45293 23480
rect 45327 23477 45339 23511
rect 45281 23471 45339 23477
rect 46106 23468 46112 23520
rect 46164 23508 46170 23520
rect 46477 23511 46535 23517
rect 46477 23508 46489 23511
rect 46164 23480 46489 23508
rect 46164 23468 46170 23480
rect 46477 23477 46489 23480
rect 46523 23477 46535 23511
rect 46477 23471 46535 23477
rect 47670 23468 47676 23520
rect 47728 23508 47734 23520
rect 47765 23511 47823 23517
rect 47765 23508 47777 23511
rect 47728 23480 47777 23508
rect 47728 23468 47734 23480
rect 47765 23477 47777 23480
rect 47811 23477 47823 23511
rect 47765 23471 47823 23477
rect 47946 23468 47952 23520
rect 48004 23508 48010 23520
rect 49050 23508 49056 23520
rect 48004 23480 49056 23508
rect 48004 23468 48010 23480
rect 49050 23468 49056 23480
rect 49108 23468 49114 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 4706 23264 4712 23316
rect 4764 23264 4770 23316
rect 5626 23304 5632 23316
rect 4816 23276 5632 23304
rect 4816 23168 4844 23276
rect 5626 23264 5632 23276
rect 5684 23264 5690 23316
rect 14182 23264 14188 23316
rect 14240 23304 14246 23316
rect 14240 23276 19196 23304
rect 14240 23264 14246 23276
rect 9214 23236 9220 23248
rect 2976 23140 4844 23168
rect 4908 23208 9220 23236
rect 2976 23109 3004 23140
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4430 23100 4436 23112
rect 4295 23072 4436 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4430 23060 4436 23072
rect 4488 23060 4494 23112
rect 4908 23109 4936 23208
rect 9214 23196 9220 23208
rect 9272 23196 9278 23248
rect 15654 23236 15660 23248
rect 10060 23208 15660 23236
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 10060 23177 10088 23208
rect 15654 23196 15660 23208
rect 15712 23196 15718 23248
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23137 10103 23171
rect 10045 23131 10103 23137
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13354 23168 13360 23180
rect 13311 23140 13360 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 15746 23128 15752 23180
rect 15804 23128 15810 23180
rect 19058 23168 19064 23180
rect 16684 23140 19064 23168
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 1762 22992 1768 23044
rect 1820 22992 1826 23044
rect 3602 22992 3608 23044
rect 3660 23032 3666 23044
rect 5368 23032 5396 23063
rect 6638 23060 6644 23112
rect 6696 23100 6702 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 6696 23072 7205 23100
rect 6696 23060 6702 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 9122 23060 9128 23112
rect 9180 23100 9186 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 9180 23072 9321 23100
rect 9180 23060 9186 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 11882 23060 11888 23112
rect 11940 23060 11946 23112
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 16684 23109 16712 23140
rect 19058 23128 19064 23140
rect 19116 23128 19122 23180
rect 19168 23168 19196 23276
rect 20254 23264 20260 23316
rect 20312 23304 20318 23316
rect 22462 23304 22468 23316
rect 20312 23276 22468 23304
rect 20312 23264 20318 23276
rect 22462 23264 22468 23276
rect 22520 23264 22526 23316
rect 23382 23264 23388 23316
rect 23440 23304 23446 23316
rect 24210 23304 24216 23316
rect 23440 23276 24216 23304
rect 23440 23264 23446 23276
rect 24210 23264 24216 23276
rect 24268 23264 24274 23316
rect 24854 23304 24860 23316
rect 24688 23276 24860 23304
rect 19610 23196 19616 23248
rect 19668 23196 19674 23248
rect 22738 23196 22744 23248
rect 22796 23236 22802 23248
rect 24581 23239 24639 23245
rect 24581 23236 24593 23239
rect 22796 23208 24593 23236
rect 22796 23196 22802 23208
rect 24581 23205 24593 23208
rect 24627 23205 24639 23239
rect 24581 23199 24639 23205
rect 19168 23140 20484 23168
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 3660 23004 5396 23032
rect 14844 23032 14872 23063
rect 17494 23060 17500 23112
rect 17552 23060 17558 23112
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23100 18935 23103
rect 19334 23100 19340 23112
rect 18923 23072 19340 23100
rect 18923 23069 18935 23072
rect 18877 23063 18935 23069
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 18601 23035 18659 23041
rect 14844 23004 17356 23032
rect 3660 22992 3666 23004
rect 4065 22967 4123 22973
rect 4065 22933 4077 22967
rect 4111 22964 4123 22967
rect 4614 22964 4620 22976
rect 4111 22936 4620 22964
rect 4111 22933 4123 22936
rect 4065 22927 4123 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 5350 22924 5356 22976
rect 5408 22964 5414 22976
rect 9217 22967 9275 22973
rect 9217 22964 9229 22967
rect 5408 22936 9229 22964
rect 5408 22924 5414 22936
rect 9217 22933 9229 22936
rect 9263 22933 9275 22967
rect 9217 22927 9275 22933
rect 14090 22924 14096 22976
rect 14148 22964 14154 22976
rect 14277 22967 14335 22973
rect 14277 22964 14289 22967
rect 14148 22936 14289 22964
rect 14148 22924 14154 22936
rect 14277 22933 14289 22936
rect 14323 22933 14335 22967
rect 14277 22927 14335 22933
rect 14642 22924 14648 22976
rect 14700 22924 14706 22976
rect 17126 22924 17132 22976
rect 17184 22924 17190 22976
rect 17328 22964 17356 23004
rect 18601 23001 18613 23035
rect 18647 23032 18659 23035
rect 18690 23032 18696 23044
rect 18647 23004 18696 23032
rect 18647 23001 18659 23004
rect 18601 22995 18659 23001
rect 18690 22992 18696 23004
rect 18748 22992 18754 23044
rect 19794 22992 19800 23044
rect 19852 22992 19858 23044
rect 17770 22964 17776 22976
rect 17328 22936 17776 22964
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 19245 22967 19303 22973
rect 19245 22964 19257 22967
rect 18932 22936 19257 22964
rect 18932 22924 18938 22936
rect 19245 22933 19257 22936
rect 19291 22933 19303 22967
rect 19245 22927 19303 22933
rect 20346 22924 20352 22976
rect 20404 22924 20410 22976
rect 20456 22964 20484 23140
rect 21174 23128 21180 23180
rect 21232 23168 21238 23180
rect 21821 23171 21879 23177
rect 21821 23168 21833 23171
rect 21232 23140 21833 23168
rect 21232 23128 21238 23140
rect 21821 23137 21833 23140
rect 21867 23168 21879 23171
rect 22186 23168 22192 23180
rect 21867 23140 22192 23168
rect 21867 23137 21879 23140
rect 21821 23131 21879 23137
rect 22186 23128 22192 23140
rect 22244 23128 22250 23180
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 24688 23168 24716 23276
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 25038 23264 25044 23316
rect 25096 23304 25102 23316
rect 27893 23307 27951 23313
rect 27893 23304 27905 23307
rect 25096 23276 27905 23304
rect 25096 23264 25102 23276
rect 27893 23273 27905 23276
rect 27939 23273 27951 23307
rect 27893 23267 27951 23273
rect 29730 23264 29736 23316
rect 29788 23264 29794 23316
rect 30834 23264 30840 23316
rect 30892 23304 30898 23316
rect 33226 23304 33232 23316
rect 30892 23276 33232 23304
rect 30892 23264 30898 23276
rect 33226 23264 33232 23276
rect 33284 23264 33290 23316
rect 33870 23264 33876 23316
rect 33928 23304 33934 23316
rect 34149 23307 34207 23313
rect 34149 23304 34161 23307
rect 33928 23276 34161 23304
rect 33928 23264 33934 23276
rect 34149 23273 34161 23276
rect 34195 23273 34207 23307
rect 34149 23267 34207 23273
rect 34238 23264 34244 23316
rect 34296 23304 34302 23316
rect 34296 23276 36400 23304
rect 34296 23264 34302 23276
rect 25222 23196 25228 23248
rect 25280 23196 25286 23248
rect 27798 23196 27804 23248
rect 27856 23236 27862 23248
rect 28997 23239 29055 23245
rect 28997 23236 29009 23239
rect 27856 23208 29009 23236
rect 27856 23196 27862 23208
rect 28997 23205 29009 23208
rect 29043 23205 29055 23239
rect 28997 23199 29055 23205
rect 29365 23239 29423 23245
rect 29365 23205 29377 23239
rect 29411 23236 29423 23239
rect 31294 23236 31300 23248
rect 29411 23208 31300 23236
rect 29411 23205 29423 23208
rect 29365 23199 29423 23205
rect 23983 23140 24716 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 24854 23128 24860 23180
rect 24912 23168 24918 23180
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 24912 23140 25973 23168
rect 24912 23128 24918 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 25961 23131 26019 23137
rect 26694 23128 26700 23180
rect 26752 23168 26758 23180
rect 28445 23171 28503 23177
rect 28445 23168 28457 23171
rect 26752 23140 28457 23168
rect 26752 23128 26758 23140
rect 28445 23137 28457 23140
rect 28491 23137 28503 23171
rect 28445 23131 28503 23137
rect 29181 23171 29239 23177
rect 29181 23137 29193 23171
rect 29227 23168 29239 23171
rect 29270 23168 29276 23180
rect 29227 23140 29276 23168
rect 29227 23137 29239 23140
rect 29181 23131 29239 23137
rect 29270 23128 29276 23140
rect 29328 23128 29334 23180
rect 22094 23060 22100 23112
rect 22152 23060 22158 23112
rect 23750 23060 23756 23112
rect 23808 23060 23814 23112
rect 24762 23060 24768 23112
rect 24820 23060 24826 23112
rect 25682 23060 25688 23112
rect 25740 23060 25746 23112
rect 28353 23103 28411 23109
rect 28353 23069 28365 23103
rect 28399 23100 28411 23103
rect 29380 23100 29408 23199
rect 31294 23196 31300 23208
rect 31352 23196 31358 23248
rect 33137 23239 33195 23245
rect 33137 23205 33149 23239
rect 33183 23236 33195 23239
rect 33962 23236 33968 23248
rect 33183 23208 33968 23236
rect 33183 23205 33195 23208
rect 33137 23199 33195 23205
rect 33962 23196 33968 23208
rect 34020 23196 34026 23248
rect 34054 23196 34060 23248
rect 34112 23236 34118 23248
rect 34425 23239 34483 23245
rect 34425 23236 34437 23239
rect 34112 23208 34437 23236
rect 34112 23196 34118 23208
rect 34425 23205 34437 23208
rect 34471 23205 34483 23239
rect 34425 23199 34483 23205
rect 30190 23128 30196 23180
rect 30248 23128 30254 23180
rect 30282 23128 30288 23180
rect 30340 23128 30346 23180
rect 31018 23128 31024 23180
rect 31076 23128 31082 23180
rect 31754 23168 31760 23180
rect 31404 23140 31760 23168
rect 28399 23072 29408 23100
rect 28399 23069 28411 23072
rect 28353 23063 28411 23069
rect 29454 23060 29460 23112
rect 29512 23100 29518 23112
rect 29512 23072 30236 23100
rect 29512 23060 29518 23072
rect 21082 22992 21088 23044
rect 21140 22992 21146 23044
rect 21910 22992 21916 23044
rect 21968 23032 21974 23044
rect 22557 23035 22615 23041
rect 22557 23032 22569 23035
rect 21968 23004 22569 23032
rect 21968 22992 21974 23004
rect 22557 23001 22569 23004
rect 22603 23001 22615 23035
rect 22557 22995 22615 23001
rect 22741 23035 22799 23041
rect 22741 23001 22753 23035
rect 22787 23032 22799 23035
rect 25130 23032 25136 23044
rect 22787 23004 25136 23032
rect 22787 23001 22799 23004
rect 22741 22995 22799 23001
rect 25130 22992 25136 23004
rect 25188 22992 25194 23044
rect 26234 23032 26240 23044
rect 25240 23004 26240 23032
rect 22830 22964 22836 22976
rect 20456 22936 22836 22964
rect 22830 22924 22836 22936
rect 22888 22924 22894 22976
rect 23290 22924 23296 22976
rect 23348 22924 23354 22976
rect 23661 22967 23719 22973
rect 23661 22933 23673 22967
rect 23707 22964 23719 22967
rect 25240 22964 25268 23004
rect 26234 22992 26240 23004
rect 26292 22992 26298 23044
rect 27246 23032 27252 23044
rect 27186 23004 27252 23032
rect 27246 22992 27252 23004
rect 27304 22992 27310 23044
rect 29914 23032 29920 23044
rect 27448 23004 29920 23032
rect 23707 22936 25268 22964
rect 23707 22933 23719 22936
rect 23661 22927 23719 22933
rect 25314 22924 25320 22976
rect 25372 22924 25378 22976
rect 26326 22924 26332 22976
rect 26384 22964 26390 22976
rect 27448 22973 27476 23004
rect 29914 22992 29920 23004
rect 29972 22992 29978 23044
rect 27433 22967 27491 22973
rect 27433 22964 27445 22967
rect 26384 22936 27445 22964
rect 26384 22924 26390 22936
rect 27433 22933 27445 22936
rect 27479 22933 27491 22967
rect 27433 22927 27491 22933
rect 28261 22967 28319 22973
rect 28261 22933 28273 22967
rect 28307 22964 28319 22967
rect 30006 22964 30012 22976
rect 28307 22936 30012 22964
rect 28307 22933 28319 22936
rect 28261 22927 28319 22933
rect 30006 22924 30012 22936
rect 30064 22924 30070 22976
rect 30098 22924 30104 22976
rect 30156 22924 30162 22976
rect 30208 22964 30236 23072
rect 30300 23032 30328 23128
rect 31404 23112 31432 23140
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 34330 23128 34336 23180
rect 34388 23168 34394 23180
rect 35069 23171 35127 23177
rect 35069 23168 35081 23171
rect 34388 23140 35081 23168
rect 34388 23128 34394 23140
rect 35069 23137 35081 23140
rect 35115 23168 35127 23171
rect 35342 23168 35348 23180
rect 35115 23140 35348 23168
rect 35115 23137 35127 23140
rect 35069 23131 35127 23137
rect 35342 23128 35348 23140
rect 35400 23128 35406 23180
rect 36372 23168 36400 23276
rect 37458 23264 37464 23316
rect 37516 23304 37522 23316
rect 38767 23307 38825 23313
rect 38767 23304 38779 23307
rect 37516 23276 38779 23304
rect 37516 23264 37522 23276
rect 38767 23273 38779 23276
rect 38813 23304 38825 23307
rect 39022 23304 39028 23316
rect 38813 23276 39028 23304
rect 38813 23273 38825 23276
rect 38767 23267 38825 23273
rect 39022 23264 39028 23276
rect 39080 23264 39086 23316
rect 39942 23264 39948 23316
rect 40000 23304 40006 23316
rect 41049 23307 41107 23313
rect 41049 23304 41061 23307
rect 40000 23276 41061 23304
rect 40000 23264 40006 23276
rect 41049 23273 41061 23276
rect 41095 23273 41107 23307
rect 41049 23267 41107 23273
rect 37277 23171 37335 23177
rect 37277 23168 37289 23171
rect 36372 23140 37289 23168
rect 37277 23137 37289 23140
rect 37323 23168 37335 23171
rect 38286 23168 38292 23180
rect 37323 23140 38292 23168
rect 37323 23137 37335 23140
rect 37277 23131 37335 23137
rect 38286 23128 38292 23140
rect 38344 23128 38350 23180
rect 38654 23128 38660 23180
rect 38712 23168 38718 23180
rect 39025 23171 39083 23177
rect 39025 23168 39037 23171
rect 38712 23140 39037 23168
rect 38712 23128 38718 23140
rect 39025 23137 39037 23140
rect 39071 23168 39083 23171
rect 39482 23168 39488 23180
rect 39071 23140 39488 23168
rect 39071 23137 39083 23140
rect 39025 23131 39083 23137
rect 39482 23128 39488 23140
rect 39540 23128 39546 23180
rect 40678 23128 40684 23180
rect 40736 23128 40742 23180
rect 41064 23168 41092 23267
rect 43990 23264 43996 23316
rect 44048 23264 44054 23316
rect 48774 23264 48780 23316
rect 48832 23304 48838 23316
rect 48869 23307 48927 23313
rect 48869 23304 48881 23307
rect 48832 23276 48881 23304
rect 48832 23264 48838 23276
rect 48869 23273 48881 23276
rect 48915 23273 48927 23307
rect 48869 23267 48927 23273
rect 49234 23264 49240 23316
rect 49292 23264 49298 23316
rect 46750 23196 46756 23248
rect 46808 23196 46814 23248
rect 42794 23168 42800 23180
rect 41064 23140 42800 23168
rect 42794 23128 42800 23140
rect 42852 23168 42858 23180
rect 43533 23171 43591 23177
rect 43533 23168 43545 23171
rect 42852 23140 43545 23168
rect 42852 23128 42858 23140
rect 43533 23137 43545 23140
rect 43579 23137 43591 23171
rect 43533 23131 43591 23137
rect 43990 23128 43996 23180
rect 44048 23168 44054 23180
rect 45189 23171 45247 23177
rect 45189 23168 45201 23171
rect 44048 23140 45201 23168
rect 44048 23128 44054 23140
rect 45189 23137 45201 23140
rect 45235 23137 45247 23171
rect 45189 23131 45247 23137
rect 46566 23128 46572 23180
rect 46624 23168 46630 23180
rect 46624 23140 48268 23168
rect 46624 23128 46630 23140
rect 31386 23060 31392 23112
rect 31444 23060 31450 23112
rect 33873 23103 33931 23109
rect 33873 23100 33885 23103
rect 33060 23072 33885 23100
rect 31665 23035 31723 23041
rect 31665 23032 31677 23035
rect 30300 23004 31677 23032
rect 31665 23001 31677 23004
rect 31711 23001 31723 23035
rect 31665 22995 31723 23001
rect 31754 22992 31760 23044
rect 31812 23032 31818 23044
rect 31812 23004 32154 23032
rect 31812 22992 31818 23004
rect 30374 22964 30380 22976
rect 30208 22936 30380 22964
rect 30374 22924 30380 22936
rect 30432 22964 30438 22976
rect 30745 22967 30803 22973
rect 30745 22964 30757 22967
rect 30432 22936 30757 22964
rect 30432 22924 30438 22936
rect 30745 22933 30757 22936
rect 30791 22933 30803 22967
rect 30745 22927 30803 22933
rect 31202 22924 31208 22976
rect 31260 22964 31266 22976
rect 33060 22964 33088 23072
rect 33873 23069 33885 23072
rect 33919 23100 33931 23103
rect 34701 23103 34759 23109
rect 34701 23100 34713 23103
rect 33919 23072 34713 23100
rect 33919 23069 33931 23072
rect 33873 23063 33931 23069
rect 34701 23069 34713 23072
rect 34747 23069 34759 23103
rect 37642 23100 37648 23112
rect 36478 23086 37648 23100
rect 34701 23063 34759 23069
rect 36464 23072 37648 23086
rect 34514 22992 34520 23044
rect 34572 23032 34578 23044
rect 35345 23035 35403 23041
rect 35345 23032 35357 23035
rect 34572 23004 35357 23032
rect 34572 22992 34578 23004
rect 35345 23001 35357 23004
rect 35391 23001 35403 23035
rect 35345 22995 35403 23001
rect 35452 23004 35834 23032
rect 31260 22936 33088 22964
rect 33689 22967 33747 22973
rect 31260 22924 31266 22936
rect 33689 22933 33701 22967
rect 33735 22964 33747 22967
rect 33778 22964 33784 22976
rect 33735 22936 33784 22964
rect 33735 22933 33747 22936
rect 33689 22927 33747 22933
rect 33778 22924 33784 22936
rect 33836 22924 33842 22976
rect 34054 22924 34060 22976
rect 34112 22964 34118 22976
rect 35452 22964 35480 23004
rect 34112 22936 35480 22964
rect 35728 22964 35756 23004
rect 36262 22964 36268 22976
rect 35728 22936 36268 22964
rect 34112 22924 34118 22936
rect 36262 22924 36268 22936
rect 36320 22964 36326 22976
rect 36464 22964 36492 23072
rect 37642 23060 37648 23072
rect 37700 23060 37706 23112
rect 39500 23100 39528 23128
rect 39942 23100 39948 23112
rect 39500 23072 39948 23100
rect 39942 23060 39948 23072
rect 40000 23060 40006 23112
rect 40034 23060 40040 23112
rect 40092 23100 40098 23112
rect 40405 23103 40463 23109
rect 40405 23100 40417 23103
rect 40092 23072 40417 23100
rect 40092 23060 40098 23072
rect 40405 23069 40417 23072
rect 40451 23069 40463 23103
rect 41322 23100 41328 23112
rect 40405 23063 40463 23069
rect 40512 23072 41328 23100
rect 38654 22992 38660 23044
rect 38712 23032 38718 23044
rect 39114 23032 39120 23044
rect 38712 23004 39120 23032
rect 38712 22992 38718 23004
rect 39114 22992 39120 23004
rect 39172 22992 39178 23044
rect 40512 23032 40540 23072
rect 41322 23060 41328 23072
rect 41380 23060 41386 23112
rect 44637 23103 44695 23109
rect 44637 23069 44649 23103
rect 44683 23100 44695 23103
rect 46474 23100 46480 23112
rect 44683 23072 46480 23100
rect 44683 23069 44695 23072
rect 44637 23063 44695 23069
rect 46474 23060 46480 23072
rect 46532 23060 46538 23112
rect 46658 23060 46664 23112
rect 46716 23100 46722 23112
rect 46937 23103 46995 23109
rect 46937 23100 46949 23103
rect 46716 23072 46949 23100
rect 46716 23060 46722 23072
rect 46937 23069 46949 23072
rect 46983 23100 46995 23103
rect 47670 23100 47676 23112
rect 46983 23072 47676 23100
rect 46983 23069 46995 23072
rect 46937 23063 46995 23069
rect 47670 23060 47676 23072
rect 47728 23060 47734 23112
rect 48240 23109 48268 23140
rect 47765 23103 47823 23109
rect 47765 23069 47777 23103
rect 47811 23069 47823 23103
rect 47765 23063 47823 23069
rect 48225 23103 48283 23109
rect 48225 23069 48237 23103
rect 48271 23069 48283 23103
rect 48225 23063 48283 23069
rect 39316 23004 40540 23032
rect 41509 23035 41567 23041
rect 36320 22936 36492 22964
rect 36320 22924 36326 22936
rect 36630 22924 36636 22976
rect 36688 22964 36694 22976
rect 36817 22967 36875 22973
rect 36817 22964 36829 22967
rect 36688 22936 36829 22964
rect 36688 22924 36694 22936
rect 36817 22933 36829 22936
rect 36863 22933 36875 22967
rect 36817 22927 36875 22933
rect 37826 22924 37832 22976
rect 37884 22964 37890 22976
rect 39316 22964 39344 23004
rect 41509 23001 41521 23035
rect 41555 23001 41567 23035
rect 41509 22995 41567 23001
rect 37884 22936 39344 22964
rect 39393 22967 39451 22973
rect 37884 22924 37890 22936
rect 39393 22933 39405 22967
rect 39439 22964 39451 22967
rect 39942 22964 39948 22976
rect 39439 22936 39948 22964
rect 39439 22933 39451 22936
rect 39393 22927 39451 22933
rect 39942 22924 39948 22936
rect 40000 22924 40006 22976
rect 40037 22967 40095 22973
rect 40037 22933 40049 22967
rect 40083 22964 40095 22967
rect 40126 22964 40132 22976
rect 40083 22936 40132 22964
rect 40083 22933 40095 22936
rect 40037 22927 40095 22933
rect 40126 22924 40132 22936
rect 40184 22924 40190 22976
rect 40494 22924 40500 22976
rect 40552 22924 40558 22976
rect 40862 22924 40868 22976
rect 40920 22964 40926 22976
rect 41524 22964 41552 22995
rect 42702 22992 42708 23044
rect 42760 22992 42766 23044
rect 43257 23035 43315 23041
rect 43257 23001 43269 23035
rect 43303 23032 43315 23035
rect 43530 23032 43536 23044
rect 43303 23004 43536 23032
rect 43303 23001 43315 23004
rect 43257 22995 43315 23001
rect 43530 22992 43536 23004
rect 43588 22992 43594 23044
rect 44726 22992 44732 23044
rect 44784 23032 44790 23044
rect 45370 23032 45376 23044
rect 44784 23004 45376 23032
rect 44784 22992 44790 23004
rect 45370 22992 45376 23004
rect 45428 22992 45434 23044
rect 46014 22992 46020 23044
rect 46072 22992 46078 23044
rect 46201 23035 46259 23041
rect 46201 23001 46213 23035
rect 46247 23032 46259 23035
rect 47302 23032 47308 23044
rect 46247 23004 47308 23032
rect 46247 23001 46259 23004
rect 46201 22995 46259 23001
rect 47302 22992 47308 23004
rect 47360 22992 47366 23044
rect 47780 23032 47808 23063
rect 48590 23032 48596 23044
rect 47780 23004 48596 23032
rect 48590 22992 48596 23004
rect 48648 22992 48654 23044
rect 43714 22964 43720 22976
rect 40920 22936 43720 22964
rect 40920 22924 40926 22936
rect 43714 22924 43720 22936
rect 43772 22924 43778 22976
rect 46934 22924 46940 22976
rect 46992 22964 46998 22976
rect 47581 22967 47639 22973
rect 47581 22964 47593 22967
rect 46992 22936 47593 22964
rect 46992 22924 46998 22936
rect 47581 22933 47593 22936
rect 47627 22933 47639 22967
rect 47581 22927 47639 22933
rect 47670 22924 47676 22976
rect 47728 22964 47734 22976
rect 47946 22964 47952 22976
rect 47728 22936 47952 22964
rect 47728 22924 47734 22936
rect 47946 22924 47952 22936
rect 48004 22924 48010 22976
rect 49326 22924 49332 22976
rect 49384 22964 49390 22976
rect 49421 22967 49479 22973
rect 49421 22964 49433 22967
rect 49384 22936 49433 22964
rect 49384 22924 49390 22936
rect 49421 22933 49433 22936
rect 49467 22933 49479 22967
rect 49421 22927 49479 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 3418 22760 3424 22772
rect 1636 22732 3424 22760
rect 1636 22720 1642 22732
rect 3418 22720 3424 22732
rect 3476 22720 3482 22772
rect 18601 22763 18659 22769
rect 3896 22732 14044 22760
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3896 22624 3924 22732
rect 4798 22652 4804 22704
rect 4856 22652 4862 22704
rect 7098 22652 7104 22704
rect 7156 22652 7162 22704
rect 9950 22652 9956 22704
rect 10008 22652 10014 22704
rect 12802 22652 12808 22704
rect 12860 22652 12866 22704
rect 14016 22692 14044 22732
rect 18601 22729 18613 22763
rect 18647 22760 18659 22763
rect 18690 22760 18696 22772
rect 18647 22732 18696 22760
rect 18647 22729 18659 22732
rect 18601 22723 18659 22729
rect 18690 22720 18696 22732
rect 18748 22720 18754 22772
rect 19153 22763 19211 22769
rect 19153 22729 19165 22763
rect 19199 22760 19211 22763
rect 19334 22760 19340 22772
rect 19199 22732 19340 22760
rect 19199 22729 19211 22732
rect 19153 22723 19211 22729
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 21174 22720 21180 22772
rect 21232 22720 21238 22772
rect 22186 22720 22192 22772
rect 22244 22760 22250 22772
rect 25038 22760 25044 22772
rect 22244 22732 25044 22760
rect 22244 22720 22250 22732
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 26234 22720 26240 22772
rect 26292 22760 26298 22772
rect 26292 22732 26556 22760
rect 26292 22720 26298 22732
rect 15010 22692 15016 22704
rect 14016 22664 15016 22692
rect 15010 22652 15016 22664
rect 15068 22652 15074 22704
rect 15102 22652 15108 22704
rect 15160 22652 15166 22704
rect 17586 22652 17592 22704
rect 17644 22652 17650 22704
rect 3007 22596 3924 22624
rect 3973 22627 4031 22633
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 3973 22593 3985 22627
rect 4019 22593 4031 22627
rect 3973 22587 4031 22593
rect 2501 22559 2559 22565
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 3988 22556 4016 22587
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 7190 22624 7196 22636
rect 6687 22596 7196 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 7466 22584 7472 22636
rect 7524 22584 7530 22636
rect 11146 22584 11152 22636
rect 11204 22584 11210 22636
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22624 11943 22627
rect 13630 22624 13636 22636
rect 11931 22596 13636 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 7282 22556 7288 22568
rect 2547 22528 2774 22556
rect 3988 22528 7288 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 2746 22500 2774 22528
rect 7282 22516 7288 22528
rect 7340 22516 7346 22568
rect 7374 22516 7380 22568
rect 7432 22556 7438 22568
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7432 22528 7941 22556
rect 7432 22516 7438 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 7929 22519 7987 22525
rect 9309 22559 9367 22565
rect 9309 22525 9321 22559
rect 9355 22556 9367 22559
rect 11900 22556 11928 22587
rect 13630 22584 13636 22596
rect 13688 22584 13694 22636
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22624 14059 22627
rect 14642 22624 14648 22636
rect 14047 22596 14648 22624
rect 14047 22593 14059 22596
rect 14001 22587 14059 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16574 22624 16580 22636
rect 16347 22596 16580 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 16850 22584 16856 22636
rect 16908 22584 16914 22636
rect 19352 22624 19380 22720
rect 21082 22692 21088 22704
rect 20930 22664 21088 22692
rect 21082 22652 21088 22664
rect 21140 22652 21146 22704
rect 24026 22652 24032 22704
rect 24084 22692 24090 22704
rect 24121 22695 24179 22701
rect 24121 22692 24133 22695
rect 24084 22664 24133 22692
rect 24084 22652 24090 22664
rect 24121 22661 24133 22664
rect 24167 22692 24179 22695
rect 24578 22692 24584 22704
rect 24167 22664 24584 22692
rect 24167 22661 24179 22664
rect 24121 22655 24179 22661
rect 24578 22652 24584 22664
rect 24636 22652 24642 22704
rect 25774 22652 25780 22704
rect 25832 22652 25838 22704
rect 26326 22652 26332 22704
rect 26384 22652 26390 22704
rect 26528 22692 26556 22732
rect 26602 22720 26608 22772
rect 26660 22760 26666 22772
rect 26660 22732 29776 22760
rect 26660 22720 26666 22732
rect 27798 22692 27804 22704
rect 26528 22664 27804 22692
rect 27798 22652 27804 22664
rect 27856 22652 27862 22704
rect 29270 22692 29276 22704
rect 29118 22664 29276 22692
rect 29270 22652 29276 22664
rect 29328 22692 29334 22704
rect 29454 22692 29460 22704
rect 29328 22664 29460 22692
rect 29328 22652 29334 22664
rect 29454 22652 29460 22664
rect 29512 22652 29518 22704
rect 29748 22692 29776 22732
rect 30466 22720 30472 22772
rect 30524 22760 30530 22772
rect 32309 22763 32367 22769
rect 32309 22760 32321 22763
rect 30524 22732 32321 22760
rect 30524 22720 30530 22732
rect 32309 22729 32321 22732
rect 32355 22729 32367 22763
rect 32309 22723 32367 22729
rect 32677 22763 32735 22769
rect 32677 22729 32689 22763
rect 32723 22760 32735 22763
rect 35250 22760 35256 22772
rect 32723 22732 35256 22760
rect 32723 22729 32735 22732
rect 32677 22723 32735 22729
rect 35250 22720 35256 22732
rect 35308 22720 35314 22772
rect 35434 22720 35440 22772
rect 35492 22720 35498 22772
rect 35526 22720 35532 22772
rect 35584 22760 35590 22772
rect 36081 22763 36139 22769
rect 36081 22760 36093 22763
rect 35584 22732 36093 22760
rect 35584 22720 35590 22732
rect 36081 22729 36093 22732
rect 36127 22729 36139 22763
rect 36081 22723 36139 22729
rect 36354 22720 36360 22772
rect 36412 22760 36418 22772
rect 37274 22760 37280 22772
rect 36412 22732 37280 22760
rect 36412 22720 36418 22732
rect 37274 22720 37280 22732
rect 37332 22720 37338 22772
rect 37458 22720 37464 22772
rect 37516 22720 37522 22772
rect 38286 22720 38292 22772
rect 38344 22760 38350 22772
rect 38838 22760 38844 22772
rect 38344 22732 38844 22760
rect 38344 22720 38350 22732
rect 38838 22720 38844 22732
rect 38896 22720 38902 22772
rect 39482 22720 39488 22772
rect 39540 22720 39546 22772
rect 39758 22720 39764 22772
rect 39816 22720 39822 22772
rect 46201 22763 46259 22769
rect 46201 22760 46213 22763
rect 40604 22732 46213 22760
rect 31386 22692 31392 22704
rect 29748 22664 31392 22692
rect 19429 22627 19487 22633
rect 19429 22624 19441 22627
rect 19352 22596 19441 22624
rect 19429 22593 19441 22596
rect 19475 22593 19487 22627
rect 21100 22624 21128 22652
rect 21634 22624 21640 22636
rect 21100 22596 21640 22624
rect 19429 22587 19487 22593
rect 21634 22584 21640 22596
rect 21692 22584 21698 22636
rect 22002 22584 22008 22636
rect 22060 22584 22066 22636
rect 23566 22624 23572 22636
rect 23414 22596 23572 22624
rect 23566 22584 23572 22596
rect 23624 22624 23630 22636
rect 24394 22624 24400 22636
rect 23624 22596 24400 22624
rect 23624 22584 23630 22596
rect 24394 22584 24400 22596
rect 24452 22624 24458 22636
rect 24452 22596 25360 22624
rect 24452 22584 24458 22596
rect 9355 22528 11928 22556
rect 9355 22525 9367 22528
rect 9309 22519 9367 22525
rect 15470 22516 15476 22568
rect 15528 22556 15534 22568
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 15528 22528 17141 22556
rect 15528 22516 15534 22528
rect 17129 22525 17141 22528
rect 17175 22525 17187 22559
rect 17129 22519 17187 22525
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 18874 22556 18880 22568
rect 17552 22528 18880 22556
rect 17552 22516 17558 22528
rect 18874 22516 18880 22528
rect 18932 22516 18938 22568
rect 19058 22516 19064 22568
rect 19116 22556 19122 22568
rect 19242 22556 19248 22568
rect 19116 22528 19248 22556
rect 19116 22516 19122 22528
rect 19242 22516 19248 22528
rect 19300 22516 19306 22568
rect 19702 22516 19708 22568
rect 19760 22516 19766 22568
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 21928 22528 22293 22556
rect 2746 22460 2780 22500
rect 2774 22448 2780 22460
rect 2832 22448 2838 22500
rect 4157 22491 4215 22497
rect 4157 22457 4169 22491
rect 4203 22488 4215 22491
rect 6362 22488 6368 22500
rect 4203 22460 6368 22488
rect 4203 22457 4215 22460
rect 4157 22451 4215 22457
rect 6362 22448 6368 22460
rect 6420 22448 6426 22500
rect 6825 22491 6883 22497
rect 6825 22457 6837 22491
rect 6871 22488 6883 22491
rect 9122 22488 9128 22500
rect 6871 22460 9128 22488
rect 6871 22457 6883 22460
rect 6825 22451 6883 22457
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 11238 22448 11244 22500
rect 11296 22488 11302 22500
rect 11701 22491 11759 22497
rect 11701 22488 11713 22491
rect 11296 22460 11713 22488
rect 11296 22448 11302 22460
rect 11701 22457 11713 22460
rect 11747 22457 11759 22491
rect 11974 22488 11980 22500
rect 11701 22451 11759 22457
rect 11808 22460 11980 22488
rect 2958 22380 2964 22432
rect 3016 22420 3022 22432
rect 5994 22420 6000 22432
rect 3016 22392 6000 22420
rect 3016 22380 3022 22392
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 9493 22423 9551 22429
rect 9493 22389 9505 22423
rect 9539 22420 9551 22423
rect 11808 22420 11836 22460
rect 11974 22448 11980 22460
rect 12032 22488 12038 22500
rect 12032 22460 16988 22488
rect 12032 22448 12038 22460
rect 9539 22392 11836 22420
rect 9539 22389 9551 22392
rect 9493 22383 9551 22389
rect 12342 22380 12348 22432
rect 12400 22380 12406 22432
rect 14090 22380 14096 22432
rect 14148 22420 14154 22432
rect 14369 22423 14427 22429
rect 14369 22420 14381 22423
rect 14148 22392 14381 22420
rect 14148 22380 14154 22392
rect 14369 22389 14381 22392
rect 14415 22389 14427 22423
rect 14369 22383 14427 22389
rect 14550 22380 14556 22432
rect 14608 22380 14614 22432
rect 16960 22420 16988 22460
rect 20806 22448 20812 22500
rect 20864 22488 20870 22500
rect 21928 22488 21956 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 25332 22556 25360 22596
rect 26602 22584 26608 22636
rect 26660 22584 26666 22636
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22624 27215 22627
rect 27706 22624 27712 22636
rect 27203 22596 27712 22624
rect 27203 22593 27215 22596
rect 27157 22587 27215 22593
rect 27706 22584 27712 22596
rect 27764 22584 27770 22636
rect 29840 22633 29868 22664
rect 31386 22652 31392 22664
rect 31444 22652 31450 22704
rect 33594 22692 33600 22704
rect 31496 22664 33600 22692
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 30650 22584 30656 22636
rect 30708 22584 30714 22636
rect 30745 22627 30803 22633
rect 30745 22593 30757 22627
rect 30791 22624 30803 22627
rect 31496 22624 31524 22664
rect 33594 22652 33600 22664
rect 33652 22652 33658 22704
rect 34238 22692 34244 22704
rect 33704 22664 34244 22692
rect 30791 22596 31524 22624
rect 30791 22593 30803 22596
rect 30745 22587 30803 22593
rect 31662 22584 31668 22636
rect 31720 22584 31726 22636
rect 32769 22627 32827 22633
rect 32769 22593 32781 22627
rect 32815 22624 32827 22627
rect 33410 22624 33416 22636
rect 32815 22596 33416 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 33410 22584 33416 22596
rect 33468 22584 33474 22636
rect 33704 22633 33732 22664
rect 34238 22652 34244 22664
rect 34296 22652 34302 22704
rect 34514 22652 34520 22704
rect 34572 22652 34578 22704
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 36354 22584 36360 22636
rect 36412 22624 36418 22636
rect 36449 22627 36507 22633
rect 36449 22624 36461 22627
rect 36412 22596 36461 22624
rect 36412 22584 36418 22596
rect 36449 22593 36461 22596
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 25774 22556 25780 22568
rect 25332 22528 25780 22556
rect 22281 22519 22339 22525
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 27614 22516 27620 22568
rect 27672 22556 27678 22568
rect 28074 22556 28080 22568
rect 27672 22528 28080 22556
rect 27672 22516 27678 22528
rect 28074 22516 28080 22528
rect 28132 22516 28138 22568
rect 29178 22516 29184 22568
rect 29236 22556 29242 22568
rect 29549 22559 29607 22565
rect 29549 22556 29561 22559
rect 29236 22528 29561 22556
rect 29236 22516 29242 22528
rect 29549 22525 29561 22528
rect 29595 22556 29607 22559
rect 29595 22528 29868 22556
rect 29595 22525 29607 22528
rect 29549 22519 29607 22525
rect 20864 22460 21956 22488
rect 20864 22448 20870 22460
rect 24210 22448 24216 22500
rect 24268 22488 24274 22500
rect 24489 22491 24547 22497
rect 24489 22488 24501 22491
rect 24268 22460 24501 22488
rect 24268 22448 24274 22460
rect 24489 22457 24501 22460
rect 24535 22457 24547 22491
rect 24489 22451 24547 22457
rect 27338 22448 27344 22500
rect 27396 22448 27402 22500
rect 27430 22448 27436 22500
rect 27488 22488 27494 22500
rect 29840 22488 29868 22528
rect 29914 22516 29920 22568
rect 29972 22556 29978 22568
rect 30837 22559 30895 22565
rect 30837 22556 30849 22559
rect 29972 22528 30849 22556
rect 29972 22516 29978 22528
rect 30837 22525 30849 22528
rect 30883 22525 30895 22559
rect 32861 22559 32919 22565
rect 30837 22519 30895 22525
rect 30944 22528 31754 22556
rect 27488 22460 28212 22488
rect 29840 22460 30420 22488
rect 27488 22448 27494 22460
rect 20990 22420 20996 22432
rect 16960 22392 20996 22420
rect 20990 22380 20996 22392
rect 21048 22380 21054 22432
rect 23753 22423 23811 22429
rect 23753 22389 23765 22423
rect 23799 22420 23811 22423
rect 24026 22420 24032 22432
rect 23799 22392 24032 22420
rect 23799 22389 23811 22392
rect 23753 22383 23811 22389
rect 24026 22380 24032 22392
rect 24084 22380 24090 22432
rect 24578 22380 24584 22432
rect 24636 22420 24642 22432
rect 24762 22420 24768 22432
rect 24636 22392 24768 22420
rect 24636 22380 24642 22392
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 24854 22380 24860 22432
rect 24912 22380 24918 22432
rect 25774 22380 25780 22432
rect 25832 22420 25838 22432
rect 27246 22420 27252 22432
rect 25832 22392 27252 22420
rect 25832 22380 25838 22392
rect 27246 22380 27252 22392
rect 27304 22420 27310 22432
rect 27709 22423 27767 22429
rect 27709 22420 27721 22423
rect 27304 22392 27721 22420
rect 27304 22380 27310 22392
rect 27709 22389 27721 22392
rect 27755 22420 27767 22423
rect 27890 22420 27896 22432
rect 27755 22392 27896 22420
rect 27755 22389 27767 22392
rect 27709 22383 27767 22389
rect 27890 22380 27896 22392
rect 27948 22380 27954 22432
rect 28184 22420 28212 22460
rect 30285 22423 30343 22429
rect 30285 22420 30297 22423
rect 28184 22392 30297 22420
rect 30285 22389 30297 22392
rect 30331 22389 30343 22423
rect 30392 22420 30420 22460
rect 30944 22420 30972 22528
rect 31018 22448 31024 22500
rect 31076 22488 31082 22500
rect 31726 22488 31754 22528
rect 32861 22525 32873 22559
rect 32907 22525 32919 22559
rect 33962 22556 33968 22568
rect 32861 22519 32919 22525
rect 33704 22528 33968 22556
rect 32876 22488 32904 22519
rect 33704 22500 33732 22528
rect 33962 22516 33968 22528
rect 34020 22516 34026 22568
rect 36262 22516 36268 22568
rect 36320 22556 36326 22568
rect 36541 22559 36599 22565
rect 36541 22556 36553 22559
rect 36320 22528 36553 22556
rect 36320 22516 36326 22528
rect 36541 22525 36553 22528
rect 36587 22525 36599 22559
rect 36541 22519 36599 22525
rect 36725 22559 36783 22565
rect 36725 22525 36737 22559
rect 36771 22556 36783 22559
rect 37476 22556 37504 22720
rect 37642 22652 37648 22704
rect 37700 22692 37706 22704
rect 37700 22664 37766 22692
rect 37700 22652 37706 22664
rect 38654 22652 38660 22704
rect 38712 22692 38718 22704
rect 38933 22695 38991 22701
rect 38933 22692 38945 22695
rect 38712 22664 38945 22692
rect 38712 22652 38718 22664
rect 38933 22661 38945 22664
rect 38979 22661 38991 22695
rect 38933 22655 38991 22661
rect 39209 22627 39267 22633
rect 39209 22593 39221 22627
rect 39255 22624 39267 22627
rect 39500 22624 39528 22720
rect 40405 22695 40463 22701
rect 40405 22692 40417 22695
rect 40328 22664 40417 22692
rect 39255 22596 39528 22624
rect 39255 22593 39267 22596
rect 39209 22587 39267 22593
rect 40218 22584 40224 22636
rect 40276 22624 40282 22636
rect 40328 22624 40356 22664
rect 40405 22661 40417 22664
rect 40451 22661 40463 22695
rect 40405 22655 40463 22661
rect 40276 22596 40356 22624
rect 40497 22627 40555 22633
rect 40276 22584 40282 22596
rect 40497 22593 40509 22627
rect 40543 22624 40555 22627
rect 40604 22624 40632 22732
rect 46201 22729 46213 22732
rect 46247 22729 46259 22763
rect 46201 22723 46259 22729
rect 47026 22720 47032 22772
rect 47084 22720 47090 22772
rect 47673 22763 47731 22769
rect 47673 22729 47685 22763
rect 47719 22760 47731 22763
rect 47762 22760 47768 22772
rect 47719 22732 47768 22760
rect 47719 22729 47731 22732
rect 47673 22723 47731 22729
rect 40862 22652 40868 22704
rect 40920 22692 40926 22704
rect 40920 22664 43576 22692
rect 40920 22652 40926 22664
rect 40543 22596 40632 22624
rect 40543 22593 40555 22596
rect 40497 22587 40555 22593
rect 41322 22584 41328 22636
rect 41380 22624 41386 22636
rect 41417 22627 41475 22633
rect 41417 22624 41429 22627
rect 41380 22596 41429 22624
rect 41380 22584 41386 22596
rect 41417 22593 41429 22596
rect 41463 22593 41475 22627
rect 41417 22587 41475 22593
rect 42058 22584 42064 22636
rect 42116 22584 42122 22636
rect 42610 22584 42616 22636
rect 42668 22584 42674 22636
rect 43548 22624 43576 22664
rect 43714 22652 43720 22704
rect 43772 22652 43778 22704
rect 44082 22652 44088 22704
rect 44140 22692 44146 22704
rect 44266 22692 44272 22704
rect 44140 22664 44272 22692
rect 44140 22652 44146 22664
rect 44266 22652 44272 22664
rect 44324 22692 44330 22704
rect 44361 22695 44419 22701
rect 44361 22692 44373 22695
rect 44324 22664 44373 22692
rect 44324 22652 44330 22664
rect 44361 22661 44373 22664
rect 44407 22661 44419 22695
rect 47688 22692 47716 22723
rect 47762 22720 47768 22732
rect 47820 22720 47826 22772
rect 48041 22763 48099 22769
rect 48041 22729 48053 22763
rect 48087 22760 48099 22763
rect 48590 22760 48596 22772
rect 48087 22732 48596 22760
rect 48087 22729 48099 22732
rect 48041 22723 48099 22729
rect 48590 22720 48596 22732
rect 48648 22720 48654 22772
rect 44361 22655 44419 22661
rect 46400 22664 47716 22692
rect 45097 22627 45155 22633
rect 45097 22624 45109 22627
rect 43548 22596 45109 22624
rect 45097 22593 45109 22596
rect 45143 22624 45155 22627
rect 45186 22624 45192 22636
rect 45143 22596 45192 22624
rect 45143 22593 45155 22596
rect 45097 22587 45155 22593
rect 45186 22584 45192 22596
rect 45244 22584 45250 22636
rect 45738 22584 45744 22636
rect 45796 22584 45802 22636
rect 46400 22633 46428 22664
rect 46385 22627 46443 22633
rect 46385 22593 46397 22627
rect 46431 22593 46443 22627
rect 46385 22587 46443 22593
rect 47210 22584 47216 22636
rect 47268 22624 47274 22636
rect 47765 22627 47823 22633
rect 47765 22624 47777 22627
rect 47268 22596 47777 22624
rect 47268 22584 47274 22596
rect 47765 22593 47777 22596
rect 47811 22593 47823 22627
rect 47765 22587 47823 22593
rect 48593 22627 48651 22633
rect 48593 22593 48605 22627
rect 48639 22624 48651 22627
rect 49234 22624 49240 22636
rect 48639 22596 49240 22624
rect 48639 22593 48651 22596
rect 48593 22587 48651 22593
rect 49234 22584 49240 22596
rect 49292 22584 49298 22636
rect 49329 22627 49387 22633
rect 49329 22593 49341 22627
rect 49375 22593 49387 22627
rect 49329 22587 49387 22593
rect 40589 22559 40647 22565
rect 40589 22556 40601 22559
rect 36771 22528 37504 22556
rect 37844 22528 40601 22556
rect 36771 22525 36783 22528
rect 36725 22519 36783 22525
rect 31076 22460 31616 22488
rect 31726 22460 32904 22488
rect 31076 22448 31082 22460
rect 30392 22392 30972 22420
rect 30285 22383 30343 22389
rect 31478 22380 31484 22432
rect 31536 22380 31542 22432
rect 31588 22420 31616 22460
rect 33686 22448 33692 22500
rect 33744 22448 33750 22500
rect 36630 22448 36636 22500
rect 36688 22488 36694 22500
rect 36906 22488 36912 22500
rect 36688 22460 36912 22488
rect 36688 22448 36694 22460
rect 36906 22448 36912 22460
rect 36964 22488 36970 22500
rect 37844 22488 37872 22528
rect 40589 22525 40601 22528
rect 40635 22525 40647 22559
rect 40589 22519 40647 22525
rect 42076 22488 42104 22584
rect 42889 22559 42947 22565
rect 42889 22525 42901 22559
rect 42935 22556 42947 22559
rect 43714 22556 43720 22568
rect 42935 22528 43720 22556
rect 42935 22525 42947 22528
rect 42889 22519 42947 22525
rect 43714 22516 43720 22528
rect 43772 22516 43778 22568
rect 47670 22516 47676 22568
rect 47728 22556 47734 22568
rect 49344 22556 49372 22587
rect 49418 22556 49424 22568
rect 47728 22528 49424 22556
rect 47728 22516 47734 22528
rect 49418 22516 49424 22528
rect 49476 22516 49482 22568
rect 36964 22460 37872 22488
rect 39592 22460 42104 22488
rect 36964 22448 36970 22460
rect 33413 22423 33471 22429
rect 33413 22420 33425 22423
rect 31588 22392 33425 22420
rect 33413 22389 33425 22392
rect 33459 22420 33471 22423
rect 35066 22420 35072 22432
rect 33459 22392 35072 22420
rect 33459 22389 33471 22392
rect 33413 22383 33471 22389
rect 35066 22380 35072 22392
rect 35124 22420 35130 22432
rect 35805 22423 35863 22429
rect 35805 22420 35817 22423
rect 35124 22392 35817 22420
rect 35124 22380 35130 22392
rect 35805 22389 35817 22392
rect 35851 22420 35863 22423
rect 38562 22420 38568 22432
rect 35851 22392 38568 22420
rect 35851 22389 35863 22392
rect 35805 22383 35863 22389
rect 38562 22380 38568 22392
rect 38620 22380 38626 22432
rect 38930 22380 38936 22432
rect 38988 22420 38994 22432
rect 39592 22420 39620 22460
rect 43438 22448 43444 22500
rect 43496 22488 43502 22500
rect 44913 22491 44971 22497
rect 44913 22488 44925 22491
rect 43496 22460 44925 22488
rect 43496 22448 43502 22460
rect 44913 22457 44925 22460
rect 44959 22457 44971 22491
rect 44913 22451 44971 22457
rect 45554 22448 45560 22500
rect 45612 22448 45618 22500
rect 38988 22392 39620 22420
rect 38988 22380 38994 22392
rect 40034 22380 40040 22432
rect 40092 22380 40098 22432
rect 40126 22380 40132 22432
rect 40184 22420 40190 22432
rect 40862 22420 40868 22432
rect 40184 22392 40868 22420
rect 40184 22380 40190 22392
rect 40862 22380 40868 22392
rect 40920 22380 40926 22432
rect 41230 22380 41236 22432
rect 41288 22380 41294 22432
rect 41874 22380 41880 22432
rect 41932 22380 41938 22432
rect 43530 22380 43536 22432
rect 43588 22420 43594 22432
rect 44269 22423 44327 22429
rect 44269 22420 44281 22423
rect 43588 22392 44281 22420
rect 43588 22380 43594 22392
rect 44269 22389 44281 22392
rect 44315 22389 44327 22423
rect 44269 22383 44327 22389
rect 48406 22380 48412 22432
rect 48464 22380 48470 22432
rect 48498 22380 48504 22432
rect 48556 22420 48562 22432
rect 49145 22423 49203 22429
rect 49145 22420 49157 22423
rect 48556 22392 49157 22420
rect 48556 22380 48562 22392
rect 49145 22389 49157 22392
rect 49191 22389 49203 22423
rect 49145 22383 49203 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 4246 22216 4252 22228
rect 2280 22188 4252 22216
rect 2280 22176 2286 22188
rect 4246 22176 4252 22188
rect 4304 22176 4310 22228
rect 11882 22176 11888 22228
rect 11940 22216 11946 22228
rect 12345 22219 12403 22225
rect 12345 22216 12357 22219
rect 11940 22188 12357 22216
rect 11940 22176 11946 22188
rect 12345 22185 12357 22188
rect 12391 22185 12403 22219
rect 15197 22219 15255 22225
rect 15197 22216 15209 22219
rect 12345 22179 12403 22185
rect 13648 22188 15209 22216
rect 3970 22108 3976 22160
rect 4028 22148 4034 22160
rect 4028 22120 6040 22148
rect 4028 22108 4034 22120
rect 6012 22089 6040 22120
rect 5997 22083 6055 22089
rect 5997 22049 6009 22083
rect 6043 22049 6055 22083
rect 9674 22080 9680 22092
rect 5997 22043 6055 22049
rect 7852 22052 9680 22080
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 21981 3019 22015
rect 2961 21975 3019 21981
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 22012 5411 22015
rect 6822 22012 6828 22024
rect 5399 21984 6828 22012
rect 5399 21981 5411 21984
rect 5353 21975 5411 21981
rect 1026 21904 1032 21956
rect 1084 21944 1090 21956
rect 1765 21947 1823 21953
rect 1765 21944 1777 21947
rect 1084 21916 1777 21944
rect 1084 21904 1090 21916
rect 1765 21913 1777 21916
rect 1811 21913 1823 21947
rect 1765 21907 1823 21913
rect 2976 21876 3004 21975
rect 6822 21972 6828 21984
rect 6880 21972 6886 22024
rect 7852 22021 7880 22052
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 11885 22083 11943 22089
rect 11885 22049 11897 22083
rect 11931 22080 11943 22083
rect 11974 22080 11980 22092
rect 11931 22052 11980 22080
rect 11931 22049 11943 22052
rect 11885 22043 11943 22049
rect 11974 22040 11980 22052
rect 12032 22040 12038 22092
rect 13262 22080 13268 22092
rect 12452 22052 13268 22080
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22012 7251 22015
rect 7837 22015 7895 22021
rect 7239 21984 7788 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 3234 21904 3240 21956
rect 3292 21944 3298 21956
rect 4157 21947 4215 21953
rect 4157 21944 4169 21947
rect 3292 21916 4169 21944
rect 3292 21904 3298 21916
rect 4157 21913 4169 21916
rect 4203 21913 4215 21947
rect 4157 21907 4215 21913
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 5684 21916 7665 21944
rect 5684 21904 5690 21916
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 7760 21944 7788 21984
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 8478 21944 8484 21956
rect 7760 21916 8484 21944
rect 7653 21907 7711 21913
rect 8478 21904 8484 21916
rect 8536 21904 8542 21956
rect 6730 21876 6736 21888
rect 2976 21848 6736 21876
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 8386 21836 8392 21888
rect 8444 21836 8450 21888
rect 8588 21876 8616 21975
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 12452 22012 12480 22052
rect 13262 22040 13268 22052
rect 13320 22040 13326 22092
rect 13648 22089 13676 22188
rect 15197 22185 15209 22188
rect 15243 22216 15255 22219
rect 15470 22216 15476 22228
rect 15243 22188 15476 22216
rect 15243 22185 15255 22188
rect 15197 22179 15255 22185
rect 15470 22176 15476 22188
rect 15528 22176 15534 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 17218 22216 17224 22228
rect 16632 22188 17224 22216
rect 16632 22176 16638 22188
rect 17218 22176 17224 22188
rect 17276 22176 17282 22228
rect 18782 22176 18788 22228
rect 18840 22216 18846 22228
rect 20806 22216 20812 22228
rect 18840 22188 20812 22216
rect 18840 22176 18846 22188
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 21634 22176 21640 22228
rect 21692 22216 21698 22228
rect 23014 22216 23020 22228
rect 21692 22188 23020 22216
rect 21692 22176 21698 22188
rect 23014 22176 23020 22188
rect 23072 22216 23078 22228
rect 23566 22216 23572 22228
rect 23072 22188 23572 22216
rect 23072 22176 23078 22188
rect 23566 22176 23572 22188
rect 23624 22176 23630 22228
rect 24581 22219 24639 22225
rect 24581 22185 24593 22219
rect 24627 22185 24639 22219
rect 24581 22179 24639 22185
rect 17034 22108 17040 22160
rect 17092 22148 17098 22160
rect 17092 22120 17632 22148
rect 17092 22108 17098 22120
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22049 13691 22083
rect 13633 22043 13691 22049
rect 14274 22040 14280 22092
rect 14332 22080 14338 22092
rect 17604 22089 17632 22120
rect 19886 22108 19892 22160
rect 19944 22148 19950 22160
rect 19944 22120 22048 22148
rect 19944 22108 19950 22120
rect 14461 22083 14519 22089
rect 14461 22080 14473 22083
rect 14332 22052 14473 22080
rect 14332 22040 14338 22052
rect 14461 22049 14473 22052
rect 14507 22049 14519 22083
rect 14461 22043 14519 22049
rect 17589 22083 17647 22089
rect 17589 22049 17601 22083
rect 17635 22049 17647 22083
rect 21910 22080 21916 22092
rect 17589 22043 17647 22049
rect 19306 22052 21916 22080
rect 11655 21984 12480 22012
rect 12529 22015 12587 22021
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 12529 21981 12541 22015
rect 12575 22008 12587 22015
rect 13538 22012 13544 22024
rect 12636 22008 13544 22012
rect 12575 21984 13544 22008
rect 12575 21981 12664 21984
rect 12529 21980 12664 21981
rect 12529 21975 12587 21980
rect 13538 21972 13544 21984
rect 13596 21972 13602 22024
rect 16942 21972 16948 22024
rect 17000 21972 17006 22024
rect 18785 22015 18843 22021
rect 18785 21981 18797 22015
rect 18831 22012 18843 22015
rect 19306 22012 19334 22052
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 22020 22089 22048 22120
rect 24302 22108 24308 22160
rect 24360 22148 24366 22160
rect 24596 22148 24624 22179
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 26694 22216 26700 22228
rect 25188 22188 26700 22216
rect 25188 22176 25194 22188
rect 26694 22176 26700 22188
rect 26752 22176 26758 22228
rect 27154 22176 27160 22228
rect 27212 22176 27218 22228
rect 27890 22176 27896 22228
rect 27948 22216 27954 22228
rect 28994 22216 29000 22228
rect 27948 22188 29000 22216
rect 27948 22176 27954 22188
rect 28994 22176 29000 22188
rect 29052 22216 29058 22228
rect 29454 22216 29460 22228
rect 29052 22188 29460 22216
rect 29052 22176 29058 22188
rect 29454 22176 29460 22188
rect 29512 22216 29518 22228
rect 30006 22216 30012 22228
rect 29512 22188 30012 22216
rect 29512 22176 29518 22188
rect 30006 22176 30012 22188
rect 30064 22176 30070 22228
rect 30190 22176 30196 22228
rect 30248 22216 30254 22228
rect 30285 22219 30343 22225
rect 30285 22216 30297 22219
rect 30248 22188 30297 22216
rect 30248 22176 30254 22188
rect 30285 22185 30297 22188
rect 30331 22216 30343 22219
rect 32122 22216 32128 22228
rect 30331 22188 32128 22216
rect 30331 22185 30343 22188
rect 30285 22179 30343 22185
rect 32122 22176 32128 22188
rect 32180 22176 32186 22228
rect 33594 22176 33600 22228
rect 33652 22216 33658 22228
rect 34698 22216 34704 22228
rect 33652 22188 34704 22216
rect 33652 22176 33658 22188
rect 34698 22176 34704 22188
rect 34756 22216 34762 22228
rect 37458 22216 37464 22228
rect 34756 22188 37464 22216
rect 34756 22176 34762 22188
rect 37458 22176 37464 22188
rect 37516 22176 37522 22228
rect 38654 22176 38660 22228
rect 38712 22216 38718 22228
rect 40221 22219 40279 22225
rect 38712 22188 40172 22216
rect 38712 22176 38718 22188
rect 24854 22148 24860 22160
rect 24360 22120 24624 22148
rect 24688 22120 24860 22148
rect 24360 22108 24366 22120
rect 22005 22083 22063 22089
rect 22005 22049 22017 22083
rect 22051 22049 22063 22083
rect 22005 22043 22063 22049
rect 22646 22040 22652 22092
rect 22704 22080 22710 22092
rect 23201 22083 23259 22089
rect 23201 22080 23213 22083
rect 22704 22052 23213 22080
rect 22704 22040 22710 22052
rect 23201 22049 23213 22052
rect 23247 22080 23259 22083
rect 24688 22080 24716 22120
rect 24854 22108 24860 22120
rect 24912 22108 24918 22160
rect 25961 22151 26019 22157
rect 25961 22117 25973 22151
rect 26007 22117 26019 22151
rect 25961 22111 26019 22117
rect 23247 22052 24716 22080
rect 23247 22049 23259 22052
rect 23201 22043 23259 22049
rect 24762 22040 24768 22092
rect 24820 22080 24826 22092
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 24820 22052 25053 22080
rect 24820 22040 24826 22052
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25041 22043 25099 22049
rect 18831 21984 19334 22012
rect 18831 21981 18843 21984
rect 18785 21975 18843 21981
rect 19426 21972 19432 22024
rect 19484 21972 19490 22024
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 22012 21235 22015
rect 22370 22012 22376 22024
rect 21223 21984 22376 22012
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 22370 21972 22376 21984
rect 22428 22012 22434 22024
rect 22830 22012 22836 22024
rect 22428 21984 22836 22012
rect 22428 21972 22434 21984
rect 22830 21972 22836 21984
rect 22888 21972 22894 22024
rect 23934 22012 23940 22024
rect 22940 21984 23940 22012
rect 13262 21904 13268 21956
rect 13320 21944 13326 21956
rect 13320 21916 14596 21944
rect 13320 21904 13326 21916
rect 12989 21879 13047 21885
rect 12989 21876 13001 21879
rect 8588 21848 13001 21876
rect 12989 21845 13001 21848
rect 13035 21845 13047 21879
rect 12989 21839 13047 21845
rect 13354 21836 13360 21888
rect 13412 21836 13418 21888
rect 13449 21879 13507 21885
rect 13449 21845 13461 21879
rect 13495 21876 13507 21879
rect 13906 21876 13912 21888
rect 13495 21848 13912 21876
rect 13495 21845 13507 21848
rect 13449 21839 13507 21845
rect 13906 21836 13912 21848
rect 13964 21836 13970 21888
rect 14090 21836 14096 21888
rect 14148 21836 14154 21888
rect 14568 21876 14596 21916
rect 14642 21904 14648 21956
rect 14700 21904 14706 21956
rect 15286 21904 15292 21956
rect 15344 21944 15350 21956
rect 15344 21916 15502 21944
rect 15344 21904 15350 21916
rect 16574 21904 16580 21956
rect 16632 21944 16638 21956
rect 16669 21947 16727 21953
rect 16669 21944 16681 21947
rect 16632 21916 16681 21944
rect 16632 21904 16638 21916
rect 16669 21913 16681 21916
rect 16715 21913 16727 21947
rect 16669 21907 16727 21913
rect 17126 21904 17132 21956
rect 17184 21944 17190 21956
rect 18874 21944 18880 21956
rect 17184 21916 18880 21944
rect 17184 21904 17190 21916
rect 18874 21904 18880 21916
rect 18932 21904 18938 21956
rect 18966 21904 18972 21956
rect 19024 21944 19030 21956
rect 20349 21947 20407 21953
rect 20349 21944 20361 21947
rect 19024 21916 20361 21944
rect 19024 21904 19030 21916
rect 20349 21913 20361 21916
rect 20395 21913 20407 21947
rect 20349 21907 20407 21913
rect 20622 21904 20628 21956
rect 20680 21944 20686 21956
rect 21821 21947 21879 21953
rect 20680 21916 21496 21944
rect 20680 21904 20686 21916
rect 21082 21876 21088 21888
rect 14568 21848 21088 21876
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 21468 21885 21496 21916
rect 21821 21913 21833 21947
rect 21867 21913 21879 21947
rect 21821 21907 21879 21913
rect 21913 21947 21971 21953
rect 21913 21913 21925 21947
rect 21959 21944 21971 21947
rect 22940 21944 22968 21984
rect 23934 21972 23940 21984
rect 23992 21972 23998 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 24946 22012 24952 22024
rect 24075 21984 24952 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25056 22012 25084 22043
rect 25130 22040 25136 22092
rect 25188 22040 25194 22092
rect 25222 22040 25228 22092
rect 25280 22080 25286 22092
rect 25976 22080 26004 22111
rect 28258 22108 28264 22160
rect 28316 22148 28322 22160
rect 28353 22151 28411 22157
rect 28353 22148 28365 22151
rect 28316 22120 28365 22148
rect 28316 22108 28322 22120
rect 28353 22117 28365 22120
rect 28399 22117 28411 22151
rect 35434 22148 35440 22160
rect 28353 22111 28411 22117
rect 33704 22120 35440 22148
rect 25280 22052 26004 22080
rect 25280 22040 25286 22052
rect 26602 22040 26608 22092
rect 26660 22040 26666 22092
rect 27522 22040 27528 22092
rect 27580 22080 27586 22092
rect 27709 22083 27767 22089
rect 27709 22080 27721 22083
rect 27580 22052 27721 22080
rect 27580 22040 27586 22052
rect 27709 22049 27721 22052
rect 27755 22049 27767 22083
rect 27709 22043 27767 22049
rect 28074 22040 28080 22092
rect 28132 22080 28138 22092
rect 28902 22080 28908 22092
rect 28132 22052 28908 22080
rect 28132 22040 28138 22052
rect 28902 22040 28908 22052
rect 28960 22040 28966 22092
rect 29178 22040 29184 22092
rect 29236 22080 29242 22092
rect 29454 22080 29460 22092
rect 29236 22052 29460 22080
rect 29236 22040 29242 22052
rect 29454 22040 29460 22052
rect 29512 22040 29518 22092
rect 30558 22080 30564 22092
rect 29840 22052 30564 22080
rect 25866 22012 25872 22024
rect 25056 21984 25872 22012
rect 25866 21972 25872 21984
rect 25924 21972 25930 22024
rect 26421 22015 26479 22021
rect 26421 21981 26433 22015
rect 26467 22012 26479 22015
rect 27430 22012 27436 22024
rect 26467 21984 27436 22012
rect 26467 21981 26479 21984
rect 26421 21975 26479 21981
rect 27430 21972 27436 21984
rect 27488 21972 27494 22024
rect 27614 21972 27620 22024
rect 27672 21972 27678 22024
rect 28721 22015 28779 22021
rect 28721 21981 28733 22015
rect 28767 22012 28779 22015
rect 29840 22012 29868 22052
rect 30558 22040 30564 22052
rect 30616 22040 30622 22092
rect 31478 22080 31484 22092
rect 30852 22052 31484 22080
rect 30852 22024 30880 22052
rect 31478 22040 31484 22052
rect 31536 22040 31542 22092
rect 33704 22089 33732 22120
rect 35434 22108 35440 22120
rect 35492 22108 35498 22160
rect 37826 22148 37832 22160
rect 36280 22120 37832 22148
rect 33689 22083 33747 22089
rect 33689 22049 33701 22083
rect 33735 22080 33747 22083
rect 34425 22083 34483 22089
rect 34425 22080 34437 22083
rect 33735 22052 33769 22080
rect 34072 22052 34437 22080
rect 33735 22049 33747 22052
rect 33689 22043 33747 22049
rect 28767 21984 29868 22012
rect 28767 21981 28779 21984
rect 28721 21975 28779 21981
rect 29914 21972 29920 22024
rect 29972 21972 29978 22024
rect 30834 21972 30840 22024
rect 30892 21972 30898 22024
rect 32398 21972 32404 22024
rect 32456 22012 32462 22024
rect 34072 22021 34100 22052
rect 34425 22049 34437 22052
rect 34471 22080 34483 22083
rect 34514 22080 34520 22092
rect 34471 22052 34520 22080
rect 34471 22049 34483 22052
rect 34425 22043 34483 22049
rect 34514 22040 34520 22052
rect 34572 22040 34578 22092
rect 35066 22040 35072 22092
rect 35124 22040 35130 22092
rect 36173 22083 36231 22089
rect 36173 22049 36185 22083
rect 36219 22080 36231 22083
rect 36280 22080 36308 22120
rect 37826 22108 37832 22120
rect 37884 22108 37890 22160
rect 39393 22151 39451 22157
rect 39393 22117 39405 22151
rect 39439 22148 39451 22151
rect 39482 22148 39488 22160
rect 39439 22120 39488 22148
rect 39439 22117 39451 22120
rect 39393 22111 39451 22117
rect 39482 22108 39488 22120
rect 39540 22148 39546 22160
rect 40144 22148 40172 22188
rect 40221 22185 40233 22219
rect 40267 22216 40279 22219
rect 40494 22216 40500 22228
rect 40267 22188 40500 22216
rect 40267 22185 40279 22188
rect 40221 22179 40279 22185
rect 40494 22176 40500 22188
rect 40552 22176 40558 22228
rect 41414 22176 41420 22228
rect 41472 22176 41478 22228
rect 43165 22219 43223 22225
rect 43165 22185 43177 22219
rect 43211 22216 43223 22219
rect 43530 22216 43536 22228
rect 43211 22188 43536 22216
rect 43211 22185 43223 22188
rect 43165 22179 43223 22185
rect 43530 22176 43536 22188
rect 43588 22176 43594 22228
rect 45186 22176 45192 22228
rect 45244 22176 45250 22228
rect 45370 22176 45376 22228
rect 45428 22176 45434 22228
rect 45649 22219 45707 22225
rect 45649 22185 45661 22219
rect 45695 22216 45707 22219
rect 45738 22216 45744 22228
rect 45695 22188 45744 22216
rect 45695 22185 45707 22188
rect 45649 22179 45707 22185
rect 45738 22176 45744 22188
rect 45796 22176 45802 22228
rect 46842 22176 46848 22228
rect 46900 22216 46906 22228
rect 47029 22219 47087 22225
rect 47029 22216 47041 22219
rect 46900 22188 47041 22216
rect 46900 22176 46906 22188
rect 47029 22185 47041 22188
rect 47075 22185 47087 22219
rect 47029 22179 47087 22185
rect 47578 22176 47584 22228
rect 47636 22176 47642 22228
rect 39540 22120 39565 22148
rect 40144 22120 42012 22148
rect 39540 22108 39546 22120
rect 38470 22080 38476 22092
rect 36219 22052 36308 22080
rect 36372 22052 38476 22080
rect 36219 22049 36231 22052
rect 36173 22043 36231 22049
rect 34057 22015 34115 22021
rect 34057 22012 34069 22015
rect 32456 21984 34069 22012
rect 32456 21972 32462 21984
rect 34057 21981 34069 21984
rect 34103 21981 34115 22015
rect 34057 21975 34115 21981
rect 34238 21972 34244 22024
rect 34296 22012 34302 22024
rect 36372 22012 36400 22052
rect 38470 22040 38476 22052
rect 38528 22040 38534 22092
rect 38838 22040 38844 22092
rect 38896 22040 38902 22092
rect 39117 22083 39175 22089
rect 39117 22049 39129 22083
rect 39163 22080 39175 22083
rect 39500 22080 39528 22108
rect 39163 22052 39528 22080
rect 39163 22049 39175 22052
rect 39117 22043 39175 22049
rect 40494 22040 40500 22092
rect 40552 22080 40558 22092
rect 40681 22083 40739 22089
rect 40681 22080 40693 22083
rect 40552 22052 40693 22080
rect 40552 22040 40558 22052
rect 40681 22049 40693 22052
rect 40727 22049 40739 22083
rect 40788 22080 40816 22120
rect 40865 22083 40923 22089
rect 40865 22080 40877 22083
rect 40788 22052 40877 22080
rect 40681 22043 40739 22049
rect 40865 22049 40877 22052
rect 40911 22049 40923 22083
rect 40865 22043 40923 22049
rect 40954 22040 40960 22092
rect 41012 22080 41018 22092
rect 41138 22080 41144 22092
rect 41012 22052 41144 22080
rect 41012 22040 41018 22052
rect 41138 22040 41144 22052
rect 41196 22040 41202 22092
rect 41874 22080 41880 22092
rect 41386 22052 41880 22080
rect 34296 21984 36400 22012
rect 36449 22015 36507 22021
rect 34296 21972 34302 21984
rect 36449 21981 36461 22015
rect 36495 22012 36507 22015
rect 37458 22012 37464 22024
rect 36495 21984 37464 22012
rect 36495 21981 36507 21984
rect 36449 21975 36507 21981
rect 37458 21972 37464 21984
rect 37516 21972 37522 22024
rect 37734 21972 37740 22024
rect 37792 21972 37798 22024
rect 41386 22012 41414 22052
rect 41874 22040 41880 22052
rect 41932 22040 41938 22092
rect 41984 22089 42012 22120
rect 42058 22108 42064 22160
rect 42116 22148 42122 22160
rect 42702 22148 42708 22160
rect 42116 22120 42708 22148
rect 42116 22108 42122 22120
rect 42702 22108 42708 22120
rect 42760 22148 42766 22160
rect 42760 22120 43944 22148
rect 42760 22108 42766 22120
rect 41969 22083 42027 22089
rect 41969 22049 41981 22083
rect 42015 22080 42027 22083
rect 42015 22052 42049 22080
rect 42015 22049 42027 22052
rect 41969 22043 42027 22049
rect 42150 22040 42156 22092
rect 42208 22080 42214 22092
rect 43254 22080 43260 22092
rect 42208 22052 43260 22080
rect 42208 22040 42214 22052
rect 43254 22040 43260 22052
rect 43312 22040 43318 22092
rect 43916 22080 43944 22120
rect 47136 22120 47440 22148
rect 47136 22094 47164 22120
rect 45005 22083 45063 22089
rect 45005 22080 45017 22083
rect 43916 22052 45017 22080
rect 45005 22049 45017 22052
rect 45051 22049 45063 22083
rect 45005 22043 45063 22049
rect 45094 22040 45100 22092
rect 45152 22080 45158 22092
rect 47044 22080 47164 22094
rect 45152 22066 47164 22080
rect 47412 22080 47440 22120
rect 48041 22083 48099 22089
rect 48041 22080 48053 22083
rect 45152 22052 47072 22066
rect 47412 22052 48053 22080
rect 45152 22040 45158 22052
rect 48041 22049 48053 22052
rect 48087 22049 48099 22083
rect 48041 22043 48099 22049
rect 39132 21984 41414 22012
rect 21959 21916 22968 21944
rect 23017 21947 23075 21953
rect 21959 21913 21971 21916
rect 21913 21907 21971 21913
rect 23017 21913 23029 21947
rect 23063 21944 23075 21947
rect 24578 21944 24584 21956
rect 23063 21916 24584 21944
rect 23063 21913 23075 21916
rect 23017 21907 23075 21913
rect 21453 21879 21511 21885
rect 21453 21845 21465 21879
rect 21499 21845 21511 21879
rect 21836 21876 21864 21907
rect 24578 21904 24584 21916
rect 24636 21904 24642 21956
rect 24762 21904 24768 21956
rect 24820 21944 24826 21956
rect 25685 21947 25743 21953
rect 25685 21944 25697 21947
rect 24820 21916 25697 21944
rect 24820 21904 24826 21916
rect 25685 21913 25697 21916
rect 25731 21944 25743 21947
rect 27525 21947 27583 21953
rect 25731 21916 26372 21944
rect 25731 21913 25743 21916
rect 25685 21907 25743 21913
rect 22462 21876 22468 21888
rect 21836 21848 22468 21876
rect 21453 21839 21511 21845
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 22612 21848 22661 21876
rect 22612 21836 22618 21848
rect 22649 21845 22661 21848
rect 22695 21845 22707 21879
rect 22649 21839 22707 21845
rect 22830 21836 22836 21888
rect 22888 21876 22894 21888
rect 23109 21879 23167 21885
rect 23109 21876 23121 21879
rect 22888 21848 23121 21876
rect 22888 21836 22894 21848
rect 23109 21845 23121 21848
rect 23155 21845 23167 21879
rect 23109 21839 23167 21845
rect 23750 21836 23756 21888
rect 23808 21876 23814 21888
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 23808 21848 23857 21876
rect 23808 21836 23814 21848
rect 23845 21845 23857 21848
rect 23891 21845 23903 21879
rect 23845 21839 23903 21845
rect 24026 21836 24032 21888
rect 24084 21876 24090 21888
rect 24670 21876 24676 21888
rect 24084 21848 24676 21876
rect 24084 21836 24090 21848
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 24854 21836 24860 21888
rect 24912 21876 24918 21888
rect 26344 21885 26372 21916
rect 27525 21913 27537 21947
rect 27571 21944 27583 21947
rect 28350 21944 28356 21956
rect 27571 21916 28356 21944
rect 27571 21913 27583 21916
rect 27525 21907 27583 21913
rect 28350 21904 28356 21916
rect 28408 21944 28414 21956
rect 28813 21947 28871 21953
rect 28408 21916 28580 21944
rect 28408 21904 28414 21916
rect 24949 21879 25007 21885
rect 24949 21876 24961 21879
rect 24912 21848 24961 21876
rect 24912 21836 24918 21848
rect 24949 21845 24961 21848
rect 24995 21845 25007 21879
rect 24949 21839 25007 21845
rect 26329 21879 26387 21885
rect 26329 21845 26341 21879
rect 26375 21876 26387 21879
rect 27614 21876 27620 21888
rect 26375 21848 27620 21876
rect 26375 21845 26387 21848
rect 26329 21839 26387 21845
rect 27614 21836 27620 21848
rect 27672 21836 27678 21888
rect 28552 21876 28580 21916
rect 28813 21913 28825 21947
rect 28859 21944 28871 21947
rect 30466 21944 30472 21956
rect 28859 21916 30472 21944
rect 28859 21913 28871 21916
rect 28813 21907 28871 21913
rect 30466 21904 30472 21916
rect 30524 21904 30530 21956
rect 30742 21904 30748 21956
rect 30800 21944 30806 21956
rect 31113 21947 31171 21953
rect 31113 21944 31125 21947
rect 30800 21916 31125 21944
rect 30800 21904 30806 21916
rect 31113 21913 31125 21916
rect 31159 21913 31171 21947
rect 31113 21907 31171 21913
rect 31386 21904 31392 21956
rect 31444 21944 31450 21956
rect 31444 21916 31602 21944
rect 31444 21904 31450 21916
rect 32766 21904 32772 21956
rect 32824 21944 32830 21956
rect 33505 21947 33563 21953
rect 33505 21944 33517 21947
rect 32824 21916 33517 21944
rect 32824 21904 32830 21916
rect 33505 21913 33517 21916
rect 33551 21913 33563 21947
rect 33505 21907 33563 21913
rect 33870 21904 33876 21956
rect 33928 21944 33934 21956
rect 35161 21947 35219 21953
rect 35161 21944 35173 21947
rect 33928 21916 35173 21944
rect 33928 21904 33934 21916
rect 35161 21913 35173 21916
rect 35207 21944 35219 21947
rect 36998 21944 37004 21956
rect 35207 21916 37004 21944
rect 35207 21913 35219 21916
rect 35161 21907 35219 21913
rect 36998 21904 37004 21916
rect 37056 21904 37062 21956
rect 37274 21904 37280 21956
rect 37332 21944 37338 21956
rect 37332 21916 37504 21944
rect 37332 21904 37338 21916
rect 29178 21876 29184 21888
rect 28552 21848 29184 21876
rect 29178 21836 29184 21848
rect 29236 21836 29242 21888
rect 29730 21836 29736 21888
rect 29788 21836 29794 21888
rect 30374 21836 30380 21888
rect 30432 21836 30438 21888
rect 30558 21836 30564 21888
rect 30616 21876 30622 21888
rect 31938 21876 31944 21888
rect 30616 21848 31944 21876
rect 30616 21836 30622 21848
rect 31938 21836 31944 21848
rect 31996 21836 32002 21888
rect 32030 21836 32036 21888
rect 32088 21876 32094 21888
rect 32582 21876 32588 21888
rect 32088 21848 32588 21876
rect 32088 21836 32094 21848
rect 32582 21836 32588 21848
rect 32640 21836 32646 21888
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32732 21848 33057 21876
rect 32732 21836 32738 21848
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 33410 21836 33416 21888
rect 33468 21836 33474 21888
rect 34330 21836 34336 21888
rect 34388 21836 34394 21888
rect 35250 21836 35256 21888
rect 35308 21836 35314 21888
rect 35621 21879 35679 21885
rect 35621 21845 35633 21879
rect 35667 21876 35679 21879
rect 35986 21876 35992 21888
rect 35667 21848 35992 21876
rect 35667 21845 35679 21848
rect 35621 21839 35679 21845
rect 35986 21836 35992 21848
rect 36044 21836 36050 21888
rect 36262 21836 36268 21888
rect 36320 21876 36326 21888
rect 36357 21879 36415 21885
rect 36357 21876 36369 21879
rect 36320 21848 36369 21876
rect 36320 21836 36326 21848
rect 36357 21845 36369 21848
rect 36403 21845 36415 21879
rect 36357 21839 36415 21845
rect 36814 21836 36820 21888
rect 36872 21836 36878 21888
rect 37366 21836 37372 21888
rect 37424 21836 37430 21888
rect 37476 21876 37504 21916
rect 39132 21876 39160 21984
rect 41506 21972 41512 22024
rect 41564 22012 41570 22024
rect 42518 22012 42524 22024
rect 41564 21984 42524 22012
rect 41564 21972 41570 21984
rect 42518 21972 42524 21984
rect 42576 21972 42582 22024
rect 42797 22015 42855 22021
rect 42797 21981 42809 22015
rect 42843 22012 42855 22015
rect 42978 22012 42984 22024
rect 42843 21984 42984 22012
rect 42843 21981 42855 21984
rect 42797 21975 42855 21981
rect 42978 21972 42984 21984
rect 43036 22012 43042 22024
rect 43714 22012 43720 22024
rect 43036 21984 43720 22012
rect 43036 21972 43042 21984
rect 43714 21972 43720 21984
rect 43772 21972 43778 22024
rect 43806 21972 43812 22024
rect 43864 21972 43870 22024
rect 44082 21972 44088 22024
rect 44140 21972 44146 22024
rect 46017 22015 46075 22021
rect 45020 21984 45232 22012
rect 40604 21916 40816 21944
rect 37476 21848 39160 21876
rect 39574 21836 39580 21888
rect 39632 21876 39638 21888
rect 39850 21876 39856 21888
rect 39632 21848 39856 21876
rect 39632 21836 39638 21848
rect 39850 21836 39856 21848
rect 39908 21836 39914 21888
rect 39942 21836 39948 21888
rect 40000 21876 40006 21888
rect 40604 21885 40632 21916
rect 40589 21879 40647 21885
rect 40589 21876 40601 21879
rect 40000 21848 40601 21876
rect 40000 21836 40006 21848
rect 40589 21845 40601 21848
rect 40635 21845 40647 21879
rect 40788 21876 40816 21916
rect 40954 21904 40960 21956
rect 41012 21944 41018 21956
rect 41785 21947 41843 21953
rect 41012 21916 41736 21944
rect 41012 21904 41018 21916
rect 41506 21876 41512 21888
rect 40788 21848 41512 21876
rect 40589 21839 40647 21845
rect 41506 21836 41512 21848
rect 41564 21836 41570 21888
rect 41708 21876 41736 21916
rect 41785 21913 41797 21947
rect 41831 21944 41843 21947
rect 45020 21944 45048 21984
rect 41831 21916 45048 21944
rect 41831 21913 41843 21916
rect 41785 21907 41843 21913
rect 41877 21879 41935 21885
rect 41877 21876 41889 21879
rect 41708 21848 41889 21876
rect 41877 21845 41889 21848
rect 41923 21876 41935 21879
rect 42150 21876 42156 21888
rect 41923 21848 42156 21876
rect 41923 21845 41935 21848
rect 41877 21839 41935 21845
rect 42150 21836 42156 21848
rect 42208 21836 42214 21888
rect 42242 21836 42248 21888
rect 42300 21876 42306 21888
rect 42613 21879 42671 21885
rect 42613 21876 42625 21879
rect 42300 21848 42625 21876
rect 42300 21836 42306 21848
rect 42613 21845 42625 21848
rect 42659 21845 42671 21879
rect 42613 21839 42671 21845
rect 43254 21836 43260 21888
rect 43312 21876 43318 21888
rect 43349 21879 43407 21885
rect 43349 21876 43361 21879
rect 43312 21848 43361 21876
rect 43312 21836 43318 21848
rect 43349 21845 43361 21848
rect 43395 21876 43407 21879
rect 43533 21879 43591 21885
rect 43533 21876 43545 21879
rect 43395 21848 43545 21876
rect 43395 21845 43407 21848
rect 43349 21839 43407 21845
rect 43533 21845 43545 21848
rect 43579 21876 43591 21879
rect 45094 21876 45100 21888
rect 43579 21848 45100 21876
rect 43579 21845 43591 21848
rect 43533 21839 43591 21845
rect 45094 21836 45100 21848
rect 45152 21836 45158 21888
rect 45204 21876 45232 21984
rect 46017 21981 46029 22015
rect 46063 22012 46075 22015
rect 46106 22012 46112 22024
rect 46063 21984 46112 22012
rect 46063 21981 46075 21984
rect 46017 21975 46075 21981
rect 46106 21972 46112 21984
rect 46164 21972 46170 22024
rect 46569 22015 46627 22021
rect 46569 21981 46581 22015
rect 46615 22012 46627 22015
rect 47213 22015 47271 22021
rect 46615 21984 47164 22012
rect 46615 21981 46627 21984
rect 46569 21975 46627 21981
rect 47136 21944 47164 21984
rect 47213 21981 47225 22015
rect 47259 22012 47271 22015
rect 47486 22012 47492 22024
rect 47259 21984 47492 22012
rect 47259 21981 47271 21984
rect 47213 21975 47271 21981
rect 47486 21972 47492 21984
rect 47544 22012 47550 22024
rect 47673 22015 47731 22021
rect 47673 22012 47685 22015
rect 47544 21984 47685 22012
rect 47544 21972 47550 21984
rect 47673 21981 47685 21984
rect 47719 21981 47731 22015
rect 47673 21975 47731 21981
rect 47578 21944 47584 21956
rect 47136 21916 47584 21944
rect 47578 21904 47584 21916
rect 47636 21904 47642 21956
rect 47854 21904 47860 21956
rect 47912 21944 47918 21956
rect 48225 21947 48283 21953
rect 48225 21944 48237 21947
rect 47912 21916 48237 21944
rect 47912 21904 47918 21916
rect 48225 21913 48237 21916
rect 48271 21913 48283 21947
rect 48225 21907 48283 21913
rect 49234 21904 49240 21956
rect 49292 21904 49298 21956
rect 46385 21879 46443 21885
rect 46385 21876 46397 21879
rect 45204 21848 46397 21876
rect 46385 21845 46397 21848
rect 46431 21845 46443 21879
rect 46385 21839 46443 21845
rect 48774 21836 48780 21888
rect 48832 21836 48838 21888
rect 48866 21836 48872 21888
rect 48924 21876 48930 21888
rect 49145 21879 49203 21885
rect 49145 21876 49157 21879
rect 48924 21848 49157 21876
rect 48924 21836 48930 21848
rect 49145 21845 49157 21848
rect 49191 21845 49203 21879
rect 49145 21839 49203 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 6730 21632 6736 21684
rect 6788 21672 6794 21684
rect 6788 21644 9168 21672
rect 6788 21632 6794 21644
rect 3326 21564 3332 21616
rect 3384 21604 3390 21616
rect 3605 21607 3663 21613
rect 3605 21604 3617 21607
rect 3384 21576 3617 21604
rect 3384 21564 3390 21576
rect 3605 21573 3617 21576
rect 3651 21573 3663 21607
rect 3605 21567 3663 21573
rect 7190 21564 7196 21616
rect 7248 21604 7254 21616
rect 9140 21604 9168 21644
rect 9490 21632 9496 21684
rect 9548 21672 9554 21684
rect 10505 21675 10563 21681
rect 10505 21672 10517 21675
rect 9548 21644 10517 21672
rect 9548 21632 9554 21644
rect 10505 21641 10517 21644
rect 10551 21641 10563 21675
rect 12526 21672 12532 21684
rect 10505 21635 10563 21641
rect 10612 21644 12532 21672
rect 10612 21604 10640 21644
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 13722 21632 13728 21684
rect 13780 21672 13786 21684
rect 13909 21675 13967 21681
rect 13909 21672 13921 21675
rect 13780 21644 13921 21672
rect 13780 21632 13786 21644
rect 13909 21641 13921 21644
rect 13955 21641 13967 21675
rect 13909 21635 13967 21641
rect 14090 21632 14096 21684
rect 14148 21672 14154 21684
rect 16666 21672 16672 21684
rect 14148 21644 16672 21672
rect 14148 21632 14154 21644
rect 7248 21576 8984 21604
rect 9140 21576 10640 21604
rect 7248 21564 7254 21576
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 1762 21428 1768 21480
rect 1820 21428 1826 21480
rect 2976 21468 3004 21499
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21536 5779 21539
rect 6546 21536 6552 21548
rect 5767 21508 6552 21536
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 6546 21496 6552 21508
rect 6604 21496 6610 21548
rect 6638 21496 6644 21548
rect 6696 21496 6702 21548
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21505 8539 21539
rect 8481 21499 8539 21505
rect 5626 21468 5632 21480
rect 2976 21440 5632 21468
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 5810 21428 5816 21480
rect 5868 21468 5874 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 5868 21440 7021 21468
rect 5868 21428 5874 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 5905 21403 5963 21409
rect 5905 21369 5917 21403
rect 5951 21400 5963 21403
rect 8496 21400 8524 21499
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21437 8907 21471
rect 8956 21468 8984 21576
rect 11422 21564 11428 21616
rect 11480 21604 11486 21616
rect 11698 21604 11704 21616
rect 11480 21576 11704 21604
rect 11480 21564 11486 21576
rect 11698 21564 11704 21576
rect 11756 21564 11762 21616
rect 11808 21576 12572 21604
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 9950 21536 9956 21548
rect 9640 21508 9956 21536
rect 9640 21496 9646 21508
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21536 10747 21539
rect 10962 21536 10968 21548
rect 10735 21508 10968 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 11808 21468 11836 21576
rect 12342 21496 12348 21548
rect 12400 21496 12406 21548
rect 12544 21536 12572 21576
rect 12618 21564 12624 21616
rect 12676 21604 12682 21616
rect 13081 21607 13139 21613
rect 13081 21604 13093 21607
rect 12676 21576 13093 21604
rect 12676 21564 12682 21576
rect 13081 21573 13093 21576
rect 13127 21573 13139 21607
rect 14182 21604 14188 21616
rect 13081 21567 13139 21573
rect 13188 21576 14188 21604
rect 13188 21536 13216 21576
rect 14182 21564 14188 21576
rect 14240 21564 14246 21616
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 14829 21607 14887 21613
rect 14829 21604 14841 21607
rect 14332 21576 14841 21604
rect 14332 21564 14338 21576
rect 14829 21573 14841 21576
rect 14875 21573 14887 21607
rect 15212 21604 15240 21644
rect 16666 21632 16672 21644
rect 16724 21672 16730 21684
rect 16853 21675 16911 21681
rect 16853 21672 16865 21675
rect 16724 21644 16865 21672
rect 16724 21632 16730 21644
rect 16853 21641 16865 21644
rect 16899 21641 16911 21675
rect 16853 21635 16911 21641
rect 17402 21632 17408 21684
rect 17460 21632 17466 21684
rect 17862 21632 17868 21684
rect 17920 21632 17926 21684
rect 19794 21672 19800 21684
rect 17972 21644 19800 21672
rect 15286 21604 15292 21616
rect 15212 21576 15292 21604
rect 14829 21567 14887 21573
rect 15286 21564 15292 21576
rect 15344 21564 15350 21616
rect 17218 21564 17224 21616
rect 17276 21604 17282 21616
rect 17972 21604 18000 21644
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 22462 21632 22468 21684
rect 22520 21672 22526 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 22520 21644 24777 21672
rect 22520 21632 22526 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 24765 21635 24823 21641
rect 25774 21632 25780 21684
rect 25832 21672 25838 21684
rect 25961 21675 26019 21681
rect 25961 21672 25973 21675
rect 25832 21644 25973 21672
rect 25832 21632 25838 21644
rect 25961 21641 25973 21644
rect 26007 21641 26019 21675
rect 25961 21635 26019 21641
rect 27157 21675 27215 21681
rect 27157 21641 27169 21675
rect 27203 21641 27215 21675
rect 27157 21635 27215 21641
rect 18782 21604 18788 21616
rect 17276 21576 18000 21604
rect 18432 21576 18788 21604
rect 17276 21564 17282 21576
rect 12544 21508 13216 21536
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 13998 21536 14004 21548
rect 13311 21508 14004 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21536 14151 21539
rect 14366 21536 14372 21548
rect 14139 21508 14372 21536
rect 14139 21505 14151 21508
rect 14093 21499 14151 21505
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 18322 21536 18328 21548
rect 17819 21508 18328 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 8956 21440 11836 21468
rect 8849 21431 8907 21437
rect 5951 21372 8524 21400
rect 5951 21369 5963 21372
rect 5905 21363 5963 21369
rect 3786 21292 3792 21344
rect 3844 21332 3850 21344
rect 8864 21332 8892 21431
rect 12434 21428 12440 21480
rect 12492 21468 12498 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12492 21440 12817 21468
rect 12492 21428 12498 21440
rect 12805 21437 12817 21440
rect 12851 21468 12863 21471
rect 14550 21468 14556 21480
rect 12851 21440 14556 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 14550 21428 14556 21440
rect 14608 21428 14614 21480
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21468 18107 21471
rect 18432 21468 18460 21576
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 20714 21564 20720 21616
rect 20772 21604 20778 21616
rect 21177 21607 21235 21613
rect 21177 21604 21189 21607
rect 20772 21576 21189 21604
rect 20772 21564 20778 21576
rect 21177 21573 21189 21576
rect 21223 21573 21235 21607
rect 21177 21567 21235 21573
rect 23014 21564 23020 21616
rect 23072 21604 23078 21616
rect 23198 21604 23204 21616
rect 23072 21576 23204 21604
rect 23072 21564 23078 21576
rect 23198 21564 23204 21576
rect 23256 21564 23262 21616
rect 24026 21564 24032 21616
rect 24084 21604 24090 21616
rect 27172 21604 27200 21635
rect 27430 21632 27436 21684
rect 27488 21672 27494 21684
rect 27617 21675 27675 21681
rect 27617 21672 27629 21675
rect 27488 21644 27629 21672
rect 27488 21632 27494 21644
rect 27617 21641 27629 21644
rect 27663 21641 27675 21675
rect 27617 21635 27675 21641
rect 27798 21632 27804 21684
rect 27856 21672 27862 21684
rect 28353 21675 28411 21681
rect 28353 21672 28365 21675
rect 27856 21644 28365 21672
rect 27856 21632 27862 21644
rect 28353 21641 28365 21644
rect 28399 21641 28411 21675
rect 28353 21635 28411 21641
rect 28810 21632 28816 21684
rect 28868 21632 28874 21684
rect 30006 21632 30012 21684
rect 30064 21672 30070 21684
rect 31386 21672 31392 21684
rect 30064 21644 31392 21672
rect 30064 21632 30070 21644
rect 31386 21632 31392 21644
rect 31444 21672 31450 21684
rect 31754 21672 31760 21684
rect 31444 21644 31760 21672
rect 31444 21632 31450 21644
rect 31754 21632 31760 21644
rect 31812 21672 31818 21684
rect 32398 21672 32404 21684
rect 31812 21644 32404 21672
rect 31812 21632 31818 21644
rect 32398 21632 32404 21644
rect 32456 21632 32462 21684
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21672 32827 21675
rect 33410 21672 33416 21684
rect 32815 21644 33416 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 33410 21632 33416 21644
rect 33468 21632 33474 21684
rect 33597 21675 33655 21681
rect 33597 21641 33609 21675
rect 33643 21672 33655 21675
rect 34606 21672 34612 21684
rect 33643 21644 34612 21672
rect 33643 21641 33655 21644
rect 33597 21635 33655 21641
rect 24084 21576 27200 21604
rect 27525 21607 27583 21613
rect 24084 21564 24090 21576
rect 27525 21573 27537 21607
rect 27571 21604 27583 21607
rect 29454 21604 29460 21616
rect 27571 21576 29460 21604
rect 27571 21573 27583 21576
rect 27525 21567 27583 21573
rect 29454 21564 29460 21576
rect 29512 21564 29518 21616
rect 30650 21604 30656 21616
rect 29840 21576 30656 21604
rect 20898 21536 20904 21548
rect 20010 21508 20904 21536
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21358 21496 21364 21548
rect 21416 21496 21422 21548
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 25777 21539 25835 21545
rect 25777 21536 25789 21539
rect 25188 21508 25789 21536
rect 25188 21496 25194 21508
rect 25777 21505 25789 21508
rect 25823 21536 25835 21539
rect 26142 21536 26148 21548
rect 25823 21508 26148 21536
rect 25823 21505 25835 21508
rect 25777 21499 25835 21505
rect 26142 21496 26148 21508
rect 26200 21496 26206 21548
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21536 26663 21539
rect 26651 21508 27844 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 18095 21440 18460 21468
rect 18601 21471 18659 21477
rect 18095 21437 18107 21440
rect 18049 21431 18107 21437
rect 18601 21437 18613 21471
rect 18647 21437 18659 21471
rect 18601 21431 18659 21437
rect 11149 21403 11207 21409
rect 11149 21369 11161 21403
rect 11195 21400 11207 21403
rect 11790 21400 11796 21412
rect 11195 21372 11796 21400
rect 11195 21369 11207 21372
rect 11149 21363 11207 21369
rect 11790 21360 11796 21372
rect 11848 21360 11854 21412
rect 11885 21403 11943 21409
rect 11885 21369 11897 21403
rect 11931 21400 11943 21403
rect 11931 21372 12434 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 3844 21304 8892 21332
rect 11333 21335 11391 21341
rect 3844 21292 3850 21304
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11698 21332 11704 21344
rect 11379 21304 11704 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 12250 21292 12256 21344
rect 12308 21292 12314 21344
rect 12406 21332 12434 21372
rect 12802 21332 12808 21344
rect 12406 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 14568 21332 14596 21428
rect 16761 21403 16819 21409
rect 16761 21400 16773 21403
rect 15856 21372 16773 21400
rect 15856 21332 15884 21372
rect 16761 21369 16773 21372
rect 16807 21400 16819 21403
rect 16850 21400 16856 21412
rect 16807 21372 16856 21400
rect 16807 21369 16819 21372
rect 16761 21363 16819 21369
rect 16850 21360 16856 21372
rect 16908 21400 16914 21412
rect 17129 21403 17187 21409
rect 17129 21400 17141 21403
rect 16908 21372 17141 21400
rect 16908 21360 16914 21372
rect 17129 21369 17141 21372
rect 17175 21400 17187 21403
rect 18616 21400 18644 21431
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 19024 21440 22094 21468
rect 19024 21428 19030 21440
rect 17175 21372 18644 21400
rect 17175 21369 17187 21372
rect 17129 21363 17187 21369
rect 14568 21304 15884 21332
rect 16301 21335 16359 21341
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 16574 21332 16580 21344
rect 16347 21304 16580 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 18616 21332 18644 21372
rect 20349 21403 20407 21409
rect 20349 21369 20361 21403
rect 20395 21400 20407 21403
rect 21450 21400 21456 21412
rect 20395 21372 21456 21400
rect 20395 21369 20407 21372
rect 20349 21363 20407 21369
rect 21450 21360 21456 21372
rect 21508 21360 21514 21412
rect 22066 21400 22094 21440
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22244 21440 22477 21468
rect 22244 21428 22250 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22465 21431 22523 21437
rect 22572 21440 22753 21468
rect 22572 21400 22600 21440
rect 22741 21437 22753 21440
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 24210 21428 24216 21480
rect 24268 21468 24274 21480
rect 25225 21471 25283 21477
rect 25225 21468 25237 21471
rect 24268 21440 25237 21468
rect 24268 21428 24274 21440
rect 25225 21437 25237 21440
rect 25271 21468 25283 21471
rect 25314 21468 25320 21480
rect 25271 21440 25320 21468
rect 25271 21437 25283 21440
rect 25225 21431 25283 21437
rect 25314 21428 25320 21440
rect 25372 21428 25378 21480
rect 25406 21428 25412 21480
rect 25464 21468 25470 21480
rect 27709 21471 27767 21477
rect 27709 21468 27721 21471
rect 25464 21440 27721 21468
rect 25464 21428 25470 21440
rect 27709 21437 27721 21440
rect 27755 21437 27767 21471
rect 27816 21468 27844 21508
rect 27890 21496 27896 21548
rect 27948 21536 27954 21548
rect 28721 21539 28779 21545
rect 28721 21536 28733 21539
rect 27948 21508 28733 21536
rect 27948 21496 27954 21508
rect 28721 21505 28733 21508
rect 28767 21505 28779 21539
rect 29840 21536 29868 21576
rect 30650 21564 30656 21576
rect 30708 21564 30714 21616
rect 31202 21564 31208 21616
rect 31260 21564 31266 21616
rect 28721 21499 28779 21505
rect 28828 21508 29868 21536
rect 28828 21468 28856 21508
rect 29914 21496 29920 21548
rect 29972 21496 29978 21548
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 30926 21536 30932 21548
rect 30055 21508 30932 21536
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 30926 21496 30932 21508
rect 30984 21496 30990 21548
rect 31113 21539 31171 21545
rect 31113 21505 31125 21539
rect 31159 21536 31171 21539
rect 31159 21508 31754 21536
rect 31159 21505 31171 21508
rect 31113 21499 31171 21505
rect 27816 21440 28856 21468
rect 27709 21431 27767 21437
rect 28902 21428 28908 21480
rect 28960 21428 28966 21480
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29012 21440 30113 21468
rect 22066 21372 22600 21400
rect 26418 21360 26424 21412
rect 26476 21360 26482 21412
rect 26878 21360 26884 21412
rect 26936 21400 26942 21412
rect 29012 21400 29040 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 30466 21428 30472 21480
rect 30524 21468 30530 21480
rect 31389 21471 31447 21477
rect 31389 21468 31401 21471
rect 30524 21440 31401 21468
rect 30524 21428 30530 21440
rect 31389 21437 31401 21440
rect 31435 21437 31447 21471
rect 31389 21431 31447 21437
rect 26936 21372 29040 21400
rect 26936 21360 26942 21372
rect 29914 21360 29920 21412
rect 29972 21400 29978 21412
rect 31110 21400 31116 21412
rect 29972 21372 31116 21400
rect 29972 21360 29978 21372
rect 31110 21360 31116 21372
rect 31168 21360 31174 21412
rect 19334 21332 19340 21344
rect 18616 21304 19340 21332
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 20717 21335 20775 21341
rect 20717 21301 20729 21335
rect 20763 21332 20775 21335
rect 20898 21332 20904 21344
rect 20763 21304 20904 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 20898 21292 20904 21304
rect 20956 21332 20962 21344
rect 21634 21332 21640 21344
rect 20956 21304 21640 21332
rect 20956 21292 20962 21304
rect 21634 21292 21640 21304
rect 21692 21332 21698 21344
rect 21913 21335 21971 21341
rect 21913 21332 21925 21335
rect 21692 21304 21925 21332
rect 21692 21292 21698 21304
rect 21913 21301 21925 21304
rect 21959 21332 21971 21335
rect 22097 21335 22155 21341
rect 22097 21332 22109 21335
rect 21959 21304 22109 21332
rect 21959 21301 21971 21304
rect 21913 21295 21971 21301
rect 22097 21301 22109 21304
rect 22143 21301 22155 21335
rect 22097 21295 22155 21301
rect 24213 21335 24271 21341
rect 24213 21301 24225 21335
rect 24259 21332 24271 21335
rect 26142 21332 26148 21344
rect 24259 21304 26148 21332
rect 24259 21301 24271 21304
rect 24213 21295 24271 21301
rect 26142 21292 26148 21304
rect 26200 21292 26206 21344
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 26970 21332 26976 21344
rect 26292 21304 26976 21332
rect 26292 21292 26298 21304
rect 26970 21292 26976 21304
rect 27028 21292 27034 21344
rect 29546 21292 29552 21344
rect 29604 21292 29610 21344
rect 30742 21292 30748 21344
rect 30800 21292 30806 21344
rect 31404 21332 31432 21431
rect 31726 21400 31754 21508
rect 31938 21496 31944 21548
rect 31996 21536 32002 21548
rect 33410 21536 33416 21548
rect 31996 21508 33416 21536
rect 31996 21496 32002 21508
rect 33410 21496 33416 21508
rect 33468 21496 33474 21548
rect 33502 21496 33508 21548
rect 33560 21496 33566 21548
rect 33318 21428 33324 21480
rect 33376 21428 33382 21480
rect 34256 21400 34284 21644
rect 34606 21632 34612 21644
rect 34664 21632 34670 21684
rect 34698 21632 34704 21684
rect 34756 21632 34762 21684
rect 34790 21632 34796 21684
rect 34848 21632 34854 21684
rect 35250 21632 35256 21684
rect 35308 21672 35314 21684
rect 36909 21675 36967 21681
rect 36909 21672 36921 21675
rect 35308 21644 36921 21672
rect 35308 21632 35314 21644
rect 36909 21641 36921 21644
rect 36955 21672 36967 21675
rect 37734 21672 37740 21684
rect 36955 21644 37740 21672
rect 36955 21641 36967 21644
rect 36909 21635 36967 21641
rect 37734 21632 37740 21644
rect 37792 21632 37798 21684
rect 38378 21632 38384 21684
rect 38436 21672 38442 21684
rect 38436 21644 39620 21672
rect 38436 21632 38442 21644
rect 36081 21607 36139 21613
rect 36081 21573 36093 21607
rect 36127 21604 36139 21607
rect 38286 21604 38292 21616
rect 36127 21576 38292 21604
rect 36127 21573 36139 21576
rect 36081 21567 36139 21573
rect 38286 21564 38292 21576
rect 38344 21564 38350 21616
rect 38562 21564 38568 21616
rect 38620 21604 38626 21616
rect 38620 21576 38778 21604
rect 38620 21564 38626 21576
rect 36725 21539 36783 21545
rect 36725 21536 36737 21539
rect 34624 21508 36737 21536
rect 34624 21477 34652 21508
rect 36725 21505 36737 21508
rect 36771 21536 36783 21539
rect 36814 21536 36820 21548
rect 36771 21508 36820 21536
rect 36771 21505 36783 21508
rect 36725 21499 36783 21505
rect 36814 21496 36820 21508
rect 36872 21496 36878 21548
rect 36998 21496 37004 21548
rect 37056 21536 37062 21548
rect 37274 21536 37280 21548
rect 37056 21508 37280 21536
rect 37056 21496 37062 21508
rect 37274 21496 37280 21508
rect 37332 21496 37338 21548
rect 39592 21536 39620 21644
rect 39850 21632 39856 21684
rect 39908 21672 39914 21684
rect 40037 21675 40095 21681
rect 40037 21672 40049 21675
rect 39908 21644 40049 21672
rect 39908 21632 39914 21644
rect 40037 21641 40049 21644
rect 40083 21672 40095 21675
rect 40221 21675 40279 21681
rect 40221 21672 40233 21675
rect 40083 21644 40233 21672
rect 40083 21641 40095 21644
rect 40037 21635 40095 21641
rect 40221 21641 40233 21644
rect 40267 21672 40279 21675
rect 40405 21675 40463 21681
rect 40405 21672 40417 21675
rect 40267 21644 40417 21672
rect 40267 21641 40279 21644
rect 40221 21635 40279 21641
rect 40405 21641 40417 21644
rect 40451 21672 40463 21675
rect 40681 21675 40739 21681
rect 40681 21672 40693 21675
rect 40451 21644 40693 21672
rect 40451 21641 40463 21644
rect 40405 21635 40463 21641
rect 40681 21641 40693 21644
rect 40727 21672 40739 21675
rect 42058 21672 42064 21684
rect 40727 21644 42064 21672
rect 40727 21641 40739 21644
rect 40681 21635 40739 21641
rect 42058 21632 42064 21644
rect 42116 21632 42122 21684
rect 42518 21632 42524 21684
rect 42576 21632 42582 21684
rect 43714 21632 43720 21684
rect 43772 21632 43778 21684
rect 44266 21632 44272 21684
rect 44324 21632 44330 21684
rect 44450 21632 44456 21684
rect 44508 21632 44514 21684
rect 45922 21632 45928 21684
rect 45980 21672 45986 21684
rect 47029 21675 47087 21681
rect 47029 21672 47041 21675
rect 45980 21644 47041 21672
rect 45980 21632 45986 21644
rect 47029 21641 47041 21644
rect 47075 21641 47087 21675
rect 47029 21635 47087 21641
rect 47854 21632 47860 21684
rect 47912 21632 47918 21684
rect 40586 21564 40592 21616
rect 40644 21604 40650 21616
rect 40770 21604 40776 21616
rect 40644 21576 40776 21604
rect 40644 21564 40650 21576
rect 40770 21564 40776 21576
rect 40828 21564 40834 21616
rect 40862 21564 40868 21616
rect 40920 21604 40926 21616
rect 40957 21607 41015 21613
rect 40957 21604 40969 21607
rect 40920 21576 40969 21604
rect 40920 21564 40926 21576
rect 40957 21573 40969 21576
rect 41003 21573 41015 21607
rect 40957 21567 41015 21573
rect 46753 21607 46811 21613
rect 46753 21573 46765 21607
rect 46799 21604 46811 21607
rect 47670 21604 47676 21616
rect 46799 21576 47676 21604
rect 46799 21573 46811 21576
rect 46753 21567 46811 21573
rect 47670 21564 47676 21576
rect 47728 21564 47734 21616
rect 43441 21539 43499 21545
rect 43441 21536 43453 21539
rect 39592 21508 43453 21536
rect 43441 21505 43453 21508
rect 43487 21536 43499 21539
rect 43901 21539 43959 21545
rect 43901 21536 43913 21539
rect 43487 21508 43913 21536
rect 43487 21505 43499 21508
rect 43441 21499 43499 21505
rect 43901 21505 43913 21508
rect 43947 21505 43959 21539
rect 43901 21499 43959 21505
rect 47213 21539 47271 21545
rect 47213 21505 47225 21539
rect 47259 21536 47271 21539
rect 47394 21536 47400 21548
rect 47259 21508 47400 21536
rect 47259 21505 47271 21508
rect 47213 21499 47271 21505
rect 47394 21496 47400 21508
rect 47452 21496 47458 21548
rect 47765 21539 47823 21545
rect 47765 21505 47777 21539
rect 47811 21536 47823 21539
rect 48222 21536 48228 21548
rect 47811 21508 48228 21536
rect 47811 21505 47823 21508
rect 47765 21499 47823 21505
rect 48222 21496 48228 21508
rect 48280 21536 48286 21548
rect 48593 21539 48651 21545
rect 48593 21536 48605 21539
rect 48280 21508 48605 21536
rect 48280 21496 48286 21508
rect 48593 21505 48605 21508
rect 48639 21505 48651 21539
rect 48593 21499 48651 21505
rect 49326 21496 49332 21548
rect 49384 21496 49390 21548
rect 34609 21471 34667 21477
rect 34609 21437 34621 21471
rect 34655 21437 34667 21471
rect 34609 21431 34667 21437
rect 36170 21428 36176 21480
rect 36228 21428 36234 21480
rect 36265 21471 36323 21477
rect 36265 21437 36277 21471
rect 36311 21437 36323 21471
rect 36265 21431 36323 21437
rect 31726 21372 34284 21400
rect 34422 21360 34428 21412
rect 34480 21400 34486 21412
rect 36280 21400 36308 21431
rect 36446 21428 36452 21480
rect 36504 21468 36510 21480
rect 36906 21468 36912 21480
rect 36504 21440 36912 21468
rect 36504 21428 36510 21440
rect 36906 21428 36912 21440
rect 36964 21428 36970 21480
rect 37550 21428 37556 21480
rect 37608 21468 37614 21480
rect 38013 21471 38071 21477
rect 38013 21468 38025 21471
rect 37608 21440 38025 21468
rect 37608 21428 37614 21440
rect 38013 21437 38025 21440
rect 38059 21437 38071 21471
rect 38286 21468 38292 21480
rect 38013 21431 38071 21437
rect 38120 21440 38292 21468
rect 34480 21372 36308 21400
rect 34480 21360 34486 21372
rect 37366 21360 37372 21412
rect 37424 21400 37430 21412
rect 38120 21400 38148 21440
rect 38286 21428 38292 21440
rect 38344 21428 38350 21480
rect 38378 21428 38384 21480
rect 38436 21468 38442 21480
rect 40034 21468 40040 21480
rect 38436 21440 40040 21468
rect 38436 21428 38442 21440
rect 40034 21428 40040 21440
rect 40092 21428 40098 21480
rect 40862 21428 40868 21480
rect 40920 21468 40926 21480
rect 41233 21471 41291 21477
rect 41233 21468 41245 21471
rect 40920 21440 41245 21468
rect 40920 21428 40926 21440
rect 41233 21437 41245 21440
rect 41279 21437 41291 21471
rect 41233 21431 41291 21437
rect 41506 21428 41512 21480
rect 41564 21428 41570 21480
rect 41874 21428 41880 21480
rect 41932 21468 41938 21480
rect 43806 21468 43812 21480
rect 41932 21440 43812 21468
rect 41932 21428 41938 21440
rect 43806 21428 43812 21440
rect 43864 21468 43870 21480
rect 44085 21471 44143 21477
rect 44085 21468 44097 21471
rect 43864 21440 44097 21468
rect 43864 21428 43870 21440
rect 44085 21437 44097 21440
rect 44131 21437 44143 21471
rect 44085 21431 44143 21437
rect 46106 21428 46112 21480
rect 46164 21468 46170 21480
rect 49234 21468 49240 21480
rect 46164 21440 49240 21468
rect 46164 21428 46170 21440
rect 49234 21428 49240 21440
rect 49292 21428 49298 21480
rect 37424 21372 38148 21400
rect 37424 21360 37430 21372
rect 39298 21360 39304 21412
rect 39356 21400 39362 21412
rect 40954 21400 40960 21412
rect 39356 21372 40960 21400
rect 39356 21360 39362 21372
rect 40954 21360 40960 21372
rect 41012 21360 41018 21412
rect 42705 21403 42763 21409
rect 42705 21400 42717 21403
rect 41064 21372 42717 21400
rect 31757 21335 31815 21341
rect 31757 21332 31769 21335
rect 31404 21304 31769 21332
rect 31757 21301 31769 21304
rect 31803 21301 31815 21335
rect 31757 21295 31815 21301
rect 33962 21292 33968 21344
rect 34020 21292 34026 21344
rect 35161 21335 35219 21341
rect 35161 21301 35173 21335
rect 35207 21332 35219 21335
rect 35618 21332 35624 21344
rect 35207 21304 35624 21332
rect 35207 21301 35219 21304
rect 35161 21295 35219 21301
rect 35618 21292 35624 21304
rect 35676 21292 35682 21344
rect 35710 21292 35716 21344
rect 35768 21292 35774 21344
rect 37550 21292 37556 21344
rect 37608 21332 37614 21344
rect 37645 21335 37703 21341
rect 37645 21332 37657 21335
rect 37608 21304 37657 21332
rect 37608 21292 37614 21304
rect 37645 21301 37657 21304
rect 37691 21301 37703 21335
rect 37645 21295 37703 21301
rect 37826 21292 37832 21344
rect 37884 21332 37890 21344
rect 39761 21335 39819 21341
rect 39761 21332 39773 21335
rect 37884 21304 39773 21332
rect 37884 21292 37890 21304
rect 39761 21301 39773 21304
rect 39807 21301 39819 21335
rect 39761 21295 39819 21301
rect 40862 21292 40868 21344
rect 40920 21332 40926 21344
rect 41064 21332 41092 21372
rect 42705 21369 42717 21372
rect 42751 21400 42763 21403
rect 48409 21403 48467 21409
rect 48409 21400 48421 21403
rect 42751 21372 48421 21400
rect 42751 21369 42763 21372
rect 42705 21363 42763 21369
rect 48409 21369 48421 21372
rect 48455 21369 48467 21403
rect 48409 21363 48467 21369
rect 40920 21304 41092 21332
rect 40920 21292 40926 21304
rect 41414 21292 41420 21344
rect 41472 21332 41478 21344
rect 42797 21335 42855 21341
rect 42797 21332 42809 21335
rect 41472 21304 42809 21332
rect 41472 21292 41478 21304
rect 42797 21301 42809 21304
rect 42843 21301 42855 21335
rect 42797 21295 42855 21301
rect 43257 21335 43315 21341
rect 43257 21301 43269 21335
rect 43303 21332 43315 21335
rect 43438 21332 43444 21344
rect 43303 21304 43444 21332
rect 43303 21301 43315 21304
rect 43257 21295 43315 21301
rect 43438 21292 43444 21304
rect 43496 21292 43502 21344
rect 48314 21292 48320 21344
rect 48372 21332 48378 21344
rect 49145 21335 49203 21341
rect 49145 21332 49157 21335
rect 48372 21304 49157 21332
rect 48372 21292 48378 21304
rect 49145 21301 49157 21304
rect 49191 21301 49203 21335
rect 49145 21295 49203 21301
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 7190 21088 7196 21140
rect 7248 21128 7254 21140
rect 7469 21131 7527 21137
rect 7469 21128 7481 21131
rect 7248 21100 7481 21128
rect 7248 21088 7254 21100
rect 7469 21097 7481 21100
rect 7515 21097 7527 21131
rect 7469 21091 7527 21097
rect 9214 21088 9220 21140
rect 9272 21088 9278 21140
rect 12250 21128 12256 21140
rect 9324 21100 12256 21128
rect 9324 21060 9352 21100
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 12434 21088 12440 21140
rect 12492 21088 12498 21140
rect 13354 21128 13360 21140
rect 12636 21100 13360 21128
rect 12636 21060 12664 21100
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 14274 21088 14280 21140
rect 14332 21088 14338 21140
rect 14366 21088 14372 21140
rect 14424 21128 14430 21140
rect 15746 21128 15752 21140
rect 14424 21100 15752 21128
rect 14424 21088 14430 21100
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 17129 21131 17187 21137
rect 17129 21128 17141 21131
rect 16356 21100 17141 21128
rect 16356 21088 16362 21100
rect 17129 21097 17141 21100
rect 17175 21128 17187 21131
rect 19702 21128 19708 21140
rect 17175 21100 19708 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 24029 21131 24087 21137
rect 19852 21100 23428 21128
rect 19852 21088 19858 21100
rect 5368 21032 9352 21060
rect 10060 21032 12664 21060
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 2866 20992 2872 21004
rect 2547 20964 2872 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 4154 20952 4160 21004
rect 4212 20952 4218 21004
rect 5368 20933 5396 21032
rect 5994 20952 6000 21004
rect 6052 20952 6058 21004
rect 9582 20992 9588 21004
rect 7116 20964 9588 20992
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20893 3019 20927
rect 2961 20887 3019 20893
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 2976 20856 3004 20887
rect 7116 20856 7144 20964
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 10060 21001 10088 21032
rect 12710 21020 12716 21072
rect 12768 21020 12774 21072
rect 13541 21063 13599 21069
rect 13541 21029 13553 21063
rect 13587 21029 13599 21063
rect 13541 21023 13599 21029
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20961 10103 20995
rect 10045 20955 10103 20961
rect 10689 20995 10747 21001
rect 10689 20961 10701 20995
rect 10735 20992 10747 20995
rect 13446 20992 13452 21004
rect 10735 20964 13452 20992
rect 10735 20961 10747 20964
rect 10689 20955 10747 20961
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 7193 20927 7251 20933
rect 7193 20893 7205 20927
rect 7239 20924 7251 20927
rect 8021 20927 8079 20933
rect 7239 20896 7880 20924
rect 7239 20893 7251 20896
rect 7193 20887 7251 20893
rect 2976 20828 7144 20856
rect 7852 20797 7880 20896
rect 8021 20893 8033 20927
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20757 7895 20791
rect 8036 20788 8064 20887
rect 8386 20884 8392 20936
rect 8444 20884 8450 20936
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20924 9459 20927
rect 11054 20924 11060 20936
rect 9447 20896 11060 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 11330 20884 11336 20936
rect 11388 20884 11394 20936
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11848 20896 11989 20924
rect 11848 20884 11854 20896
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 8536 20828 11928 20856
rect 8536 20816 8542 20828
rect 10870 20788 10876 20800
rect 8036 20760 10876 20788
rect 7837 20751 7895 20757
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 11146 20748 11152 20800
rect 11204 20748 11210 20800
rect 11900 20797 11928 20828
rect 11885 20791 11943 20797
rect 11885 20757 11897 20791
rect 11931 20757 11943 20791
rect 11992 20788 12020 20887
rect 12066 20884 12072 20936
rect 12124 20924 12130 20936
rect 13556 20924 13584 21023
rect 16666 21020 16672 21072
rect 16724 21060 16730 21072
rect 17494 21060 17500 21072
rect 16724 21032 17500 21060
rect 16724 21020 16730 21032
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 19058 21020 19064 21072
rect 19116 21060 19122 21072
rect 23400 21069 23428 21100
rect 24029 21097 24041 21131
rect 24075 21128 24087 21131
rect 24118 21128 24124 21140
rect 24075 21100 24124 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 24118 21088 24124 21100
rect 24176 21088 24182 21140
rect 26050 21088 26056 21140
rect 26108 21128 26114 21140
rect 26881 21131 26939 21137
rect 26881 21128 26893 21131
rect 26108 21100 26893 21128
rect 26108 21088 26114 21100
rect 26881 21097 26893 21100
rect 26927 21097 26939 21131
rect 26881 21091 26939 21097
rect 29638 21088 29644 21140
rect 29696 21128 29702 21140
rect 29733 21131 29791 21137
rect 29733 21128 29745 21131
rect 29696 21100 29745 21128
rect 29696 21088 29702 21100
rect 29733 21097 29745 21100
rect 29779 21097 29791 21131
rect 29733 21091 29791 21097
rect 30006 21088 30012 21140
rect 30064 21128 30070 21140
rect 30193 21131 30251 21137
rect 30193 21128 30205 21131
rect 30064 21100 30205 21128
rect 30064 21088 30070 21100
rect 30193 21097 30205 21100
rect 30239 21097 30251 21131
rect 35710 21128 35716 21140
rect 30193 21091 30251 21097
rect 31312 21100 35716 21128
rect 19337 21063 19395 21069
rect 19337 21060 19349 21063
rect 19116 21032 19349 21060
rect 19116 21020 19122 21032
rect 19337 21029 19349 21032
rect 19383 21029 19395 21063
rect 19337 21023 19395 21029
rect 19981 21063 20039 21069
rect 19981 21029 19993 21063
rect 20027 21029 20039 21063
rect 21177 21063 21235 21069
rect 21177 21060 21189 21063
rect 19981 21023 20039 21029
rect 20548 21032 21189 21060
rect 19996 20992 20024 21023
rect 20548 21001 20576 21032
rect 21177 21029 21189 21032
rect 21223 21029 21235 21063
rect 21177 21023 21235 21029
rect 23385 21063 23443 21069
rect 23385 21029 23397 21063
rect 23431 21029 23443 21063
rect 23385 21023 23443 21029
rect 23934 21020 23940 21072
rect 23992 21060 23998 21072
rect 25685 21063 25743 21069
rect 25685 21060 25697 21063
rect 23992 21032 25697 21060
rect 23992 21020 23998 21032
rect 25685 21029 25697 21032
rect 25731 21029 25743 21063
rect 25685 21023 25743 21029
rect 26510 21020 26516 21072
rect 26568 21060 26574 21072
rect 29546 21060 29552 21072
rect 26568 21032 29552 21060
rect 26568 21020 26574 21032
rect 29546 21020 29552 21032
rect 29604 21020 29610 21072
rect 29822 21020 29828 21072
rect 29880 21060 29886 21072
rect 30377 21063 30435 21069
rect 30377 21060 30389 21063
rect 29880 21032 30389 21060
rect 29880 21020 29886 21032
rect 30377 21029 30389 21032
rect 30423 21029 30435 21063
rect 30377 21023 30435 21029
rect 20533 20995 20591 21001
rect 20533 20992 20545 20995
rect 13740 20964 20024 20992
rect 20272 20964 20545 20992
rect 13740 20933 13768 20964
rect 12124 20896 13584 20924
rect 13725 20927 13783 20933
rect 12124 20884 12130 20896
rect 13725 20893 13737 20927
rect 13771 20893 13783 20927
rect 13725 20887 13783 20893
rect 16025 20927 16083 20933
rect 16025 20893 16037 20927
rect 16071 20924 16083 20927
rect 16850 20924 16856 20936
rect 16071 20896 16856 20924
rect 16071 20893 16083 20896
rect 16025 20887 16083 20893
rect 16850 20884 16856 20896
rect 16908 20884 16914 20936
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20924 18935 20927
rect 19334 20924 19340 20936
rect 18923 20896 19340 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 19334 20884 19340 20896
rect 19392 20924 19398 20936
rect 19392 20896 19564 20924
rect 19392 20884 19398 20896
rect 12618 20816 12624 20868
rect 12676 20856 12682 20868
rect 12897 20859 12955 20865
rect 12897 20856 12909 20859
rect 12676 20828 12909 20856
rect 12676 20816 12682 20828
rect 12897 20825 12909 20828
rect 12943 20825 12955 20859
rect 12897 20819 12955 20825
rect 13170 20816 13176 20868
rect 13228 20856 13234 20868
rect 14090 20856 14096 20868
rect 13228 20828 14096 20856
rect 13228 20816 13234 20828
rect 14090 20816 14096 20828
rect 14148 20856 14154 20868
rect 15749 20859 15807 20865
rect 14148 20828 14582 20856
rect 14148 20816 14154 20828
rect 15749 20825 15761 20859
rect 15795 20856 15807 20859
rect 16114 20856 16120 20868
rect 15795 20828 16120 20856
rect 15795 20825 15807 20828
rect 15749 20819 15807 20825
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 16669 20859 16727 20865
rect 16669 20825 16681 20859
rect 16715 20856 16727 20859
rect 18601 20859 18659 20865
rect 16715 20828 17356 20856
rect 16715 20825 16727 20828
rect 16669 20819 16727 20825
rect 13814 20788 13820 20800
rect 11992 20760 13820 20788
rect 11885 20751 11943 20757
rect 13814 20748 13820 20760
rect 13872 20748 13878 20800
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 16758 20788 16764 20800
rect 13964 20760 16764 20788
rect 13964 20748 13970 20760
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 17328 20788 17356 20828
rect 18601 20825 18613 20859
rect 18647 20856 18659 20859
rect 19426 20856 19432 20868
rect 18647 20828 19432 20856
rect 18647 20825 18659 20828
rect 18601 20819 18659 20825
rect 19426 20816 19432 20828
rect 19484 20816 19490 20868
rect 18506 20788 18512 20800
rect 17328 20760 18512 20788
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 19536 20797 19564 20896
rect 19794 20884 19800 20936
rect 19852 20924 19858 20936
rect 20272 20924 20300 20964
rect 20533 20961 20545 20964
rect 20579 20961 20591 20995
rect 22554 20992 22560 21004
rect 20533 20955 20591 20961
rect 21192 20964 22560 20992
rect 19852 20896 20300 20924
rect 20349 20927 20407 20933
rect 19852 20884 19858 20896
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 21192 20924 21220 20964
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 22646 20952 22652 21004
rect 22704 20952 22710 21004
rect 23290 20952 23296 21004
rect 23348 20992 23354 21004
rect 24210 20992 24216 21004
rect 23348 20964 24216 20992
rect 23348 20952 23354 20964
rect 24210 20952 24216 20964
rect 24268 20992 24274 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 24268 20964 25145 20992
rect 24268 20952 24274 20964
rect 25133 20961 25145 20964
rect 25179 20992 25191 20995
rect 25317 20995 25375 21001
rect 25317 20992 25329 20995
rect 25179 20964 25329 20992
rect 25179 20961 25191 20964
rect 25133 20955 25191 20961
rect 25317 20961 25329 20964
rect 25363 20961 25375 20995
rect 25317 20955 25375 20961
rect 25590 20952 25596 21004
rect 25648 20992 25654 21004
rect 26237 20995 26295 21001
rect 26237 20992 26249 20995
rect 25648 20964 26249 20992
rect 25648 20952 25654 20964
rect 26237 20961 26249 20964
rect 26283 20961 26295 20995
rect 26237 20955 26295 20961
rect 26326 20952 26332 21004
rect 26384 20992 26390 21004
rect 26384 20964 27568 20992
rect 26384 20952 26390 20964
rect 20395 20896 21220 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 22922 20884 22928 20936
rect 22980 20884 22986 20936
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24176 20896 24593 20924
rect 24176 20884 24182 20896
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 27430 20884 27436 20936
rect 27488 20884 27494 20936
rect 27540 20924 27568 20964
rect 27890 20952 27896 21004
rect 27948 20952 27954 21004
rect 31312 21001 31340 21100
rect 35710 21088 35716 21100
rect 35768 21088 35774 21140
rect 36630 21088 36636 21140
rect 36688 21128 36694 21140
rect 40037 21131 40095 21137
rect 36688 21100 39988 21128
rect 36688 21088 36694 21100
rect 34238 21020 34244 21072
rect 34296 21020 34302 21072
rect 39960 21060 39988 21100
rect 40037 21097 40049 21131
rect 40083 21128 40095 21131
rect 40310 21128 40316 21140
rect 40083 21100 40316 21128
rect 40083 21097 40095 21100
rect 40037 21091 40095 21097
rect 40310 21088 40316 21100
rect 40368 21088 40374 21140
rect 42242 21128 42248 21140
rect 40420 21100 42248 21128
rect 40420 21060 40448 21100
rect 42242 21088 42248 21100
rect 42300 21088 42306 21140
rect 42521 21131 42579 21137
rect 42521 21097 42533 21131
rect 42567 21128 42579 21131
rect 42794 21128 42800 21140
rect 42567 21100 42800 21128
rect 42567 21097 42579 21100
rect 42521 21091 42579 21097
rect 42794 21088 42800 21100
rect 42852 21088 42858 21140
rect 42889 21131 42947 21137
rect 42889 21097 42901 21131
rect 42935 21128 42947 21131
rect 43346 21128 43352 21140
rect 42935 21100 43352 21128
rect 42935 21097 42947 21100
rect 42889 21091 42947 21097
rect 43346 21088 43352 21100
rect 43404 21088 43410 21140
rect 47305 21131 47363 21137
rect 47305 21097 47317 21131
rect 47351 21128 47363 21131
rect 47762 21128 47768 21140
rect 47351 21100 47768 21128
rect 47351 21097 47363 21100
rect 47305 21091 47363 21097
rect 47762 21088 47768 21100
rect 47820 21088 47826 21140
rect 49145 21131 49203 21137
rect 49145 21128 49157 21131
rect 48286 21100 49157 21128
rect 39960 21032 40448 21060
rect 40678 21020 40684 21072
rect 40736 21060 40742 21072
rect 42613 21063 42671 21069
rect 42613 21060 42625 21063
rect 40736 21032 42625 21060
rect 40736 21020 40742 21032
rect 42613 21029 42625 21032
rect 42659 21029 42671 21063
rect 42613 21023 42671 21029
rect 42702 21020 42708 21072
rect 42760 21060 42766 21072
rect 48286 21060 48314 21100
rect 49145 21097 49157 21100
rect 49191 21097 49203 21131
rect 49145 21091 49203 21097
rect 42760 21032 48314 21060
rect 48409 21063 48467 21069
rect 42760 21020 42766 21032
rect 48409 21029 48421 21063
rect 48455 21029 48467 21063
rect 48409 21023 48467 21029
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20992 28595 20995
rect 31297 20995 31355 21001
rect 28583 20964 30144 20992
rect 28583 20961 28595 20964
rect 28537 20955 28595 20961
rect 29546 20924 29552 20936
rect 27540 20896 29552 20924
rect 29546 20884 29552 20896
rect 29604 20884 29610 20936
rect 29914 20884 29920 20936
rect 29972 20884 29978 20936
rect 30116 20924 30144 20964
rect 31297 20961 31309 20995
rect 31343 20961 31355 20995
rect 31297 20955 31355 20961
rect 31481 20995 31539 21001
rect 31481 20961 31493 20995
rect 31527 20992 31539 20995
rect 32306 20992 32312 21004
rect 31527 20964 32312 20992
rect 31527 20961 31539 20964
rect 31481 20955 31539 20961
rect 32306 20952 32312 20964
rect 32364 20992 32370 21004
rect 32769 20995 32827 21001
rect 32769 20992 32781 20995
rect 32364 20964 32781 20992
rect 32364 20952 32370 20964
rect 32769 20961 32781 20964
rect 32815 20961 32827 20995
rect 32769 20955 32827 20961
rect 32858 20952 32864 21004
rect 32916 20992 32922 21004
rect 34256 20992 34284 21020
rect 32916 20964 34284 20992
rect 32916 20952 32922 20964
rect 34330 20952 34336 21004
rect 34388 20992 34394 21004
rect 37093 20995 37151 21001
rect 34388 20964 36676 20992
rect 34388 20952 34394 20964
rect 32030 20924 32036 20936
rect 30116 20896 32036 20924
rect 32030 20884 32036 20896
rect 32088 20884 32094 20936
rect 32490 20884 32496 20936
rect 32548 20884 32554 20936
rect 34514 20884 34520 20936
rect 34572 20924 34578 20936
rect 35066 20924 35072 20936
rect 34572 20896 35072 20924
rect 34572 20884 34578 20896
rect 35066 20884 35072 20896
rect 35124 20924 35130 20936
rect 36648 20933 36676 20964
rect 37093 20961 37105 20995
rect 37139 20992 37151 20995
rect 37550 20992 37556 21004
rect 37139 20964 37556 20992
rect 37139 20961 37151 20964
rect 37093 20955 37151 20961
rect 36633 20927 36691 20933
rect 35124 20896 35282 20924
rect 35124 20884 35130 20896
rect 36633 20893 36645 20927
rect 36679 20924 36691 20927
rect 37108 20924 37136 20955
rect 37550 20952 37556 20964
rect 37608 20992 37614 21004
rect 39393 20995 39451 21001
rect 39393 20992 39405 20995
rect 37608 20964 39405 20992
rect 37608 20952 37614 20964
rect 39393 20961 39405 20964
rect 39439 20992 39451 20995
rect 39482 20992 39488 21004
rect 39439 20964 39488 20992
rect 39439 20961 39451 20964
rect 39393 20955 39451 20961
rect 39482 20952 39488 20964
rect 39540 20952 39546 21004
rect 39666 20952 39672 21004
rect 39724 20992 39730 21004
rect 40497 20995 40555 21001
rect 40497 20992 40509 20995
rect 39724 20964 40509 20992
rect 39724 20952 39730 20964
rect 40497 20961 40509 20964
rect 40543 20961 40555 20995
rect 40497 20955 40555 20961
rect 40589 20995 40647 21001
rect 40589 20961 40601 20995
rect 40635 20961 40647 20995
rect 40589 20955 40647 20961
rect 41785 20995 41843 21001
rect 41785 20961 41797 20995
rect 41831 20961 41843 20995
rect 41785 20955 41843 20961
rect 40604 20924 40632 20955
rect 36679 20896 37136 20924
rect 40328 20896 40632 20924
rect 36679 20893 36691 20896
rect 36633 20887 36691 20893
rect 21358 20816 21364 20868
rect 21416 20856 21422 20868
rect 21416 20828 21482 20856
rect 21416 20816 21422 20828
rect 23566 20816 23572 20868
rect 23624 20816 23630 20868
rect 25222 20856 25228 20868
rect 23676 20828 25228 20856
rect 19521 20791 19579 20797
rect 19521 20757 19533 20791
rect 19567 20788 19579 20791
rect 19610 20788 19616 20800
rect 19567 20760 19616 20788
rect 19567 20757 19579 20760
rect 19521 20751 19579 20757
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 20441 20791 20499 20797
rect 20441 20757 20453 20791
rect 20487 20788 20499 20791
rect 23676 20788 23704 20828
rect 25222 20816 25228 20828
rect 25280 20816 25286 20868
rect 26786 20856 26792 20868
rect 26068 20828 26792 20856
rect 20487 20760 23704 20788
rect 24765 20791 24823 20797
rect 20487 20757 20499 20760
rect 20441 20751 20499 20757
rect 24765 20757 24777 20791
rect 24811 20788 24823 20791
rect 25774 20788 25780 20800
rect 24811 20760 25780 20788
rect 24811 20757 24823 20760
rect 24765 20751 24823 20757
rect 25774 20748 25780 20760
rect 25832 20748 25838 20800
rect 26068 20797 26096 20828
rect 26786 20816 26792 20828
rect 26844 20816 26850 20868
rect 27706 20816 27712 20868
rect 27764 20856 27770 20868
rect 27764 20828 30880 20856
rect 27764 20816 27770 20828
rect 26053 20791 26111 20797
rect 26053 20757 26065 20791
rect 26099 20757 26111 20791
rect 26053 20751 26111 20757
rect 26145 20791 26203 20797
rect 26145 20757 26157 20791
rect 26191 20788 26203 20791
rect 26510 20788 26516 20800
rect 26191 20760 26516 20788
rect 26191 20757 26203 20760
rect 26145 20751 26203 20757
rect 26510 20748 26516 20760
rect 26568 20748 26574 20800
rect 26697 20791 26755 20797
rect 26697 20757 26709 20791
rect 26743 20788 26755 20791
rect 26970 20788 26976 20800
rect 26743 20760 26976 20788
rect 26743 20757 26755 20760
rect 26697 20751 26755 20757
rect 26970 20748 26976 20760
rect 27028 20748 27034 20800
rect 27062 20748 27068 20800
rect 27120 20788 27126 20800
rect 28629 20791 28687 20797
rect 28629 20788 28641 20791
rect 27120 20760 28641 20788
rect 27120 20748 27126 20760
rect 28629 20757 28641 20760
rect 28675 20757 28687 20791
rect 28629 20751 28687 20757
rect 28718 20748 28724 20800
rect 28776 20748 28782 20800
rect 29089 20791 29147 20797
rect 29089 20757 29101 20791
rect 29135 20788 29147 20791
rect 30098 20788 30104 20800
rect 29135 20760 30104 20788
rect 29135 20757 29147 20760
rect 29089 20751 29147 20757
rect 30098 20748 30104 20760
rect 30156 20748 30162 20800
rect 30852 20797 30880 20828
rect 30926 20816 30932 20868
rect 30984 20856 30990 20868
rect 31754 20856 31760 20868
rect 30984 20828 31760 20856
rect 30984 20816 30990 20828
rect 31754 20816 31760 20828
rect 31812 20816 31818 20868
rect 32398 20816 32404 20868
rect 32456 20856 32462 20868
rect 36357 20859 36415 20865
rect 32456 20828 33258 20856
rect 34348 20828 35020 20856
rect 32456 20816 32462 20828
rect 30837 20791 30895 20797
rect 30837 20757 30849 20791
rect 30883 20757 30895 20791
rect 30837 20751 30895 20757
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 31294 20748 31300 20800
rect 31352 20788 31358 20800
rect 31941 20791 31999 20797
rect 31941 20788 31953 20791
rect 31352 20760 31953 20788
rect 31352 20748 31358 20760
rect 31941 20757 31953 20760
rect 31987 20788 31999 20791
rect 34348 20788 34376 20828
rect 31987 20760 34376 20788
rect 31987 20757 31999 20760
rect 31941 20751 31999 20757
rect 34422 20748 34428 20800
rect 34480 20788 34486 20800
rect 34885 20791 34943 20797
rect 34885 20788 34897 20791
rect 34480 20760 34897 20788
rect 34480 20748 34486 20760
rect 34885 20757 34897 20760
rect 34931 20757 34943 20791
rect 34992 20788 35020 20828
rect 36357 20825 36369 20859
rect 36403 20856 36415 20859
rect 36446 20856 36452 20868
rect 36403 20828 36452 20856
rect 36403 20825 36415 20828
rect 36357 20819 36415 20825
rect 36446 20816 36452 20828
rect 36504 20816 36510 20868
rect 36722 20816 36728 20868
rect 36780 20856 36786 20868
rect 37277 20859 37335 20865
rect 37277 20856 37289 20859
rect 36780 20828 37289 20856
rect 36780 20816 36786 20828
rect 37277 20825 37289 20828
rect 37323 20825 37335 20859
rect 37277 20819 37335 20825
rect 38378 20816 38384 20868
rect 38436 20816 38442 20868
rect 39117 20859 39175 20865
rect 39117 20825 39129 20859
rect 39163 20856 39175 20859
rect 40328 20856 40356 20896
rect 40678 20884 40684 20936
rect 40736 20924 40742 20936
rect 41322 20924 41328 20936
rect 40736 20896 41328 20924
rect 40736 20884 40742 20896
rect 41322 20884 41328 20896
rect 41380 20924 41386 20936
rect 41380 20884 41414 20924
rect 41598 20884 41604 20936
rect 41656 20924 41662 20936
rect 41800 20924 41828 20955
rect 41966 20952 41972 21004
rect 42024 20992 42030 21004
rect 48424 20992 48452 21023
rect 42024 20964 48452 20992
rect 42024 20952 42030 20964
rect 41656 20896 41828 20924
rect 41656 20884 41662 20896
rect 47118 20884 47124 20936
rect 47176 20924 47182 20936
rect 47854 20924 47860 20936
rect 47176 20896 47860 20924
rect 47176 20884 47182 20896
rect 47854 20884 47860 20896
rect 47912 20924 47918 20936
rect 47949 20927 48007 20933
rect 47949 20924 47961 20927
rect 47912 20896 47961 20924
rect 47912 20884 47918 20896
rect 47949 20893 47961 20896
rect 47995 20893 48007 20927
rect 47949 20887 48007 20893
rect 48593 20927 48651 20933
rect 48593 20893 48605 20927
rect 48639 20924 48651 20927
rect 48774 20924 48780 20936
rect 48639 20896 48780 20924
rect 48639 20893 48651 20896
rect 48593 20887 48651 20893
rect 48774 20884 48780 20896
rect 48832 20884 48838 20936
rect 49326 20884 49332 20936
rect 49384 20884 49390 20936
rect 39163 20828 40356 20856
rect 40405 20859 40463 20865
rect 39163 20825 39175 20828
rect 39117 20819 39175 20825
rect 40405 20825 40417 20859
rect 40451 20856 40463 20859
rect 41386 20856 41414 20884
rect 41693 20859 41751 20865
rect 41693 20856 41705 20859
rect 40451 20828 41276 20856
rect 41386 20828 41705 20856
rect 40451 20825 40463 20828
rect 40405 20819 40463 20825
rect 36630 20788 36636 20800
rect 34992 20760 36636 20788
rect 34885 20751 34943 20757
rect 36630 20748 36636 20760
rect 36688 20748 36694 20800
rect 36906 20748 36912 20800
rect 36964 20748 36970 20800
rect 37182 20748 37188 20800
rect 37240 20788 37246 20800
rect 37642 20788 37648 20800
rect 37240 20760 37648 20788
rect 37240 20748 37246 20760
rect 37642 20748 37648 20760
rect 37700 20748 37706 20800
rect 37826 20748 37832 20800
rect 37884 20788 37890 20800
rect 39132 20788 39160 20819
rect 37884 20760 39160 20788
rect 37884 20748 37890 20760
rect 40218 20748 40224 20800
rect 40276 20788 40282 20800
rect 40862 20788 40868 20800
rect 40276 20760 40868 20788
rect 40276 20748 40282 20760
rect 40862 20748 40868 20760
rect 40920 20748 40926 20800
rect 41248 20797 41276 20828
rect 41693 20825 41705 20828
rect 41739 20856 41751 20859
rect 41782 20856 41788 20868
rect 41739 20828 41788 20856
rect 41739 20825 41751 20828
rect 41693 20819 41751 20825
rect 41782 20816 41788 20828
rect 41840 20816 41846 20868
rect 42058 20816 42064 20868
rect 42116 20856 42122 20868
rect 42337 20859 42395 20865
rect 42337 20856 42349 20859
rect 42116 20828 42349 20856
rect 42116 20816 42122 20828
rect 42337 20825 42349 20828
rect 42383 20856 42395 20859
rect 46014 20856 46020 20868
rect 42383 20828 46020 20856
rect 42383 20825 42395 20828
rect 42337 20819 42395 20825
rect 46014 20816 46020 20828
rect 46072 20816 46078 20868
rect 47489 20859 47547 20865
rect 47489 20825 47501 20859
rect 47535 20856 47547 20859
rect 49344 20856 49372 20884
rect 47535 20828 49372 20856
rect 47535 20825 47547 20828
rect 47489 20819 47547 20825
rect 41233 20791 41291 20797
rect 41233 20757 41245 20791
rect 41279 20757 41291 20791
rect 41233 20751 41291 20757
rect 41598 20748 41604 20800
rect 41656 20748 41662 20800
rect 43622 20748 43628 20800
rect 43680 20788 43686 20800
rect 47765 20791 47823 20797
rect 47765 20788 47777 20791
rect 43680 20760 47777 20788
rect 43680 20748 43686 20760
rect 47765 20757 47777 20760
rect 47811 20757 47823 20791
rect 47765 20751 47823 20757
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5445 20587 5503 20593
rect 5445 20553 5457 20587
rect 5491 20584 5503 20587
rect 6638 20584 6644 20596
rect 5491 20556 6644 20584
rect 5491 20553 5503 20556
rect 5445 20547 5503 20553
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 13725 20587 13783 20593
rect 13725 20584 13737 20587
rect 11112 20556 13737 20584
rect 11112 20544 11118 20556
rect 13725 20553 13737 20556
rect 13771 20553 13783 20587
rect 14093 20587 14151 20593
rect 14093 20584 14105 20587
rect 13725 20547 13783 20553
rect 13832 20556 14105 20584
rect 1302 20476 1308 20528
rect 1360 20516 1366 20528
rect 3605 20519 3663 20525
rect 3605 20516 3617 20519
rect 1360 20488 3617 20516
rect 1360 20476 1366 20488
rect 3605 20485 3617 20488
rect 3651 20485 3663 20519
rect 3605 20479 3663 20485
rect 4724 20488 6684 20516
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 4724 20448 4752 20488
rect 3007 20420 4752 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 4798 20408 4804 20460
rect 4856 20408 4862 20460
rect 5258 20408 5264 20460
rect 5316 20408 5322 20460
rect 6362 20408 6368 20460
rect 6420 20448 6426 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6420 20420 6561 20448
rect 6420 20408 6426 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6656 20448 6684 20488
rect 6822 20476 6828 20528
rect 6880 20516 6886 20528
rect 6880 20488 11468 20516
rect 6880 20476 6886 20488
rect 9217 20451 9275 20457
rect 6656 20420 7604 20448
rect 6549 20411 6607 20417
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 2547 20352 2774 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 2746 20324 2774 20352
rect 5902 20340 5908 20392
rect 5960 20380 5966 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 5960 20352 7021 20380
rect 5960 20340 5966 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7576 20380 7604 20420
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9766 20448 9772 20460
rect 9263 20420 9772 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 9858 20408 9864 20460
rect 9916 20408 9922 20460
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 11440 20448 11468 20488
rect 12526 20476 12532 20528
rect 12584 20476 12590 20528
rect 12621 20519 12679 20525
rect 12621 20485 12633 20519
rect 12667 20516 12679 20519
rect 12802 20516 12808 20528
rect 12667 20488 12808 20516
rect 12667 20485 12679 20488
rect 12621 20479 12679 20485
rect 12802 20476 12808 20488
rect 12860 20476 12866 20528
rect 13446 20476 13452 20528
rect 13504 20516 13510 20528
rect 13832 20516 13860 20556
rect 14093 20553 14105 20556
rect 14139 20553 14151 20587
rect 14093 20547 14151 20553
rect 14918 20544 14924 20596
rect 14976 20544 14982 20596
rect 15562 20544 15568 20596
rect 15620 20544 15626 20596
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15712 20556 15945 20584
rect 15712 20544 15718 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 16022 20544 16028 20596
rect 16080 20544 16086 20596
rect 17126 20544 17132 20596
rect 17184 20544 17190 20596
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 18785 20587 18843 20593
rect 17552 20556 18644 20584
rect 17552 20544 17558 20556
rect 17144 20516 17172 20544
rect 13504 20488 13860 20516
rect 16224 20488 17172 20516
rect 17512 20516 17540 20544
rect 18616 20516 18644 20556
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 18874 20584 18880 20596
rect 18831 20556 18880 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 19484 20556 19717 20584
rect 19484 20544 19490 20556
rect 19705 20553 19717 20556
rect 19751 20584 19763 20587
rect 19886 20584 19892 20596
rect 19751 20556 19892 20584
rect 19751 20553 19763 20556
rect 19705 20547 19763 20553
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 21358 20584 21364 20596
rect 20916 20556 21364 20584
rect 20916 20528 20944 20556
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 25682 20584 25688 20596
rect 22980 20556 25688 20584
rect 22980 20544 22986 20556
rect 19058 20516 19064 20528
rect 17512 20488 17802 20516
rect 18616 20488 19064 20516
rect 13504 20476 13510 20488
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 10551 20420 11376 20448
rect 11440 20420 11713 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 11054 20380 11060 20392
rect 7576 20352 11060 20380
rect 7009 20343 7067 20349
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11149 20383 11207 20389
rect 11149 20349 11161 20383
rect 11195 20349 11207 20383
rect 11348 20380 11376 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11882 20408 11888 20460
rect 11940 20408 11946 20460
rect 12437 20451 12495 20457
rect 12437 20417 12449 20451
rect 12483 20448 12495 20451
rect 12544 20448 12572 20476
rect 12483 20420 12572 20448
rect 14185 20451 14243 20457
rect 12483 20417 12495 20420
rect 12437 20411 12495 20417
rect 14185 20417 14197 20451
rect 14231 20448 14243 20451
rect 14231 20420 15056 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 12526 20380 12532 20392
rect 11348 20352 12532 20380
rect 11149 20343 11207 20349
rect 2746 20284 2780 20324
rect 2774 20272 2780 20284
rect 2832 20272 2838 20324
rect 3326 20272 3332 20324
rect 3384 20312 3390 20324
rect 10778 20312 10784 20324
rect 3384 20284 10784 20312
rect 3384 20272 3390 20284
rect 10778 20272 10784 20284
rect 10836 20272 10842 20324
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 9033 20247 9091 20253
rect 9033 20244 9045 20247
rect 4212 20216 9045 20244
rect 4212 20204 4218 20216
rect 9033 20213 9045 20216
rect 9079 20213 9091 20247
rect 11164 20244 11192 20343
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 14274 20340 14280 20392
rect 14332 20340 14338 20392
rect 15028 20380 15056 20420
rect 15102 20408 15108 20460
rect 15160 20408 15166 20460
rect 15930 20380 15936 20392
rect 15028 20352 15936 20380
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 16224 20389 16252 20488
rect 19058 20476 19064 20488
rect 19116 20476 19122 20528
rect 20898 20516 20904 20528
rect 20746 20488 20904 20516
rect 20898 20476 20904 20488
rect 20956 20476 20962 20528
rect 21177 20519 21235 20525
rect 21177 20485 21189 20519
rect 21223 20516 21235 20519
rect 21542 20516 21548 20528
rect 21223 20488 21548 20516
rect 21223 20485 21235 20488
rect 21177 20479 21235 20485
rect 21542 20476 21548 20488
rect 21600 20476 21606 20528
rect 22373 20519 22431 20525
rect 22373 20485 22385 20519
rect 22419 20516 22431 20519
rect 23750 20516 23756 20528
rect 22419 20488 23756 20516
rect 22419 20485 22431 20488
rect 22373 20479 22431 20485
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 23952 20516 23980 20556
rect 25682 20544 25688 20556
rect 25740 20544 25746 20596
rect 25774 20544 25780 20596
rect 25832 20584 25838 20596
rect 27062 20584 27068 20596
rect 25832 20556 27068 20584
rect 25832 20544 25838 20556
rect 27062 20544 27068 20556
rect 27120 20544 27126 20596
rect 30834 20584 30840 20596
rect 27264 20556 30840 20584
rect 23860 20488 23980 20516
rect 16850 20408 16856 20460
rect 16908 20448 16914 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16908 20420 17049 20448
rect 16908 20408 16914 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 21453 20451 21511 20457
rect 21453 20417 21465 20451
rect 21499 20448 21511 20451
rect 22186 20448 22192 20460
rect 21499 20420 22192 20448
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 23382 20408 23388 20460
rect 23440 20408 23446 20460
rect 23860 20457 23888 20488
rect 24210 20476 24216 20528
rect 24268 20516 24274 20528
rect 26878 20516 26884 20528
rect 24268 20488 24610 20516
rect 25976 20488 26884 20516
rect 24268 20476 24274 20488
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20349 16267 20383
rect 17313 20383 17371 20389
rect 17313 20380 17325 20383
rect 16209 20343 16267 20349
rect 16868 20352 17325 20380
rect 16868 20324 16896 20352
rect 17313 20349 17325 20352
rect 17359 20380 17371 20383
rect 20162 20380 20168 20392
rect 17359 20352 20168 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 20162 20340 20168 20352
rect 20220 20340 20226 20392
rect 21542 20340 21548 20392
rect 21600 20340 21606 20392
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 24121 20383 24179 20389
rect 24121 20349 24133 20383
rect 24167 20380 24179 20383
rect 24670 20380 24676 20392
rect 24167 20352 24676 20380
rect 24167 20349 24179 20352
rect 24121 20343 24179 20349
rect 16850 20272 16856 20324
rect 16908 20272 16914 20324
rect 21560 20312 21588 20340
rect 18984 20284 20208 20312
rect 11790 20244 11796 20256
rect 11164 20216 11796 20244
rect 9033 20207 9091 20213
rect 11790 20204 11796 20216
rect 11848 20204 11854 20256
rect 12802 20204 12808 20256
rect 12860 20244 12866 20256
rect 12989 20247 13047 20253
rect 12989 20244 13001 20247
rect 12860 20216 13001 20244
rect 12860 20204 12866 20216
rect 12989 20213 13001 20216
rect 13035 20244 13047 20247
rect 13170 20244 13176 20256
rect 13035 20216 13176 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 13449 20247 13507 20253
rect 13449 20213 13461 20247
rect 13495 20244 13507 20247
rect 15470 20244 15476 20256
rect 13495 20216 15476 20244
rect 13495 20213 13507 20216
rect 13449 20207 13507 20213
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 16761 20247 16819 20253
rect 16761 20213 16773 20247
rect 16807 20244 16819 20247
rect 17034 20244 17040 20256
rect 16807 20216 17040 20244
rect 16807 20213 16819 20216
rect 16761 20207 16819 20213
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 18984 20244 19012 20284
rect 17184 20216 19012 20244
rect 19337 20247 19395 20253
rect 17184 20204 17190 20216
rect 19337 20213 19349 20247
rect 19383 20244 19395 20247
rect 19610 20244 19616 20256
rect 19383 20216 19616 20244
rect 19383 20213 19395 20216
rect 19337 20207 19395 20213
rect 19610 20204 19616 20216
rect 19668 20204 19674 20256
rect 20180 20244 20208 20284
rect 21376 20284 21588 20312
rect 21376 20256 21404 20284
rect 22278 20272 22284 20324
rect 22336 20312 22342 20324
rect 22572 20312 22600 20343
rect 24670 20340 24676 20352
rect 24728 20380 24734 20392
rect 25976 20380 26004 20488
rect 26878 20476 26884 20488
rect 26936 20476 26942 20528
rect 26050 20408 26056 20460
rect 26108 20408 26114 20460
rect 27264 20457 27292 20556
rect 30834 20544 30840 20556
rect 30892 20584 30898 20596
rect 31478 20584 31484 20596
rect 30892 20556 31484 20584
rect 30892 20544 30898 20556
rect 31478 20544 31484 20556
rect 31536 20584 31542 20596
rect 32490 20584 32496 20596
rect 31536 20556 32496 20584
rect 31536 20544 31542 20556
rect 32490 20544 32496 20556
rect 32548 20584 32554 20596
rect 34054 20584 34060 20596
rect 32548 20556 34060 20584
rect 32548 20544 32554 20556
rect 34054 20544 34060 20556
rect 34112 20544 34118 20596
rect 35253 20587 35311 20593
rect 35253 20553 35265 20587
rect 35299 20584 35311 20587
rect 36170 20584 36176 20596
rect 35299 20556 36176 20584
rect 35299 20553 35311 20556
rect 35253 20547 35311 20553
rect 36170 20544 36176 20556
rect 36228 20544 36234 20596
rect 36446 20544 36452 20596
rect 36504 20544 36510 20596
rect 37458 20544 37464 20596
rect 37516 20584 37522 20596
rect 41141 20587 41199 20593
rect 41141 20584 41153 20587
rect 37516 20556 41153 20584
rect 37516 20544 37522 20556
rect 41141 20553 41153 20556
rect 41187 20553 41199 20587
rect 41141 20547 41199 20553
rect 47854 20544 47860 20596
rect 47912 20584 47918 20596
rect 48041 20587 48099 20593
rect 48041 20584 48053 20587
rect 47912 20556 48053 20584
rect 47912 20544 47918 20556
rect 48041 20553 48053 20556
rect 48087 20553 48099 20587
rect 48041 20547 48099 20553
rect 28902 20516 28908 20528
rect 28750 20488 28908 20516
rect 28902 20476 28908 20488
rect 28960 20476 28966 20528
rect 29178 20476 29184 20528
rect 29236 20516 29242 20528
rect 29825 20519 29883 20525
rect 29825 20516 29837 20519
rect 29236 20488 29837 20516
rect 29236 20476 29242 20488
rect 29825 20485 29837 20488
rect 29871 20485 29883 20519
rect 29825 20479 29883 20485
rect 31018 20476 31024 20528
rect 31076 20476 31082 20528
rect 31113 20519 31171 20525
rect 31113 20485 31125 20519
rect 31159 20516 31171 20519
rect 31294 20516 31300 20528
rect 31159 20488 31300 20516
rect 31159 20485 31171 20488
rect 31113 20479 31171 20485
rect 31294 20476 31300 20488
rect 31352 20476 31358 20528
rect 31757 20519 31815 20525
rect 31757 20485 31769 20519
rect 31803 20516 31815 20519
rect 32122 20516 32128 20528
rect 31803 20488 32128 20516
rect 31803 20485 31815 20488
rect 31757 20479 31815 20485
rect 32122 20476 32128 20488
rect 32180 20476 32186 20528
rect 32398 20476 32404 20528
rect 32456 20516 32462 20528
rect 32456 20488 32614 20516
rect 32456 20476 32462 20488
rect 33686 20476 33692 20528
rect 33744 20516 33750 20528
rect 33781 20519 33839 20525
rect 33781 20516 33793 20519
rect 33744 20488 33793 20516
rect 33744 20476 33750 20488
rect 33781 20485 33793 20488
rect 33827 20516 33839 20519
rect 34422 20516 34428 20528
rect 33827 20488 34428 20516
rect 33827 20485 33839 20488
rect 33781 20479 33839 20485
rect 34422 20476 34428 20488
rect 34480 20476 34486 20528
rect 36464 20516 36492 20544
rect 34808 20488 36492 20516
rect 27249 20451 27307 20457
rect 27249 20417 27261 20451
rect 27295 20417 27307 20451
rect 27249 20411 27307 20417
rect 29733 20451 29791 20457
rect 29733 20417 29745 20451
rect 29779 20448 29791 20451
rect 30190 20448 30196 20460
rect 29779 20420 30196 20448
rect 29779 20417 29791 20420
rect 29733 20411 29791 20417
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 32490 20448 32496 20460
rect 31726 20420 32496 20448
rect 24728 20352 26004 20380
rect 24728 20340 24734 20352
rect 26142 20340 26148 20392
rect 26200 20380 26206 20392
rect 27525 20383 27583 20389
rect 27525 20380 27537 20383
rect 26200 20352 27537 20380
rect 26200 20340 26206 20352
rect 27525 20349 27537 20352
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 28997 20383 29055 20389
rect 28997 20349 29009 20383
rect 29043 20380 29055 20383
rect 29270 20380 29276 20392
rect 29043 20352 29276 20380
rect 29043 20349 29055 20352
rect 28997 20343 29055 20349
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 29546 20340 29552 20392
rect 29604 20340 29610 20392
rect 30558 20380 30564 20392
rect 30024 20352 30564 20380
rect 22336 20284 22600 20312
rect 22336 20272 22342 20284
rect 22738 20272 22744 20324
rect 22796 20312 22802 20324
rect 23201 20315 23259 20321
rect 23201 20312 23213 20315
rect 22796 20284 23213 20312
rect 22796 20272 22802 20284
rect 23201 20281 23213 20284
rect 23247 20281 23259 20315
rect 23201 20275 23259 20281
rect 26050 20272 26056 20324
rect 26108 20312 26114 20324
rect 26605 20315 26663 20321
rect 26605 20312 26617 20315
rect 26108 20284 26617 20312
rect 26108 20272 26114 20284
rect 26605 20281 26617 20284
rect 26651 20281 26663 20315
rect 26605 20275 26663 20281
rect 20622 20244 20628 20256
rect 20180 20216 20628 20244
rect 20622 20204 20628 20216
rect 20680 20204 20686 20256
rect 21358 20204 21364 20256
rect 21416 20204 21422 20256
rect 21542 20204 21548 20256
rect 21600 20244 21606 20256
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 21600 20216 22017 20244
rect 21600 20204 21606 20216
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22005 20207 22063 20213
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 25590 20244 25596 20256
rect 24912 20216 25596 20244
rect 24912 20204 24918 20216
rect 25590 20204 25596 20216
rect 25648 20204 25654 20256
rect 26237 20247 26295 20253
rect 26237 20213 26249 20247
rect 26283 20244 26295 20247
rect 26510 20244 26516 20256
rect 26283 20216 26516 20244
rect 26283 20213 26295 20216
rect 26237 20207 26295 20213
rect 26510 20204 26516 20216
rect 26568 20204 26574 20256
rect 26620 20244 26648 20275
rect 28902 20272 28908 20324
rect 28960 20312 28966 20324
rect 30024 20312 30052 20352
rect 30558 20340 30564 20352
rect 30616 20340 30622 20392
rect 31110 20340 31116 20392
rect 31168 20380 31174 20392
rect 31205 20383 31263 20389
rect 31205 20380 31217 20383
rect 31168 20352 31217 20380
rect 31168 20340 31174 20352
rect 31205 20349 31217 20352
rect 31251 20349 31263 20383
rect 31205 20343 31263 20349
rect 31726 20312 31754 20420
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 34808 20448 34836 20488
rect 36722 20476 36728 20528
rect 36780 20516 36786 20528
rect 37366 20516 37372 20528
rect 36780 20488 37372 20516
rect 36780 20476 36786 20488
rect 37366 20476 37372 20488
rect 37424 20516 37430 20528
rect 37918 20516 37924 20528
rect 37424 20488 37924 20516
rect 37424 20476 37430 20488
rect 37918 20476 37924 20488
rect 37976 20516 37982 20528
rect 37976 20488 38042 20516
rect 37976 20476 37982 20488
rect 39758 20476 39764 20528
rect 39816 20516 39822 20528
rect 40221 20519 40279 20525
rect 40221 20516 40233 20519
rect 39816 20488 40233 20516
rect 39816 20476 39822 20488
rect 40221 20485 40233 20488
rect 40267 20516 40279 20519
rect 41785 20519 41843 20525
rect 41785 20516 41797 20519
rect 40267 20488 41797 20516
rect 40267 20485 40279 20488
rect 40221 20479 40279 20485
rect 41785 20485 41797 20488
rect 41831 20485 41843 20519
rect 41785 20479 41843 20485
rect 34716 20420 34836 20448
rect 32306 20340 32312 20392
rect 32364 20340 32370 20392
rect 34054 20340 34060 20392
rect 34112 20340 34118 20392
rect 34716 20389 34744 20420
rect 34882 20408 34888 20460
rect 34940 20408 34946 20460
rect 35066 20408 35072 20460
rect 35124 20448 35130 20460
rect 35713 20451 35771 20457
rect 35713 20448 35725 20451
rect 35124 20420 35725 20448
rect 35124 20408 35130 20420
rect 35713 20417 35725 20420
rect 35759 20417 35771 20451
rect 35713 20411 35771 20417
rect 36446 20408 36452 20460
rect 36504 20408 36510 20460
rect 36541 20451 36599 20457
rect 36541 20417 36553 20451
rect 36587 20448 36599 20451
rect 37182 20448 37188 20460
rect 36587 20420 37188 20448
rect 36587 20417 36599 20420
rect 36541 20411 36599 20417
rect 37182 20408 37188 20420
rect 37240 20408 37246 20460
rect 39482 20408 39488 20460
rect 39540 20408 39546 20460
rect 39666 20408 39672 20460
rect 39724 20448 39730 20460
rect 40313 20451 40371 20457
rect 40313 20448 40325 20451
rect 39724 20420 40325 20448
rect 39724 20408 39730 20420
rect 40313 20417 40325 20420
rect 40359 20448 40371 20451
rect 48593 20451 48651 20457
rect 40359 20420 41736 20448
rect 40359 20417 40371 20420
rect 40313 20411 40371 20417
rect 34701 20383 34759 20389
rect 34701 20349 34713 20383
rect 34747 20349 34759 20383
rect 34701 20343 34759 20349
rect 34793 20383 34851 20389
rect 34793 20349 34805 20383
rect 34839 20380 34851 20383
rect 34974 20380 34980 20392
rect 34839 20352 34980 20380
rect 34839 20349 34851 20352
rect 34793 20343 34851 20349
rect 34974 20340 34980 20352
rect 35032 20340 35038 20392
rect 36725 20383 36783 20389
rect 35084 20352 36216 20380
rect 28960 20284 30052 20312
rect 30116 20284 31754 20312
rect 28960 20272 28966 20284
rect 30116 20244 30144 20284
rect 31938 20272 31944 20324
rect 31996 20272 32002 20324
rect 26620 20216 30144 20244
rect 30193 20247 30251 20253
rect 30193 20213 30205 20247
rect 30239 20244 30251 20247
rect 30558 20244 30564 20256
rect 30239 20216 30564 20244
rect 30239 20213 30251 20216
rect 30193 20207 30251 20213
rect 30558 20204 30564 20216
rect 30616 20204 30622 20256
rect 30653 20247 30711 20253
rect 30653 20213 30665 20247
rect 30699 20244 30711 20247
rect 30834 20244 30840 20256
rect 30699 20216 30840 20244
rect 30699 20213 30711 20216
rect 30653 20207 30711 20213
rect 30834 20204 30840 20216
rect 30892 20204 30898 20256
rect 31386 20204 31392 20256
rect 31444 20244 31450 20256
rect 35084 20244 35112 20352
rect 35526 20272 35532 20324
rect 35584 20272 35590 20324
rect 35986 20272 35992 20324
rect 36044 20312 36050 20324
rect 36081 20315 36139 20321
rect 36081 20312 36093 20315
rect 36044 20284 36093 20312
rect 36044 20272 36050 20284
rect 36081 20281 36093 20284
rect 36127 20281 36139 20315
rect 36188 20312 36216 20352
rect 36725 20349 36737 20383
rect 36771 20380 36783 20383
rect 37458 20380 37464 20392
rect 36771 20352 37464 20380
rect 36771 20349 36783 20352
rect 36725 20343 36783 20349
rect 37458 20340 37464 20352
rect 37516 20340 37522 20392
rect 37642 20340 37648 20392
rect 37700 20380 37706 20392
rect 39209 20383 39267 20389
rect 39209 20380 39221 20383
rect 37700 20352 39221 20380
rect 37700 20340 37706 20352
rect 39209 20349 39221 20352
rect 39255 20349 39267 20383
rect 39209 20343 39267 20349
rect 40126 20340 40132 20392
rect 40184 20340 40190 20392
rect 41046 20340 41052 20392
rect 41104 20380 41110 20392
rect 41104 20352 41414 20380
rect 41104 20340 41110 20352
rect 36188 20284 37872 20312
rect 36081 20275 36139 20281
rect 31444 20216 35112 20244
rect 37369 20247 37427 20253
rect 31444 20204 31450 20216
rect 37369 20213 37381 20247
rect 37415 20244 37427 20247
rect 37642 20244 37648 20256
rect 37415 20216 37648 20244
rect 37415 20213 37427 20216
rect 37369 20207 37427 20213
rect 37642 20204 37648 20216
rect 37700 20204 37706 20256
rect 37734 20204 37740 20256
rect 37792 20204 37798 20256
rect 37844 20244 37872 20284
rect 39206 20244 39212 20256
rect 37844 20216 39212 20244
rect 39206 20204 39212 20216
rect 39264 20204 39270 20256
rect 40678 20204 40684 20256
rect 40736 20204 40742 20256
rect 41386 20244 41414 20352
rect 41708 20321 41736 20420
rect 48593 20417 48605 20451
rect 48639 20448 48651 20451
rect 48774 20448 48780 20460
rect 48639 20420 48780 20448
rect 48639 20417 48651 20420
rect 48593 20411 48651 20417
rect 48774 20408 48780 20420
rect 48832 20408 48838 20460
rect 49329 20451 49387 20457
rect 49329 20417 49341 20451
rect 49375 20448 49387 20451
rect 49418 20448 49424 20460
rect 49375 20420 49424 20448
rect 49375 20417 49387 20420
rect 49329 20411 49387 20417
rect 47949 20383 48007 20389
rect 47949 20349 47961 20383
rect 47995 20380 48007 20383
rect 49344 20380 49372 20411
rect 49418 20408 49424 20420
rect 49476 20408 49482 20460
rect 47995 20352 49372 20380
rect 47995 20349 48007 20352
rect 47949 20343 48007 20349
rect 41693 20315 41751 20321
rect 41693 20281 41705 20315
rect 41739 20312 41751 20315
rect 49145 20315 49203 20321
rect 49145 20312 49157 20315
rect 41739 20284 49157 20312
rect 41739 20281 41751 20284
rect 41693 20275 41751 20281
rect 49145 20281 49157 20284
rect 49191 20281 49203 20315
rect 49145 20275 49203 20281
rect 48314 20244 48320 20256
rect 41386 20216 48320 20244
rect 48314 20204 48320 20216
rect 48372 20204 48378 20256
rect 48406 20204 48412 20256
rect 48464 20204 48470 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 4798 20000 4804 20052
rect 4856 20040 4862 20052
rect 11333 20043 11391 20049
rect 11333 20040 11345 20043
rect 4856 20012 11345 20040
rect 4856 20000 4862 20012
rect 11333 20009 11345 20012
rect 11379 20009 11391 20043
rect 11333 20003 11391 20009
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12434 20040 12440 20052
rect 12032 20012 12440 20040
rect 12032 20000 12038 20012
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 14458 20000 14464 20052
rect 14516 20000 14522 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 14568 20012 16865 20040
rect 5258 19932 5264 19984
rect 5316 19972 5322 19984
rect 8294 19972 8300 19984
rect 5316 19944 8300 19972
rect 5316 19932 5322 19944
rect 8294 19932 8300 19944
rect 8352 19932 8358 19984
rect 9950 19932 9956 19984
rect 10008 19972 10014 19984
rect 10778 19972 10784 19984
rect 10008 19944 10784 19972
rect 10008 19932 10014 19944
rect 10778 19932 10784 19944
rect 10836 19932 10842 19984
rect 14568 19972 14596 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 18322 20040 18328 20052
rect 18187 20012 18328 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 20346 20040 20352 20052
rect 19168 20012 20352 20040
rect 11900 19944 12112 19972
rect 4246 19864 4252 19916
rect 4304 19864 4310 19916
rect 5718 19864 5724 19916
rect 5776 19904 5782 19916
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5776 19876 6009 19904
rect 5776 19864 5782 19876
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 11900 19904 11928 19944
rect 5997 19867 6055 19873
rect 10152 19876 11928 19904
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 3326 19836 3332 19848
rect 3007 19808 3332 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 5350 19796 5356 19848
rect 5408 19796 5414 19848
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19836 7251 19839
rect 7929 19839 7987 19845
rect 7239 19808 7420 19836
rect 7239 19805 7251 19808
rect 7193 19799 7251 19805
rect 1486 19728 1492 19780
rect 1544 19768 1550 19780
rect 1765 19771 1823 19777
rect 1765 19768 1777 19771
rect 1544 19740 1777 19768
rect 1544 19728 1550 19740
rect 1765 19737 1777 19740
rect 1811 19737 1823 19771
rect 1765 19731 1823 19737
rect 7392 19700 7420 19808
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 9950 19836 9956 19848
rect 7975 19808 9956 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10152 19845 10180 19876
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 12084 19904 12112 19944
rect 13556 19944 14596 19972
rect 13556 19904 13584 19944
rect 14918 19932 14924 19984
rect 14976 19932 14982 19984
rect 15657 19975 15715 19981
rect 15657 19941 15669 19975
rect 15703 19941 15715 19975
rect 18874 19972 18880 19984
rect 15657 19935 15715 19941
rect 17512 19944 18880 19972
rect 15672 19904 15700 19935
rect 12084 19876 13584 19904
rect 13648 19876 15700 19904
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19836 10839 19839
rect 10827 19808 11652 19836
rect 10827 19805 10839 19808
rect 10781 19799 10839 19805
rect 11422 19728 11428 19780
rect 11480 19728 11486 19780
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7392 19672 7757 19700
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 10597 19703 10655 19709
rect 10597 19669 10609 19703
rect 10643 19700 10655 19703
rect 10870 19700 10876 19712
rect 10643 19672 10876 19700
rect 10643 19669 10655 19672
rect 10597 19663 10655 19669
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 11624 19700 11652 19808
rect 11698 19728 11704 19780
rect 11756 19768 11762 19780
rect 12253 19771 12311 19777
rect 12253 19768 12265 19771
rect 11756 19740 12265 19768
rect 11756 19728 11762 19740
rect 12253 19737 12265 19740
rect 12299 19737 12311 19771
rect 12253 19731 12311 19737
rect 12894 19728 12900 19780
rect 12952 19728 12958 19780
rect 13648 19700 13676 19876
rect 16298 19864 16304 19916
rect 16356 19864 16362 19916
rect 17512 19913 17540 19944
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 17586 19864 17592 19916
rect 17644 19904 17650 19916
rect 18785 19907 18843 19913
rect 17644 19876 18736 19904
rect 17644 19864 17650 19876
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19836 15163 19839
rect 15470 19836 15476 19848
rect 15151 19808 15476 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 16114 19836 16120 19848
rect 15672 19808 16120 19836
rect 11624 19672 13676 19700
rect 13725 19703 13783 19709
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 15672 19700 15700 19808
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19836 18567 19839
rect 18598 19836 18604 19848
rect 18555 19808 18604 19836
rect 18555 19805 18567 19808
rect 18509 19799 18567 19805
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 18708 19836 18736 19876
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 19168 19904 19196 20012
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 22370 20040 22376 20052
rect 20456 20012 22376 20040
rect 19242 19932 19248 19984
rect 19300 19972 19306 19984
rect 19613 19975 19671 19981
rect 19613 19972 19625 19975
rect 19300 19944 19625 19972
rect 19300 19932 19306 19944
rect 19613 19941 19625 19944
rect 19659 19941 19671 19975
rect 20456 19972 20484 20012
rect 22370 20000 22376 20012
rect 22428 20000 22434 20052
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 25593 20043 25651 20049
rect 25593 20040 25605 20043
rect 22520 20012 25605 20040
rect 22520 20000 22526 20012
rect 25593 20009 25605 20012
rect 25639 20009 25651 20043
rect 25593 20003 25651 20009
rect 26068 20012 26740 20040
rect 24029 19975 24087 19981
rect 19613 19935 19671 19941
rect 19720 19944 20484 19972
rect 22204 19944 23980 19972
rect 18831 19876 19196 19904
rect 19337 19907 19395 19913
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19337 19873 19349 19907
rect 19383 19904 19395 19907
rect 19720 19904 19748 19944
rect 20990 19904 20996 19916
rect 19383 19876 19748 19904
rect 20180 19876 20996 19904
rect 19383 19873 19395 19876
rect 19337 19867 19395 19873
rect 19352 19836 19380 19867
rect 20180 19836 20208 19876
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 21634 19904 21640 19916
rect 21508 19876 21640 19904
rect 21508 19864 21514 19876
rect 21634 19864 21640 19876
rect 21692 19904 21698 19916
rect 22204 19904 22232 19944
rect 21692 19876 22232 19904
rect 22281 19907 22339 19913
rect 21692 19864 21698 19876
rect 22281 19873 22293 19907
rect 22327 19904 22339 19907
rect 22830 19904 22836 19916
rect 22327 19876 22836 19904
rect 22327 19873 22339 19876
rect 22281 19867 22339 19873
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 23385 19907 23443 19913
rect 23385 19904 23397 19907
rect 22940 19876 23397 19904
rect 18708 19808 19380 19836
rect 19720 19808 20208 19836
rect 20257 19839 20315 19845
rect 16025 19771 16083 19777
rect 16025 19737 16037 19771
rect 16071 19768 16083 19771
rect 18322 19768 18328 19780
rect 16071 19740 18328 19768
rect 16071 19737 16083 19740
rect 16025 19731 16083 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 19720 19768 19748 19808
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 20346 19836 20352 19848
rect 20303 19808 20352 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 20898 19796 20904 19848
rect 20956 19796 20962 19848
rect 22741 19839 22799 19845
rect 22741 19805 22753 19839
rect 22787 19836 22799 19839
rect 22940 19836 22968 19876
rect 23385 19873 23397 19876
rect 23431 19873 23443 19907
rect 23385 19867 23443 19873
rect 22787 19808 22968 19836
rect 22787 19805 22799 19808
rect 22741 19799 22799 19805
rect 23014 19796 23020 19848
rect 23072 19796 23078 19848
rect 18616 19740 19748 19768
rect 19797 19771 19855 19777
rect 13771 19672 15700 19700
rect 16117 19703 16175 19709
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 16117 19669 16129 19703
rect 16163 19700 16175 19703
rect 17126 19700 17132 19712
rect 16163 19672 17132 19700
rect 16163 19669 16175 19672
rect 16117 19663 16175 19669
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 17218 19660 17224 19712
rect 17276 19660 17282 19712
rect 17310 19660 17316 19712
rect 17368 19660 17374 19712
rect 18616 19709 18644 19740
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 20714 19768 20720 19780
rect 19843 19740 20720 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 22005 19771 22063 19777
rect 22005 19737 22017 19771
rect 22051 19768 22063 19771
rect 22094 19768 22100 19780
rect 22051 19740 22100 19768
rect 22051 19737 22063 19740
rect 22005 19731 22063 19737
rect 22094 19728 22100 19740
rect 22152 19728 22158 19780
rect 22370 19728 22376 19780
rect 22428 19768 22434 19780
rect 23400 19768 23428 19867
rect 23474 19864 23480 19916
rect 23532 19864 23538 19916
rect 23569 19907 23627 19913
rect 23569 19873 23581 19907
rect 23615 19904 23627 19907
rect 23842 19904 23848 19916
rect 23615 19876 23848 19904
rect 23615 19873 23627 19876
rect 23569 19867 23627 19873
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 23952 19904 23980 19944
rect 24029 19941 24041 19975
rect 24075 19972 24087 19975
rect 25774 19972 25780 19984
rect 24075 19944 25780 19972
rect 24075 19941 24087 19944
rect 24029 19935 24087 19941
rect 25774 19932 25780 19944
rect 25832 19932 25838 19984
rect 24302 19904 24308 19916
rect 23952 19876 24308 19904
rect 24302 19864 24308 19876
rect 24360 19864 24366 19916
rect 24578 19864 24584 19916
rect 24636 19864 24642 19916
rect 26068 19904 26096 20012
rect 24964 19876 26096 19904
rect 26237 19907 26295 19913
rect 23492 19836 23520 19864
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23492 19808 23673 19836
rect 23661 19805 23673 19808
rect 23707 19805 23719 19839
rect 23661 19799 23719 19805
rect 24964 19768 24992 19876
rect 26237 19873 26249 19907
rect 26283 19873 26295 19907
rect 26237 19867 26295 19873
rect 25222 19796 25228 19848
rect 25280 19836 25286 19848
rect 26252 19836 26280 19867
rect 25280 19808 26280 19836
rect 26712 19836 26740 20012
rect 26786 20000 26792 20052
rect 26844 20000 26850 20052
rect 27062 20000 27068 20052
rect 27120 20040 27126 20052
rect 28997 20043 29055 20049
rect 28997 20040 29009 20043
rect 27120 20012 29009 20040
rect 27120 20000 27126 20012
rect 28997 20009 29009 20012
rect 29043 20040 29055 20043
rect 30374 20040 30380 20052
rect 29043 20012 30380 20040
rect 29043 20009 29055 20012
rect 28997 20003 29055 20009
rect 30374 20000 30380 20012
rect 30432 20000 30438 20052
rect 31665 20043 31723 20049
rect 31665 20009 31677 20043
rect 31711 20040 31723 20043
rect 32766 20040 32772 20052
rect 31711 20012 32772 20040
rect 31711 20009 31723 20012
rect 31665 20003 31723 20009
rect 32766 20000 32772 20012
rect 32824 20000 32830 20052
rect 34330 20040 34336 20052
rect 33612 20012 34336 20040
rect 28902 19972 28908 19984
rect 27724 19944 28908 19972
rect 26878 19864 26884 19916
rect 26936 19904 26942 19916
rect 27341 19907 27399 19913
rect 27341 19904 27353 19907
rect 26936 19876 27353 19904
rect 26936 19864 26942 19876
rect 27341 19873 27353 19876
rect 27387 19873 27399 19907
rect 27341 19867 27399 19873
rect 27724 19836 27752 19944
rect 28902 19932 28908 19944
rect 28960 19972 28966 19984
rect 29273 19975 29331 19981
rect 29273 19972 29285 19975
rect 28960 19944 29285 19972
rect 28960 19932 28966 19944
rect 29273 19941 29285 19944
rect 29319 19941 29331 19975
rect 29273 19935 29331 19941
rect 30300 19944 32720 19972
rect 30300 19916 30328 19944
rect 28350 19864 28356 19916
rect 28408 19904 28414 19916
rect 28537 19907 28595 19913
rect 28537 19904 28549 19907
rect 28408 19876 28549 19904
rect 28408 19864 28414 19876
rect 28537 19873 28549 19876
rect 28583 19873 28595 19907
rect 28537 19867 28595 19873
rect 30006 19864 30012 19916
rect 30064 19904 30070 19916
rect 30190 19904 30196 19916
rect 30064 19876 30196 19904
rect 30064 19864 30070 19876
rect 30190 19864 30196 19876
rect 30248 19864 30254 19916
rect 30282 19864 30288 19916
rect 30340 19864 30346 19916
rect 32692 19913 32720 19944
rect 33612 19913 33640 20012
rect 34330 20000 34336 20012
rect 34388 20000 34394 20052
rect 34882 20000 34888 20052
rect 34940 20040 34946 20052
rect 36906 20040 36912 20052
rect 34940 20012 36912 20040
rect 34940 20000 34946 20012
rect 36906 20000 36912 20012
rect 36964 20000 36970 20052
rect 37826 20000 37832 20052
rect 37884 20040 37890 20052
rect 39025 20043 39083 20049
rect 39025 20040 39037 20043
rect 37884 20012 39037 20040
rect 37884 20000 37890 20012
rect 39025 20009 39037 20012
rect 39071 20040 39083 20043
rect 39942 20040 39948 20052
rect 39071 20012 39948 20040
rect 39071 20009 39083 20012
rect 39025 20003 39083 20009
rect 39942 20000 39948 20012
rect 40000 20000 40006 20052
rect 40494 20000 40500 20052
rect 40552 20040 40558 20052
rect 41233 20043 41291 20049
rect 41233 20040 41245 20043
rect 40552 20012 41245 20040
rect 40552 20000 40558 20012
rect 41233 20009 41245 20012
rect 41279 20009 41291 20043
rect 41233 20003 41291 20009
rect 48774 20000 48780 20052
rect 48832 20000 48838 20052
rect 34149 19975 34207 19981
rect 34149 19941 34161 19975
rect 34195 19972 34207 19975
rect 34698 19972 34704 19984
rect 34195 19944 34704 19972
rect 34195 19941 34207 19944
rect 34149 19935 34207 19941
rect 34698 19932 34704 19944
rect 34756 19932 34762 19984
rect 43438 19972 43444 19984
rect 34900 19944 43444 19972
rect 31113 19907 31171 19913
rect 31113 19873 31125 19907
rect 31159 19904 31171 19907
rect 32677 19907 32735 19913
rect 31159 19876 32444 19904
rect 31159 19873 31171 19876
rect 31113 19867 31171 19873
rect 28626 19836 28632 19848
rect 26712 19808 27752 19836
rect 27816 19808 28632 19836
rect 25280 19796 25286 19808
rect 27816 19780 27844 19808
rect 28626 19796 28632 19808
rect 28684 19796 28690 19848
rect 30098 19836 30104 19848
rect 29012 19808 30104 19836
rect 22428 19740 22876 19768
rect 23400 19740 24992 19768
rect 25133 19771 25191 19777
rect 22428 19728 22434 19740
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19669 18659 19703
rect 18601 19663 18659 19669
rect 19058 19660 19064 19712
rect 19116 19700 19122 19712
rect 19978 19700 19984 19712
rect 19116 19672 19984 19700
rect 19116 19660 19122 19672
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 20254 19660 20260 19712
rect 20312 19700 20318 19712
rect 20533 19703 20591 19709
rect 20533 19700 20545 19703
rect 20312 19672 20545 19700
rect 20312 19660 20318 19672
rect 20533 19669 20545 19672
rect 20579 19669 20591 19703
rect 20533 19663 20591 19669
rect 22646 19660 22652 19712
rect 22704 19660 22710 19712
rect 22848 19700 22876 19740
rect 25133 19737 25145 19771
rect 25179 19768 25191 19771
rect 25961 19771 26019 19777
rect 25179 19740 25912 19768
rect 25179 19737 25191 19740
rect 25133 19731 25191 19737
rect 25038 19700 25044 19712
rect 22848 19672 25044 19700
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 25314 19660 25320 19712
rect 25372 19660 25378 19712
rect 25884 19700 25912 19740
rect 25961 19737 25973 19771
rect 26007 19768 26019 19771
rect 27798 19768 27804 19780
rect 26007 19740 27804 19768
rect 26007 19737 26019 19740
rect 25961 19731 26019 19737
rect 27798 19728 27804 19740
rect 27856 19728 27862 19780
rect 28445 19771 28503 19777
rect 28445 19737 28457 19771
rect 28491 19768 28503 19771
rect 29012 19768 29040 19808
rect 30098 19796 30104 19808
rect 30156 19796 30162 19848
rect 31570 19836 31576 19848
rect 30576 19808 31576 19836
rect 30576 19768 30604 19808
rect 31570 19796 31576 19808
rect 31628 19796 31634 19848
rect 28491 19740 29040 19768
rect 29104 19740 30604 19768
rect 31205 19771 31263 19777
rect 28491 19737 28503 19740
rect 28445 19731 28503 19737
rect 26053 19703 26111 19709
rect 26053 19700 26065 19703
rect 25884 19672 26065 19700
rect 26053 19669 26065 19672
rect 26099 19700 26111 19703
rect 26694 19700 26700 19712
rect 26099 19672 26700 19700
rect 26099 19669 26111 19672
rect 26053 19663 26111 19669
rect 26694 19660 26700 19672
rect 26752 19660 26758 19712
rect 27062 19660 27068 19712
rect 27120 19700 27126 19712
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 27120 19672 27169 19700
rect 27120 19660 27126 19672
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 27157 19663 27215 19669
rect 27246 19660 27252 19712
rect 27304 19660 27310 19712
rect 27614 19660 27620 19712
rect 27672 19700 27678 19712
rect 27985 19703 28043 19709
rect 27985 19700 27997 19703
rect 27672 19672 27997 19700
rect 27672 19660 27678 19672
rect 27985 19669 27997 19672
rect 28031 19669 28043 19703
rect 27985 19663 28043 19669
rect 28353 19703 28411 19709
rect 28353 19669 28365 19703
rect 28399 19700 28411 19703
rect 29104 19700 29132 19740
rect 31205 19737 31217 19771
rect 31251 19768 31263 19771
rect 31938 19768 31944 19780
rect 31251 19740 31944 19768
rect 31251 19737 31263 19740
rect 31205 19731 31263 19737
rect 31938 19728 31944 19740
rect 31996 19728 32002 19780
rect 28399 19672 29132 19700
rect 28399 19669 28411 19672
rect 28353 19663 28411 19669
rect 29178 19660 29184 19712
rect 29236 19700 29242 19712
rect 29546 19700 29552 19712
rect 29236 19672 29552 19700
rect 29236 19660 29242 19672
rect 29546 19660 29552 19672
rect 29604 19660 29610 19712
rect 29730 19660 29736 19712
rect 29788 19660 29794 19712
rect 30098 19660 30104 19712
rect 30156 19660 30162 19712
rect 31294 19660 31300 19712
rect 31352 19660 31358 19712
rect 32122 19660 32128 19712
rect 32180 19660 32186 19712
rect 32416 19700 32444 19876
rect 32677 19873 32689 19907
rect 32723 19873 32735 19907
rect 32677 19867 32735 19873
rect 33597 19907 33655 19913
rect 33597 19873 33609 19907
rect 33643 19873 33655 19907
rect 33597 19867 33655 19873
rect 33689 19907 33747 19913
rect 33689 19873 33701 19907
rect 33735 19904 33747 19907
rect 34900 19904 34928 19944
rect 43438 19932 43444 19944
rect 43496 19932 43502 19984
rect 33735 19876 34928 19904
rect 33735 19873 33747 19876
rect 33689 19867 33747 19873
rect 32493 19839 32551 19845
rect 32493 19805 32505 19839
rect 32539 19836 32551 19839
rect 33778 19836 33784 19848
rect 32539 19808 33784 19836
rect 32539 19805 32551 19808
rect 32493 19799 32551 19805
rect 33778 19796 33784 19808
rect 33836 19796 33842 19848
rect 32585 19771 32643 19777
rect 32585 19737 32597 19771
rect 32631 19768 32643 19771
rect 33888 19768 33916 19876
rect 35066 19864 35072 19916
rect 35124 19864 35130 19916
rect 36722 19864 36728 19916
rect 36780 19864 36786 19916
rect 38013 19907 38071 19913
rect 38013 19873 38025 19907
rect 38059 19904 38071 19907
rect 38378 19904 38384 19916
rect 38059 19876 38384 19904
rect 38059 19873 38071 19876
rect 38013 19867 38071 19873
rect 38378 19864 38384 19876
rect 38436 19864 38442 19916
rect 39390 19864 39396 19916
rect 39448 19904 39454 19916
rect 40129 19907 40187 19913
rect 40129 19904 40141 19907
rect 39448 19876 40141 19904
rect 39448 19864 39454 19876
rect 40129 19873 40141 19876
rect 40175 19873 40187 19907
rect 40129 19867 40187 19873
rect 40313 19907 40371 19913
rect 40313 19873 40325 19907
rect 40359 19904 40371 19907
rect 40494 19904 40500 19916
rect 40359 19876 40500 19904
rect 40359 19873 40371 19876
rect 40313 19867 40371 19873
rect 40494 19864 40500 19876
rect 40552 19864 40558 19916
rect 35158 19796 35164 19848
rect 35216 19836 35222 19848
rect 35253 19839 35311 19845
rect 35253 19836 35265 19839
rect 35216 19808 35265 19836
rect 35216 19796 35222 19808
rect 35253 19805 35265 19808
rect 35299 19805 35311 19839
rect 35253 19799 35311 19805
rect 37826 19796 37832 19848
rect 37884 19836 37890 19848
rect 38105 19839 38163 19845
rect 38105 19836 38117 19839
rect 37884 19808 38117 19836
rect 37884 19796 37890 19808
rect 38105 19805 38117 19808
rect 38151 19805 38163 19839
rect 38105 19799 38163 19805
rect 38194 19796 38200 19848
rect 38252 19836 38258 19848
rect 38841 19839 38899 19845
rect 38841 19836 38853 19839
rect 38252 19808 38853 19836
rect 38252 19796 38258 19808
rect 38841 19805 38853 19808
rect 38887 19836 38899 19839
rect 40218 19836 40224 19848
rect 38887 19808 40224 19836
rect 38887 19805 38899 19808
rect 38841 19799 38899 19805
rect 40218 19796 40224 19808
rect 40276 19796 40282 19848
rect 40402 19796 40408 19848
rect 40460 19836 40466 19848
rect 41049 19839 41107 19845
rect 41049 19836 41061 19839
rect 40460 19808 41061 19836
rect 40460 19796 40466 19808
rect 41049 19805 41061 19808
rect 41095 19836 41107 19839
rect 42702 19836 42708 19848
rect 41095 19808 42708 19836
rect 41095 19805 41107 19808
rect 41049 19799 41107 19805
rect 42702 19796 42708 19808
rect 42760 19796 42766 19848
rect 32631 19740 33916 19768
rect 32631 19737 32643 19740
rect 32585 19731 32643 19737
rect 34238 19728 34244 19780
rect 34296 19768 34302 19780
rect 36262 19768 36268 19780
rect 34296 19740 36268 19768
rect 34296 19728 34302 19740
rect 36262 19728 36268 19740
rect 36320 19728 36326 19780
rect 36449 19771 36507 19777
rect 36449 19737 36461 19771
rect 36495 19768 36507 19771
rect 40034 19768 40040 19780
rect 36495 19740 40040 19768
rect 36495 19737 36507 19740
rect 36449 19731 36507 19737
rect 40034 19728 40040 19740
rect 40092 19728 40098 19780
rect 48593 19771 48651 19777
rect 48593 19737 48605 19771
rect 48639 19768 48651 19771
rect 49237 19771 49295 19777
rect 49237 19768 49249 19771
rect 48639 19740 49249 19768
rect 48639 19737 48651 19740
rect 48593 19731 48651 19737
rect 49237 19737 49249 19740
rect 49283 19768 49295 19771
rect 49326 19768 49332 19780
rect 49283 19740 49332 19768
rect 49283 19737 49295 19740
rect 49237 19731 49295 19737
rect 49326 19728 49332 19740
rect 49384 19728 49390 19780
rect 33594 19700 33600 19712
rect 32416 19672 33600 19700
rect 33594 19660 33600 19672
rect 33652 19660 33658 19712
rect 34330 19660 34336 19712
rect 34388 19700 34394 19712
rect 34425 19703 34483 19709
rect 34425 19700 34437 19703
rect 34388 19672 34437 19700
rect 34388 19660 34394 19672
rect 34425 19669 34437 19672
rect 34471 19669 34483 19703
rect 34425 19663 34483 19669
rect 35161 19703 35219 19709
rect 35161 19669 35173 19703
rect 35207 19700 35219 19703
rect 35342 19700 35348 19712
rect 35207 19672 35348 19700
rect 35207 19669 35219 19672
rect 35161 19663 35219 19669
rect 35342 19660 35348 19672
rect 35400 19660 35406 19712
rect 35621 19703 35679 19709
rect 35621 19669 35633 19703
rect 35667 19700 35679 19703
rect 35802 19700 35808 19712
rect 35667 19672 35808 19700
rect 35667 19669 35679 19672
rect 35621 19663 35679 19669
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 35894 19660 35900 19712
rect 35952 19700 35958 19712
rect 36081 19703 36139 19709
rect 36081 19700 36093 19703
rect 35952 19672 36093 19700
rect 35952 19660 35958 19672
rect 36081 19669 36093 19672
rect 36127 19669 36139 19703
rect 36081 19663 36139 19669
rect 36538 19660 36544 19712
rect 36596 19660 36602 19712
rect 37369 19703 37427 19709
rect 37369 19669 37381 19703
rect 37415 19700 37427 19703
rect 37550 19700 37556 19712
rect 37415 19672 37556 19700
rect 37415 19669 37427 19672
rect 37369 19663 37427 19669
rect 37550 19660 37556 19672
rect 37608 19660 37614 19712
rect 38470 19660 38476 19712
rect 38528 19700 38534 19712
rect 38565 19703 38623 19709
rect 38565 19700 38577 19703
rect 38528 19672 38577 19700
rect 38528 19660 38534 19672
rect 38565 19669 38577 19672
rect 38611 19669 38623 19703
rect 38565 19663 38623 19669
rect 39574 19660 39580 19712
rect 39632 19660 39638 19712
rect 40773 19703 40831 19709
rect 40773 19669 40785 19703
rect 40819 19700 40831 19703
rect 40862 19700 40868 19712
rect 40819 19672 40868 19700
rect 40819 19669 40831 19672
rect 40773 19663 40831 19669
rect 40862 19660 40868 19672
rect 40920 19660 40926 19712
rect 49142 19660 49148 19712
rect 49200 19660 49206 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 7282 19456 7288 19508
rect 7340 19496 7346 19508
rect 7742 19496 7748 19508
rect 7340 19468 7748 19496
rect 7340 19456 7346 19468
rect 7742 19456 7748 19468
rect 7800 19496 7806 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 7800 19468 10977 19496
rect 7800 19456 7806 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 13504 19468 14504 19496
rect 13504 19456 13510 19468
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 3476 19400 3617 19428
rect 3476 19388 3482 19400
rect 3605 19397 3617 19400
rect 3651 19397 3663 19431
rect 9214 19428 9220 19440
rect 3605 19391 3663 19397
rect 4540 19400 9220 19428
rect 1762 19320 1768 19372
rect 1820 19320 1826 19372
rect 2961 19363 3019 19369
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 4540 19360 4568 19400
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 10505 19431 10563 19437
rect 10505 19397 10517 19431
rect 10551 19428 10563 19431
rect 12802 19428 12808 19440
rect 10551 19400 12808 19428
rect 10551 19397 10563 19400
rect 10505 19391 10563 19397
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 14476 19428 14504 19468
rect 15010 19456 15016 19508
rect 15068 19496 15074 19508
rect 15381 19499 15439 19505
rect 15381 19496 15393 19499
rect 15068 19468 15393 19496
rect 15068 19456 15074 19468
rect 15381 19465 15393 19468
rect 15427 19465 15439 19499
rect 15381 19459 15439 19465
rect 15930 19456 15936 19508
rect 15988 19496 15994 19508
rect 16853 19499 16911 19505
rect 16853 19496 16865 19499
rect 15988 19468 16865 19496
rect 15988 19456 15994 19468
rect 16853 19465 16865 19468
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 17310 19456 17316 19508
rect 17368 19496 17374 19508
rect 19886 19496 19892 19508
rect 17368 19468 19892 19496
rect 17368 19456 17374 19468
rect 19886 19456 19892 19468
rect 19944 19456 19950 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 23934 19496 23940 19508
rect 21223 19468 23940 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 24302 19456 24308 19508
rect 24360 19496 24366 19508
rect 25222 19496 25228 19508
rect 24360 19468 25228 19496
rect 24360 19456 24366 19468
rect 25222 19456 25228 19468
rect 25280 19456 25286 19508
rect 26050 19456 26056 19508
rect 26108 19496 26114 19508
rect 26145 19499 26203 19505
rect 26145 19496 26157 19499
rect 26108 19468 26157 19496
rect 26108 19456 26114 19468
rect 26145 19465 26157 19468
rect 26191 19465 26203 19499
rect 28350 19496 28356 19508
rect 26145 19459 26203 19465
rect 26620 19468 28356 19496
rect 16022 19428 16028 19440
rect 3007 19332 4568 19360
rect 4801 19363 4859 19369
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 5445 19363 5503 19369
rect 4847 19332 5396 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 5261 19295 5319 19301
rect 5261 19292 5273 19295
rect 3936 19264 5273 19292
rect 3936 19252 3942 19264
rect 5261 19261 5273 19264
rect 5307 19261 5319 19295
rect 5368 19292 5396 19332
rect 5445 19329 5457 19363
rect 5491 19360 5503 19363
rect 5810 19360 5816 19372
rect 5491 19332 5816 19360
rect 5491 19329 5503 19332
rect 5445 19323 5503 19329
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 11149 19363 11207 19369
rect 9640 19332 11100 19360
rect 9640 19320 9646 19332
rect 6822 19292 6828 19304
rect 5368 19264 6828 19292
rect 5261 19255 5319 19261
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 9858 19252 9864 19304
rect 9916 19252 9922 19304
rect 11072 19292 11100 19332
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 11606 19360 11612 19372
rect 11195 19332 11612 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 12158 19360 12164 19372
rect 11747 19332 12164 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12894 19360 12900 19372
rect 12492 19332 12900 19360
rect 12492 19320 12498 19332
rect 12894 19320 12900 19332
rect 12952 19360 12958 19372
rect 13004 19360 13032 19414
rect 14476 19400 16028 19428
rect 14476 19369 14504 19400
rect 16022 19388 16028 19400
rect 16080 19428 16086 19440
rect 16942 19428 16948 19440
rect 16080 19400 16948 19428
rect 16080 19388 16086 19400
rect 16942 19388 16948 19400
rect 17000 19388 17006 19440
rect 17494 19388 17500 19440
rect 17552 19428 17558 19440
rect 17552 19400 18630 19428
rect 17552 19388 17558 19400
rect 19702 19388 19708 19440
rect 19760 19428 19766 19440
rect 20346 19428 20352 19440
rect 19760 19400 20352 19428
rect 19760 19388 19766 19400
rect 20346 19388 20352 19400
rect 20404 19428 20410 19440
rect 23474 19428 23480 19440
rect 20404 19400 23480 19428
rect 20404 19388 20410 19400
rect 23474 19388 23480 19400
rect 23532 19388 23538 19440
rect 24210 19388 24216 19440
rect 24268 19388 24274 19440
rect 26237 19431 26295 19437
rect 26237 19397 26249 19431
rect 26283 19428 26295 19431
rect 26510 19428 26516 19440
rect 26283 19400 26516 19428
rect 26283 19397 26295 19400
rect 26237 19391 26295 19397
rect 26510 19388 26516 19400
rect 26568 19388 26574 19440
rect 12952 19332 13032 19360
rect 14461 19363 14519 19369
rect 12952 19320 12958 19332
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 15194 19360 15200 19372
rect 14461 19323 14519 19329
rect 15120 19332 15200 19360
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11072 19264 11989 19292
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 11977 19255 12035 19261
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 15013 19295 15071 19301
rect 14231 19264 14964 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 12250 19184 12256 19236
rect 12308 19224 12314 19236
rect 14936 19224 14964 19264
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15120 19292 15148 19332
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15059 19264 15148 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15286 19252 15292 19304
rect 15344 19292 15350 19304
rect 15488 19292 15516 19323
rect 16206 19320 16212 19372
rect 16264 19320 16270 19372
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 17092 19332 17233 19360
rect 17092 19320 17098 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17586 19360 17592 19372
rect 17359 19332 17592 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19360 18107 19363
rect 21085 19363 21143 19369
rect 18095 19332 18644 19360
rect 18095 19329 18107 19332
rect 18049 19323 18107 19329
rect 18616 19304 18644 19332
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 22554 19360 22560 19372
rect 21131 19332 22560 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 22554 19320 22560 19332
rect 22612 19320 22618 19372
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 22925 19363 22983 19369
rect 22925 19360 22937 19363
rect 22704 19332 22937 19360
rect 22704 19320 22710 19332
rect 22925 19329 22937 19332
rect 22971 19360 22983 19363
rect 23290 19360 23296 19372
rect 22971 19332 23296 19360
rect 22971 19329 22983 19332
rect 22925 19323 22983 19329
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19360 25283 19363
rect 25682 19360 25688 19372
rect 25271 19332 25688 19360
rect 25271 19329 25283 19332
rect 25225 19323 25283 19329
rect 25682 19320 25688 19332
rect 25740 19320 25746 19372
rect 26620 19360 26648 19468
rect 28350 19456 28356 19468
rect 28408 19456 28414 19508
rect 28445 19499 28503 19505
rect 28445 19465 28457 19499
rect 28491 19496 28503 19499
rect 28718 19496 28724 19508
rect 28491 19468 28724 19496
rect 28491 19465 28503 19468
rect 28445 19459 28503 19465
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 28810 19456 28816 19508
rect 28868 19496 28874 19508
rect 31386 19496 31392 19508
rect 28868 19468 31392 19496
rect 28868 19456 28874 19468
rect 31386 19456 31392 19468
rect 31444 19456 31450 19508
rect 31662 19456 31668 19508
rect 31720 19496 31726 19508
rect 32677 19499 32735 19505
rect 32677 19496 32689 19499
rect 31720 19468 32689 19496
rect 31720 19456 31726 19468
rect 32677 19465 32689 19468
rect 32723 19465 32735 19499
rect 32677 19459 32735 19465
rect 32858 19456 32864 19508
rect 32916 19496 32922 19508
rect 33045 19499 33103 19505
rect 33045 19496 33057 19499
rect 32916 19468 33057 19496
rect 32916 19456 32922 19468
rect 33045 19465 33057 19468
rect 33091 19465 33103 19499
rect 33045 19459 33103 19465
rect 33781 19499 33839 19505
rect 33781 19465 33793 19499
rect 33827 19496 33839 19499
rect 34514 19496 34520 19508
rect 33827 19468 34520 19496
rect 33827 19465 33839 19468
rect 33781 19459 33839 19465
rect 26694 19388 26700 19440
rect 26752 19428 26758 19440
rect 29638 19428 29644 19440
rect 26752 19400 29644 19428
rect 26752 19388 26758 19400
rect 29638 19388 29644 19400
rect 29696 19388 29702 19440
rect 31478 19388 31484 19440
rect 31536 19388 31542 19440
rect 32490 19388 32496 19440
rect 32548 19428 32554 19440
rect 33796 19428 33824 19459
rect 34514 19456 34520 19468
rect 34572 19456 34578 19508
rect 34882 19456 34888 19508
rect 34940 19496 34946 19508
rect 35069 19499 35127 19505
rect 35069 19496 35081 19499
rect 34940 19468 35081 19496
rect 34940 19456 34946 19468
rect 35069 19465 35081 19468
rect 35115 19465 35127 19499
rect 35069 19459 35127 19465
rect 35437 19499 35495 19505
rect 35437 19465 35449 19499
rect 35483 19496 35495 19499
rect 36538 19496 36544 19508
rect 35483 19468 36544 19496
rect 35483 19465 35495 19468
rect 35437 19459 35495 19465
rect 36538 19456 36544 19468
rect 36596 19456 36602 19508
rect 36906 19456 36912 19508
rect 36964 19496 36970 19508
rect 37277 19499 37335 19505
rect 37277 19496 37289 19499
rect 36964 19468 37289 19496
rect 36964 19456 36970 19468
rect 37277 19465 37289 19468
rect 37323 19465 37335 19499
rect 37277 19459 37335 19465
rect 37366 19456 37372 19508
rect 37424 19496 37430 19508
rect 37461 19499 37519 19505
rect 37461 19496 37473 19499
rect 37424 19468 37473 19496
rect 37424 19456 37430 19468
rect 37461 19465 37473 19468
rect 37507 19496 37519 19499
rect 37918 19496 37924 19508
rect 37507 19468 37924 19496
rect 37507 19465 37519 19468
rect 37461 19459 37519 19465
rect 37918 19456 37924 19468
rect 37976 19496 37982 19508
rect 39574 19496 39580 19508
rect 37976 19468 39580 19496
rect 37976 19456 37982 19468
rect 32548 19400 33824 19428
rect 32548 19388 32554 19400
rect 33962 19388 33968 19440
rect 34020 19428 34026 19440
rect 36173 19431 36231 19437
rect 36173 19428 36185 19431
rect 34020 19400 36185 19428
rect 34020 19388 34026 19400
rect 36173 19397 36185 19400
rect 36219 19397 36231 19431
rect 38120 19428 38148 19468
rect 39574 19456 39580 19468
rect 39632 19456 39638 19508
rect 40034 19456 40040 19508
rect 40092 19496 40098 19508
rect 40129 19499 40187 19505
rect 40129 19496 40141 19499
rect 40092 19468 40141 19496
rect 40092 19456 40098 19468
rect 40129 19465 40141 19468
rect 40175 19465 40187 19499
rect 40129 19459 40187 19465
rect 40589 19499 40647 19505
rect 40589 19465 40601 19499
rect 40635 19496 40647 19499
rect 41046 19496 41052 19508
rect 40635 19468 41052 19496
rect 40635 19465 40647 19468
rect 40589 19459 40647 19465
rect 41046 19456 41052 19468
rect 41104 19496 41110 19508
rect 41325 19499 41383 19505
rect 41325 19496 41337 19499
rect 41104 19468 41337 19496
rect 41104 19456 41110 19468
rect 41325 19465 41337 19468
rect 41371 19465 41383 19499
rect 41325 19459 41383 19465
rect 38120 19400 38226 19428
rect 36173 19391 36231 19397
rect 39482 19388 39488 19440
rect 39540 19428 39546 19440
rect 40497 19431 40555 19437
rect 39540 19400 39712 19428
rect 39540 19388 39546 19400
rect 25792 19332 26648 19360
rect 15344 19264 15516 19292
rect 15344 19252 15350 19264
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 16025 19295 16083 19301
rect 16025 19292 16037 19295
rect 15620 19264 16037 19292
rect 15620 19252 15626 19264
rect 16025 19261 16037 19264
rect 16071 19261 16083 19295
rect 16025 19255 16083 19261
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 16172 19264 17417 19292
rect 16172 19252 16178 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 18598 19252 18604 19304
rect 18656 19252 18662 19304
rect 19794 19252 19800 19304
rect 19852 19252 19858 19304
rect 20073 19295 20131 19301
rect 20073 19261 20085 19295
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 20441 19295 20499 19301
rect 20441 19261 20453 19295
rect 20487 19292 20499 19295
rect 20898 19292 20904 19304
rect 20487 19264 20904 19292
rect 20487 19261 20499 19264
rect 20441 19255 20499 19261
rect 15930 19224 15936 19236
rect 12308 19196 13216 19224
rect 14936 19196 15936 19224
rect 12308 19184 12314 19196
rect 5810 19116 5816 19168
rect 5868 19116 5874 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 11882 19156 11888 19168
rect 8352 19128 11888 19156
rect 8352 19116 8358 19128
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12710 19116 12716 19168
rect 12768 19116 12774 19168
rect 13188 19156 13216 19196
rect 15930 19184 15936 19196
rect 15988 19184 15994 19236
rect 14458 19156 14464 19168
rect 13188 19128 14464 19156
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19156 14887 19159
rect 15286 19156 15292 19168
rect 14875 19128 15292 19156
rect 14875 19125 14887 19128
rect 14829 19119 14887 19125
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 19610 19116 19616 19168
rect 19668 19156 19674 19168
rect 20088 19156 20116 19255
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 21407 19264 22094 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 20622 19184 20628 19236
rect 20680 19224 20686 19236
rect 21542 19224 21548 19236
rect 20680 19196 21548 19224
rect 20680 19184 20686 19196
rect 21542 19184 21548 19196
rect 21600 19184 21606 19236
rect 19668 19128 20116 19156
rect 19668 19116 19674 19128
rect 20438 19116 20444 19168
rect 20496 19156 20502 19168
rect 20717 19159 20775 19165
rect 20717 19156 20729 19159
rect 20496 19128 20729 19156
rect 20496 19116 20502 19128
rect 20717 19125 20729 19128
rect 20763 19125 20775 19159
rect 22066 19156 22094 19264
rect 22186 19252 22192 19304
rect 22244 19252 22250 19304
rect 24854 19252 24860 19304
rect 24912 19292 24918 19304
rect 24949 19295 25007 19301
rect 24949 19292 24961 19295
rect 24912 19264 24961 19292
rect 24912 19252 24918 19264
rect 24949 19261 24961 19264
rect 24995 19261 25007 19295
rect 25792 19292 25820 19332
rect 26436 19301 26464 19332
rect 26970 19320 26976 19372
rect 27028 19360 27034 19372
rect 27246 19360 27252 19372
rect 27028 19332 27252 19360
rect 27028 19320 27034 19332
rect 27246 19320 27252 19332
rect 27304 19320 27310 19372
rect 27617 19363 27675 19369
rect 27617 19329 27629 19363
rect 27663 19360 27675 19363
rect 28166 19360 28172 19372
rect 27663 19332 28172 19360
rect 27663 19329 27675 19332
rect 27617 19323 27675 19329
rect 28166 19320 28172 19332
rect 28224 19360 28230 19372
rect 28442 19360 28448 19372
rect 28224 19332 28448 19360
rect 28224 19320 28230 19332
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28813 19363 28871 19369
rect 28813 19329 28825 19363
rect 28859 19360 28871 19363
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 28859 19332 29745 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29932 19332 30328 19360
rect 24949 19255 25007 19261
rect 25148 19264 25820 19292
rect 26421 19295 26479 19301
rect 22646 19184 22652 19236
rect 22704 19224 22710 19236
rect 22704 19196 23980 19224
rect 22704 19184 22710 19196
rect 23477 19159 23535 19165
rect 23477 19156 23489 19159
rect 22066 19128 23489 19156
rect 20717 19119 20775 19125
rect 23477 19125 23489 19128
rect 23523 19156 23535 19159
rect 23842 19156 23848 19168
rect 23523 19128 23848 19156
rect 23523 19125 23535 19128
rect 23477 19119 23535 19125
rect 23842 19116 23848 19128
rect 23900 19116 23906 19168
rect 23952 19156 23980 19196
rect 25148 19156 25176 19264
rect 26421 19261 26433 19295
rect 26467 19261 26479 19295
rect 26421 19255 26479 19261
rect 27709 19295 27767 19301
rect 27709 19261 27721 19295
rect 27755 19261 27767 19295
rect 27709 19255 27767 19261
rect 27893 19295 27951 19301
rect 27893 19261 27905 19295
rect 27939 19292 27951 19295
rect 27982 19292 27988 19304
rect 27939 19264 27988 19292
rect 27939 19261 27951 19264
rect 27893 19255 27951 19261
rect 25866 19184 25872 19236
rect 25924 19224 25930 19236
rect 27724 19224 27752 19255
rect 27982 19252 27988 19264
rect 28040 19252 28046 19304
rect 28350 19252 28356 19304
rect 28408 19292 28414 19304
rect 28905 19295 28963 19301
rect 28905 19292 28917 19295
rect 28408 19264 28917 19292
rect 28408 19252 28414 19264
rect 28905 19261 28917 19264
rect 28951 19261 28963 19295
rect 28905 19255 28963 19261
rect 28994 19252 29000 19304
rect 29052 19252 29058 19304
rect 29086 19252 29092 19304
rect 29144 19292 29150 19304
rect 29932 19292 29960 19332
rect 29144 19264 29960 19292
rect 30300 19292 30328 19332
rect 30374 19320 30380 19372
rect 30432 19360 30438 19372
rect 30745 19363 30803 19369
rect 30745 19360 30757 19363
rect 30432 19332 30757 19360
rect 30432 19320 30438 19332
rect 30745 19329 30757 19332
rect 30791 19329 30803 19363
rect 30745 19323 30803 19329
rect 32582 19320 32588 19372
rect 32640 19320 32646 19372
rect 33873 19363 33931 19369
rect 33873 19329 33885 19363
rect 33919 19360 33931 19363
rect 34146 19360 34152 19372
rect 33919 19332 34152 19360
rect 33919 19329 33931 19332
rect 33873 19323 33931 19329
rect 34146 19320 34152 19332
rect 34204 19320 34210 19372
rect 34808 19332 35112 19360
rect 30466 19292 30472 19304
rect 30300 19264 30472 19292
rect 29144 19252 29150 19264
rect 30466 19252 30472 19264
rect 30524 19252 30530 19304
rect 32490 19252 32496 19304
rect 32548 19252 32554 19304
rect 33689 19295 33747 19301
rect 33689 19261 33701 19295
rect 33735 19292 33747 19295
rect 34808 19292 34836 19332
rect 33735 19264 34836 19292
rect 34885 19295 34943 19301
rect 33735 19261 33747 19264
rect 33689 19255 33747 19261
rect 34885 19261 34897 19295
rect 34931 19261 34943 19295
rect 34885 19255 34943 19261
rect 28534 19224 28540 19236
rect 25924 19196 27660 19224
rect 27724 19196 28540 19224
rect 25924 19184 25930 19196
rect 23952 19128 25176 19156
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 27246 19116 27252 19168
rect 27304 19116 27310 19168
rect 27632 19156 27660 19196
rect 28534 19184 28540 19196
rect 28592 19224 28598 19236
rect 31018 19224 31024 19236
rect 28592 19196 31024 19224
rect 28592 19184 28598 19196
rect 31018 19184 31024 19196
rect 31076 19184 31082 19236
rect 34238 19184 34244 19236
rect 34296 19184 34302 19236
rect 34900 19224 34928 19255
rect 34974 19252 34980 19304
rect 35032 19252 35038 19304
rect 35084 19292 35112 19332
rect 35912 19332 36124 19360
rect 35912 19292 35940 19332
rect 35084 19264 35940 19292
rect 35986 19252 35992 19304
rect 36044 19252 36050 19304
rect 36096 19292 36124 19332
rect 36262 19320 36268 19372
rect 36320 19320 36326 19372
rect 39684 19369 39712 19400
rect 40497 19397 40509 19431
rect 40543 19428 40555 19431
rect 48406 19428 48412 19440
rect 40543 19400 48412 19428
rect 40543 19397 40555 19400
rect 40497 19391 40555 19397
rect 48406 19388 48412 19400
rect 48464 19388 48470 19440
rect 39669 19363 39727 19369
rect 39669 19329 39681 19363
rect 39715 19329 39727 19363
rect 39669 19323 39727 19329
rect 48593 19363 48651 19369
rect 48593 19329 48605 19363
rect 48639 19360 48651 19363
rect 49234 19360 49240 19372
rect 48639 19332 49240 19360
rect 48639 19329 48651 19332
rect 48593 19323 48651 19329
rect 49234 19320 49240 19332
rect 49292 19320 49298 19372
rect 37274 19292 37280 19304
rect 36096 19264 37280 19292
rect 37274 19252 37280 19264
rect 37332 19252 37338 19304
rect 39390 19252 39396 19304
rect 39448 19252 39454 19304
rect 40681 19295 40739 19301
rect 40681 19292 40693 19295
rect 39592 19264 40693 19292
rect 37366 19224 37372 19236
rect 34900 19196 37372 19224
rect 37366 19184 37372 19196
rect 37424 19224 37430 19236
rect 37734 19224 37740 19236
rect 37424 19196 37740 19224
rect 37424 19184 37430 19196
rect 37734 19184 37740 19196
rect 37792 19224 37798 19236
rect 37792 19196 38056 19224
rect 37792 19184 37798 19196
rect 29270 19156 29276 19168
rect 27632 19128 29276 19156
rect 29270 19116 29276 19128
rect 29328 19116 29334 19168
rect 30098 19116 30104 19168
rect 30156 19156 30162 19168
rect 30193 19159 30251 19165
rect 30193 19156 30205 19159
rect 30156 19128 30205 19156
rect 30156 19116 30162 19128
rect 30193 19125 30205 19128
rect 30239 19125 30251 19159
rect 30193 19119 30251 19125
rect 30374 19116 30380 19168
rect 30432 19116 30438 19168
rect 33962 19116 33968 19168
rect 34020 19156 34026 19168
rect 35066 19156 35072 19168
rect 34020 19128 35072 19156
rect 34020 19116 34026 19128
rect 35066 19116 35072 19128
rect 35124 19116 35130 19168
rect 36630 19116 36636 19168
rect 36688 19116 36694 19168
rect 36906 19116 36912 19168
rect 36964 19116 36970 19168
rect 37826 19116 37832 19168
rect 37884 19156 37890 19168
rect 37921 19159 37979 19165
rect 37921 19156 37933 19159
rect 37884 19128 37933 19156
rect 37884 19116 37890 19128
rect 37921 19125 37933 19128
rect 37967 19125 37979 19159
rect 38028 19156 38056 19196
rect 39592 19156 39620 19264
rect 40681 19261 40693 19264
rect 40727 19261 40739 19295
rect 40681 19255 40739 19261
rect 41046 19252 41052 19304
rect 41104 19292 41110 19304
rect 42058 19292 42064 19304
rect 41104 19264 42064 19292
rect 41104 19252 41110 19264
rect 42058 19252 42064 19264
rect 42116 19252 42122 19304
rect 40218 19184 40224 19236
rect 40276 19224 40282 19236
rect 49053 19227 49111 19233
rect 49053 19224 49065 19227
rect 40276 19196 49065 19224
rect 40276 19184 40282 19196
rect 49053 19193 49065 19196
rect 49099 19193 49111 19227
rect 49053 19187 49111 19193
rect 38028 19128 39620 19156
rect 37921 19119 37979 19125
rect 40034 19116 40040 19168
rect 40092 19156 40098 19168
rect 41046 19156 41052 19168
rect 40092 19128 41052 19156
rect 40092 19116 40098 19128
rect 41046 19116 41052 19128
rect 41104 19156 41110 19168
rect 41141 19159 41199 19165
rect 41141 19156 41153 19159
rect 41104 19128 41153 19156
rect 41104 19116 41110 19128
rect 41141 19125 41153 19128
rect 41187 19125 41199 19159
rect 41141 19119 41199 19125
rect 48777 19159 48835 19165
rect 48777 19125 48789 19159
rect 48823 19156 48835 19159
rect 49418 19156 49424 19168
rect 48823 19128 49424 19156
rect 48823 19125 48835 19128
rect 48777 19119 48835 19125
rect 49418 19116 49424 19128
rect 49476 19116 49482 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 6880 18924 9229 18952
rect 6880 18912 6886 18924
rect 9217 18921 9229 18924
rect 9263 18952 9275 18955
rect 10962 18952 10968 18964
rect 9263 18924 10968 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 10962 18912 10968 18924
rect 11020 18912 11026 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11112 18924 11560 18952
rect 11112 18912 11118 18924
rect 11146 18884 11152 18896
rect 10888 18856 11152 18884
rect 3510 18776 3516 18828
rect 3568 18816 3574 18828
rect 4157 18819 4215 18825
rect 4157 18816 4169 18819
rect 3568 18788 4169 18816
rect 3568 18776 3574 18788
rect 4157 18785 4169 18788
rect 4203 18785 4215 18819
rect 10888 18816 10916 18856
rect 11146 18844 11152 18856
rect 11204 18844 11210 18896
rect 11532 18884 11560 18924
rect 11882 18912 11888 18964
rect 11940 18912 11946 18964
rect 14292 18924 15884 18952
rect 12526 18884 12532 18896
rect 11532 18856 12532 18884
rect 12526 18844 12532 18856
rect 12584 18844 12590 18896
rect 12710 18844 12716 18896
rect 12768 18884 12774 18896
rect 12768 18856 13124 18884
rect 12768 18844 12774 18856
rect 13096 18825 13124 18856
rect 13354 18844 13360 18896
rect 13412 18884 13418 18896
rect 13630 18884 13636 18896
rect 13412 18856 13636 18884
rect 13412 18844 13418 18856
rect 13630 18844 13636 18856
rect 13688 18844 13694 18896
rect 4157 18779 4215 18785
rect 8312 18788 10916 18816
rect 10965 18819 11023 18825
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18717 3019 18751
rect 2961 18711 3019 18717
rect 1394 18640 1400 18692
rect 1452 18680 1458 18692
rect 1765 18683 1823 18689
rect 1765 18680 1777 18683
rect 1452 18652 1777 18680
rect 1452 18640 1458 18652
rect 1765 18649 1777 18652
rect 1811 18649 1823 18683
rect 1765 18643 1823 18649
rect 2976 18612 3004 18711
rect 5350 18708 5356 18760
rect 5408 18708 5414 18760
rect 8312 18757 8340 18788
rect 10965 18785 10977 18819
rect 11011 18816 11023 18819
rect 13081 18819 13139 18825
rect 11011 18788 13032 18816
rect 11011 18785 11023 18788
rect 10965 18779 11023 18785
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 13004 18748 13032 18788
rect 13081 18785 13093 18819
rect 13127 18816 13139 18819
rect 13170 18816 13176 18828
rect 13127 18788 13176 18816
rect 13127 18785 13139 18788
rect 13081 18779 13139 18785
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 14292 18825 14320 18924
rect 15856 18884 15884 18924
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 16025 18955 16083 18961
rect 16025 18952 16037 18955
rect 15988 18924 16037 18952
rect 15988 18912 15994 18924
rect 16025 18921 16037 18924
rect 16071 18952 16083 18955
rect 16114 18952 16120 18964
rect 16071 18924 16120 18952
rect 16071 18921 16083 18924
rect 16025 18915 16083 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 16393 18955 16451 18961
rect 16393 18921 16405 18955
rect 16439 18952 16451 18955
rect 16666 18952 16672 18964
rect 16439 18924 16672 18952
rect 16439 18921 16451 18924
rect 16393 18915 16451 18921
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 16758 18912 16764 18964
rect 16816 18952 16822 18964
rect 16945 18955 17003 18961
rect 16945 18952 16957 18955
rect 16816 18924 16957 18952
rect 16816 18912 16822 18924
rect 16945 18921 16957 18924
rect 16991 18921 17003 18955
rect 16945 18915 17003 18921
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 18322 18952 18328 18964
rect 18187 18924 18328 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 19886 18912 19892 18964
rect 19944 18912 19950 18964
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 21048 18924 21097 18952
rect 21048 18912 21054 18924
rect 21085 18921 21097 18924
rect 21131 18921 21143 18955
rect 21085 18915 21143 18921
rect 22462 18912 22468 18964
rect 22520 18952 22526 18964
rect 27154 18952 27160 18964
rect 22520 18924 27160 18952
rect 22520 18912 22526 18924
rect 27154 18912 27160 18924
rect 27212 18912 27218 18964
rect 27525 18955 27583 18961
rect 27525 18921 27537 18955
rect 27571 18952 27583 18955
rect 29086 18952 29092 18964
rect 27571 18924 29092 18952
rect 27571 18921 27583 18924
rect 27525 18915 27583 18921
rect 29086 18912 29092 18924
rect 29144 18952 29150 18964
rect 30282 18952 30288 18964
rect 29144 18924 30288 18952
rect 29144 18912 29150 18924
rect 30282 18912 30288 18924
rect 30340 18912 30346 18964
rect 30650 18912 30656 18964
rect 30708 18952 30714 18964
rect 31481 18955 31539 18961
rect 31481 18952 31493 18955
rect 30708 18924 31493 18952
rect 30708 18912 30714 18924
rect 31481 18921 31493 18924
rect 31527 18921 31539 18955
rect 36078 18952 36084 18964
rect 31481 18915 31539 18921
rect 33520 18924 36084 18952
rect 16298 18884 16304 18896
rect 15856 18856 16304 18884
rect 16298 18844 16304 18856
rect 16356 18844 16362 18896
rect 16574 18844 16580 18896
rect 16632 18884 16638 18896
rect 20806 18884 20812 18896
rect 16632 18856 17540 18884
rect 16632 18844 16638 18856
rect 17512 18825 17540 18856
rect 18616 18856 20812 18884
rect 18616 18825 18644 18856
rect 20806 18844 20812 18856
rect 20864 18844 20870 18896
rect 24320 18856 25912 18884
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18785 14335 18819
rect 14277 18779 14335 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 19426 18816 19432 18828
rect 18831 18788 19432 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 20162 18776 20168 18828
rect 20220 18816 20226 18828
rect 20441 18819 20499 18825
rect 20441 18816 20453 18819
rect 20220 18788 20453 18816
rect 20220 18776 20226 18788
rect 20441 18785 20453 18788
rect 20487 18785 20499 18819
rect 20441 18779 20499 18785
rect 21174 18776 21180 18828
rect 21232 18816 21238 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21232 18788 21649 18816
rect 21232 18776 21238 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 21637 18779 21695 18785
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22281 18819 22339 18825
rect 22281 18816 22293 18819
rect 22152 18788 22293 18816
rect 22152 18776 22158 18788
rect 22281 18785 22293 18788
rect 22327 18816 22339 18819
rect 24320 18816 24348 18856
rect 22327 18788 24348 18816
rect 22327 18785 22339 18788
rect 22281 18779 22339 18785
rect 25038 18776 25044 18828
rect 25096 18776 25102 18828
rect 25240 18825 25268 18856
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 25740 18788 25789 18816
rect 25740 18776 25746 18788
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 25884 18816 25912 18856
rect 27982 18844 27988 18896
rect 28040 18884 28046 18896
rect 28169 18887 28227 18893
rect 28169 18884 28181 18887
rect 28040 18856 28181 18884
rect 28040 18844 28046 18856
rect 28169 18853 28181 18856
rect 28215 18884 28227 18887
rect 28902 18884 28908 18896
rect 28215 18856 28908 18884
rect 28215 18853 28227 18856
rect 28169 18847 28227 18853
rect 28902 18844 28908 18856
rect 28960 18844 28966 18896
rect 28994 18844 29000 18896
rect 29052 18844 29058 18896
rect 30098 18884 30104 18896
rect 29288 18856 30104 18884
rect 27522 18816 27528 18828
rect 25884 18788 27528 18816
rect 25777 18779 25835 18785
rect 27522 18776 27528 18788
rect 27580 18776 27586 18828
rect 27706 18776 27712 18828
rect 27764 18816 27770 18828
rect 28077 18819 28135 18825
rect 28077 18816 28089 18819
rect 27764 18788 28089 18816
rect 27764 18776 27770 18788
rect 28077 18785 28089 18788
rect 28123 18816 28135 18819
rect 29288 18816 29316 18856
rect 30098 18844 30104 18856
rect 30156 18844 30162 18896
rect 30926 18844 30932 18896
rect 30984 18844 30990 18896
rect 33413 18887 33471 18893
rect 33413 18853 33425 18887
rect 33459 18884 33471 18887
rect 33520 18884 33548 18924
rect 36078 18912 36084 18924
rect 36136 18912 36142 18964
rect 37369 18955 37427 18961
rect 37369 18921 37381 18955
rect 37415 18952 37427 18955
rect 39390 18952 39396 18964
rect 37415 18924 39396 18952
rect 37415 18921 37427 18924
rect 37369 18915 37427 18921
rect 39390 18912 39396 18924
rect 39448 18912 39454 18964
rect 42058 18912 42064 18964
rect 42116 18912 42122 18964
rect 33459 18856 33548 18884
rect 33459 18853 33471 18856
rect 33413 18847 33471 18853
rect 33594 18844 33600 18896
rect 33652 18884 33658 18896
rect 34149 18887 34207 18893
rect 34149 18884 34161 18887
rect 33652 18856 34161 18884
rect 33652 18844 33658 18856
rect 34149 18853 34161 18856
rect 34195 18884 34207 18887
rect 34238 18884 34244 18896
rect 34195 18856 34244 18884
rect 34195 18853 34207 18856
rect 34149 18847 34207 18853
rect 34238 18844 34244 18856
rect 34296 18844 34302 18896
rect 34514 18844 34520 18896
rect 34572 18844 34578 18896
rect 37182 18844 37188 18896
rect 37240 18884 37246 18896
rect 37734 18884 37740 18896
rect 37240 18856 37740 18884
rect 37240 18844 37246 18856
rect 37734 18844 37740 18856
rect 37792 18844 37798 18896
rect 38010 18844 38016 18896
rect 38068 18844 38074 18896
rect 42702 18844 42708 18896
rect 42760 18884 42766 18896
rect 49145 18887 49203 18893
rect 49145 18884 49157 18887
rect 42760 18856 49157 18884
rect 42760 18844 42766 18856
rect 49145 18853 49157 18856
rect 49191 18853 49203 18887
rect 49145 18847 49203 18853
rect 28123 18788 29316 18816
rect 28123 18785 28135 18788
rect 28077 18779 28135 18785
rect 29546 18776 29552 18828
rect 29604 18816 29610 18828
rect 29825 18819 29883 18825
rect 29825 18816 29837 18819
rect 29604 18788 29837 18816
rect 29604 18776 29610 18788
rect 29825 18785 29837 18788
rect 29871 18785 29883 18819
rect 29825 18779 29883 18785
rect 29914 18776 29920 18828
rect 29972 18816 29978 18828
rect 30009 18819 30067 18825
rect 30009 18816 30021 18819
rect 29972 18788 30021 18816
rect 29972 18776 29978 18788
rect 30009 18785 30021 18788
rect 30055 18816 30067 18819
rect 30650 18816 30656 18828
rect 30055 18788 30656 18816
rect 30055 18785 30067 18788
rect 30009 18779 30067 18785
rect 30650 18776 30656 18788
rect 30708 18776 30714 18828
rect 32125 18819 32183 18825
rect 32125 18785 32137 18819
rect 32171 18785 32183 18819
rect 32125 18779 32183 18785
rect 13446 18748 13452 18760
rect 12115 18720 12756 18748
rect 13004 18720 13452 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 8113 18683 8171 18689
rect 8113 18680 8125 18683
rect 4396 18652 8125 18680
rect 4396 18640 4402 18652
rect 8113 18649 8125 18652
rect 8159 18649 8171 18683
rect 8113 18643 8171 18649
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10284 18652 10640 18680
rect 10284 18640 10290 18652
rect 7834 18612 7840 18624
rect 2976 18584 7840 18612
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 10612 18612 10640 18652
rect 10686 18640 10692 18692
rect 10744 18640 10750 18692
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 10612 18584 11345 18612
rect 11333 18581 11345 18584
rect 11379 18612 11391 18615
rect 11609 18615 11667 18621
rect 11609 18612 11621 18615
rect 11379 18584 11621 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11609 18581 11621 18584
rect 11655 18612 11667 18615
rect 11974 18612 11980 18624
rect 11655 18584 11980 18612
rect 11655 18581 11667 18584
rect 11609 18575 11667 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12342 18572 12348 18624
rect 12400 18612 12406 18624
rect 12529 18615 12587 18621
rect 12529 18612 12541 18615
rect 12400 18584 12541 18612
rect 12400 18572 12406 18584
rect 12529 18581 12541 18584
rect 12575 18581 12587 18615
rect 12728 18612 12756 18720
rect 13446 18708 13452 18720
rect 13504 18708 13510 18760
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 16666 18748 16672 18760
rect 15712 18720 16672 18748
rect 15712 18708 15718 18720
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 22002 18748 22008 18760
rect 18564 18720 22008 18748
rect 18564 18708 18570 18720
rect 22002 18708 22008 18720
rect 22060 18708 22066 18760
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18748 24087 18751
rect 24118 18748 24124 18760
rect 24075 18720 24124 18748
rect 24075 18717 24087 18720
rect 24029 18711 24087 18717
rect 24118 18708 24124 18720
rect 24176 18748 24182 18760
rect 25700 18748 25728 18776
rect 24176 18720 25728 18748
rect 27893 18751 27951 18757
rect 24176 18708 24182 18720
rect 27893 18717 27905 18751
rect 27939 18748 27951 18751
rect 28810 18748 28816 18760
rect 27939 18720 28816 18748
rect 27939 18717 27951 18720
rect 27893 18711 27951 18717
rect 28810 18708 28816 18720
rect 28868 18708 28874 18760
rect 29181 18751 29239 18757
rect 29181 18717 29193 18751
rect 29227 18717 29239 18751
rect 29181 18711 29239 18717
rect 12802 18640 12808 18692
rect 12860 18680 12866 18692
rect 12897 18683 12955 18689
rect 12897 18680 12909 18683
rect 12860 18652 12909 18680
rect 12860 18640 12866 18652
rect 12897 18649 12909 18652
rect 12943 18649 12955 18683
rect 12897 18643 12955 18649
rect 12989 18683 13047 18689
rect 12989 18649 13001 18683
rect 13035 18680 13047 18683
rect 13035 18652 14504 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 13262 18612 13268 18624
rect 12728 18584 13268 18612
rect 12529 18575 12587 18581
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 13906 18572 13912 18624
rect 13964 18572 13970 18624
rect 14476 18612 14504 18652
rect 14550 18640 14556 18692
rect 14608 18640 14614 18692
rect 17402 18640 17408 18692
rect 17460 18640 17466 18692
rect 19334 18640 19340 18692
rect 19392 18640 19398 18692
rect 20257 18683 20315 18689
rect 20257 18649 20269 18683
rect 20303 18680 20315 18683
rect 20303 18652 22508 18680
rect 20303 18649 20315 18652
rect 20257 18643 20315 18649
rect 15562 18612 15568 18624
rect 14476 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 16669 18615 16727 18621
rect 16669 18581 16681 18615
rect 16715 18612 16727 18615
rect 16758 18612 16764 18624
rect 16715 18584 16764 18612
rect 16715 18581 16727 18584
rect 16669 18575 16727 18581
rect 16758 18572 16764 18584
rect 16816 18612 16822 18624
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 16816 18584 17325 18612
rect 16816 18572 16822 18584
rect 17313 18581 17325 18584
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 18414 18572 18420 18624
rect 18472 18612 18478 18624
rect 18509 18615 18567 18621
rect 18509 18612 18521 18615
rect 18472 18584 18521 18612
rect 18472 18572 18478 18584
rect 18509 18581 18521 18584
rect 18555 18581 18567 18615
rect 18509 18575 18567 18581
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 19518 18612 19524 18624
rect 18656 18584 19524 18612
rect 18656 18572 18662 18584
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 19610 18572 19616 18624
rect 19668 18572 19674 18624
rect 20346 18572 20352 18624
rect 20404 18572 20410 18624
rect 21450 18572 21456 18624
rect 21508 18572 21514 18624
rect 21545 18615 21603 18621
rect 21545 18581 21557 18615
rect 21591 18612 21603 18615
rect 21910 18612 21916 18624
rect 21591 18584 21916 18612
rect 21591 18581 21603 18584
rect 21545 18575 21603 18581
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 22480 18612 22508 18652
rect 22738 18640 22744 18692
rect 22796 18640 22802 18692
rect 23474 18640 23480 18692
rect 23532 18680 23538 18692
rect 23753 18683 23811 18689
rect 23753 18680 23765 18683
rect 23532 18652 23765 18680
rect 23532 18640 23538 18652
rect 23753 18649 23765 18652
rect 23799 18649 23811 18683
rect 23753 18643 23811 18649
rect 23842 18640 23848 18692
rect 23900 18680 23906 18692
rect 26053 18683 26111 18689
rect 26053 18680 26065 18683
rect 23900 18652 26065 18680
rect 23900 18640 23906 18652
rect 26053 18649 26065 18652
rect 26099 18649 26111 18683
rect 27430 18680 27436 18692
rect 27278 18652 27436 18680
rect 26053 18643 26111 18649
rect 27430 18640 27436 18652
rect 27488 18640 27494 18692
rect 27522 18640 27528 18692
rect 27580 18680 27586 18692
rect 29196 18680 29224 18711
rect 29454 18708 29460 18760
rect 29512 18748 29518 18760
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 29512 18720 30113 18748
rect 29512 18708 29518 18720
rect 30101 18717 30113 18720
rect 30147 18717 30159 18751
rect 32140 18748 32168 18779
rect 32766 18776 32772 18828
rect 32824 18776 32830 18828
rect 32950 18776 32956 18828
rect 33008 18776 33014 18828
rect 33042 18776 33048 18828
rect 33100 18816 33106 18828
rect 33873 18819 33931 18825
rect 33873 18816 33885 18819
rect 33100 18788 33885 18816
rect 33100 18776 33106 18788
rect 33873 18785 33885 18788
rect 33919 18785 33931 18819
rect 33873 18779 33931 18785
rect 34054 18776 34060 18828
rect 34112 18816 34118 18828
rect 35621 18819 35679 18825
rect 35621 18816 35633 18819
rect 34112 18788 35633 18816
rect 34112 18776 34118 18788
rect 35621 18785 35633 18788
rect 35667 18785 35679 18819
rect 35621 18779 35679 18785
rect 37090 18776 37096 18828
rect 37148 18816 37154 18828
rect 37918 18816 37924 18828
rect 37148 18788 37924 18816
rect 37148 18776 37154 18788
rect 37918 18776 37924 18788
rect 37976 18776 37982 18828
rect 38562 18776 38568 18828
rect 38620 18776 38626 18828
rect 41785 18819 41843 18825
rect 41785 18816 41797 18819
rect 39776 18788 41797 18816
rect 35342 18748 35348 18760
rect 32140 18720 35348 18748
rect 30101 18711 30159 18717
rect 35342 18708 35348 18720
rect 35400 18748 35406 18760
rect 35400 18720 35664 18748
rect 35400 18708 35406 18720
rect 35526 18680 35532 18692
rect 27580 18652 28672 18680
rect 29196 18652 35532 18680
rect 27580 18640 27586 18652
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 22480 18584 24593 18612
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 24762 18572 24768 18624
rect 24820 18612 24826 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24820 18584 24961 18612
rect 24820 18572 24826 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 26786 18572 26792 18624
rect 26844 18612 26850 18624
rect 27982 18612 27988 18624
rect 26844 18584 27988 18612
rect 26844 18572 26850 18584
rect 27982 18572 27988 18584
rect 28040 18572 28046 18624
rect 28166 18572 28172 18624
rect 28224 18612 28230 18624
rect 28353 18615 28411 18621
rect 28353 18612 28365 18615
rect 28224 18584 28365 18612
rect 28224 18572 28230 18584
rect 28353 18581 28365 18584
rect 28399 18581 28411 18615
rect 28353 18575 28411 18581
rect 28442 18572 28448 18624
rect 28500 18612 28506 18624
rect 28537 18615 28595 18621
rect 28537 18612 28549 18615
rect 28500 18584 28549 18612
rect 28500 18572 28506 18584
rect 28537 18581 28549 18584
rect 28583 18581 28595 18615
rect 28644 18612 28672 18652
rect 35526 18640 35532 18652
rect 35584 18640 35590 18692
rect 35636 18680 35664 18720
rect 35897 18683 35955 18689
rect 35897 18680 35909 18683
rect 35636 18652 35909 18680
rect 35897 18649 35909 18652
rect 35943 18649 35955 18683
rect 37108 18666 37136 18776
rect 37642 18708 37648 18760
rect 37700 18748 37706 18760
rect 38381 18751 38439 18757
rect 38381 18748 38393 18751
rect 37700 18720 38393 18748
rect 37700 18708 37706 18720
rect 38381 18717 38393 18720
rect 38427 18717 38439 18751
rect 38381 18711 38439 18717
rect 39776 18692 39804 18788
rect 41785 18785 41797 18788
rect 41831 18785 41843 18819
rect 41785 18779 41843 18785
rect 40034 18708 40040 18760
rect 40092 18748 40098 18760
rect 48593 18751 48651 18757
rect 40092 18720 40434 18748
rect 40092 18708 40098 18720
rect 48593 18717 48605 18751
rect 48639 18748 48651 18751
rect 48774 18748 48780 18760
rect 48639 18720 48780 18748
rect 48639 18717 48651 18720
rect 48593 18711 48651 18717
rect 48774 18708 48780 18720
rect 48832 18708 48838 18760
rect 49329 18751 49387 18757
rect 49329 18717 49341 18751
rect 49375 18748 49387 18751
rect 49418 18748 49424 18760
rect 49375 18720 49424 18748
rect 49375 18717 49387 18720
rect 49329 18711 49387 18717
rect 49418 18708 49424 18720
rect 49476 18708 49482 18760
rect 39577 18683 39635 18689
rect 39577 18680 39589 18683
rect 35897 18643 35955 18649
rect 37660 18652 39589 18680
rect 29362 18612 29368 18624
rect 28644 18584 29368 18612
rect 28537 18575 28595 18581
rect 29362 18572 29368 18584
rect 29420 18572 29426 18624
rect 30466 18572 30472 18624
rect 30524 18572 30530 18624
rect 30650 18572 30656 18624
rect 30708 18612 30714 18624
rect 30837 18615 30895 18621
rect 30837 18612 30849 18615
rect 30708 18584 30849 18612
rect 30708 18572 30714 18584
rect 30837 18581 30849 18584
rect 30883 18612 30895 18615
rect 30926 18612 30932 18624
rect 30883 18584 30932 18612
rect 30883 18581 30895 18584
rect 30837 18575 30895 18581
rect 30926 18572 30932 18584
rect 30984 18572 30990 18624
rect 31205 18615 31263 18621
rect 31205 18581 31217 18615
rect 31251 18612 31263 18615
rect 31386 18612 31392 18624
rect 31251 18584 31392 18612
rect 31251 18581 31263 18584
rect 31205 18575 31263 18581
rect 31386 18572 31392 18584
rect 31444 18572 31450 18624
rect 31662 18572 31668 18624
rect 31720 18612 31726 18624
rect 31849 18615 31907 18621
rect 31849 18612 31861 18615
rect 31720 18584 31861 18612
rect 31720 18572 31726 18584
rect 31849 18581 31861 18584
rect 31895 18581 31907 18615
rect 31849 18575 31907 18581
rect 31938 18572 31944 18624
rect 31996 18572 32002 18624
rect 32030 18572 32036 18624
rect 32088 18612 32094 18624
rect 33045 18615 33103 18621
rect 33045 18612 33057 18615
rect 32088 18584 33057 18612
rect 32088 18572 32094 18584
rect 33045 18581 33057 18584
rect 33091 18612 33103 18615
rect 33689 18615 33747 18621
rect 33689 18612 33701 18615
rect 33091 18584 33701 18612
rect 33091 18581 33103 18584
rect 33045 18575 33103 18581
rect 33689 18581 33701 18584
rect 33735 18581 33747 18615
rect 33689 18575 33747 18581
rect 34146 18572 34152 18624
rect 34204 18612 34210 18624
rect 34241 18615 34299 18621
rect 34241 18612 34253 18615
rect 34204 18584 34253 18612
rect 34204 18572 34210 18584
rect 34241 18581 34253 18584
rect 34287 18581 34299 18615
rect 34241 18575 34299 18581
rect 35161 18615 35219 18621
rect 35161 18581 35173 18615
rect 35207 18612 35219 18615
rect 36262 18612 36268 18624
rect 35207 18584 36268 18612
rect 35207 18581 35219 18584
rect 35161 18575 35219 18581
rect 36262 18572 36268 18584
rect 36320 18572 36326 18624
rect 37550 18572 37556 18624
rect 37608 18612 37614 18624
rect 37660 18621 37688 18652
rect 39577 18649 39589 18652
rect 39623 18680 39635 18683
rect 39758 18680 39764 18692
rect 39623 18652 39764 18680
rect 39623 18649 39635 18652
rect 39577 18643 39635 18649
rect 39758 18640 39764 18652
rect 39816 18640 39822 18692
rect 41509 18683 41567 18689
rect 41509 18680 41521 18683
rect 41386 18652 41521 18680
rect 37645 18615 37703 18621
rect 37645 18612 37657 18615
rect 37608 18584 37657 18612
rect 37608 18572 37614 18584
rect 37645 18581 37657 18584
rect 37691 18581 37703 18615
rect 37645 18575 37703 18581
rect 38473 18615 38531 18621
rect 38473 18581 38485 18615
rect 38519 18612 38531 18615
rect 39942 18612 39948 18624
rect 38519 18584 39948 18612
rect 38519 18581 38531 18584
rect 38473 18575 38531 18581
rect 39942 18572 39948 18584
rect 40000 18572 40006 18624
rect 40037 18615 40095 18621
rect 40037 18581 40049 18615
rect 40083 18612 40095 18615
rect 40126 18612 40132 18624
rect 40083 18584 40132 18612
rect 40083 18581 40095 18584
rect 40037 18575 40095 18581
rect 40126 18572 40132 18584
rect 40184 18572 40190 18624
rect 40218 18572 40224 18624
rect 40276 18612 40282 18624
rect 41386 18612 41414 18652
rect 41509 18649 41521 18652
rect 41555 18649 41567 18683
rect 41509 18643 41567 18649
rect 40276 18584 41414 18612
rect 40276 18572 40282 18584
rect 48406 18572 48412 18624
rect 48464 18572 48470 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 3602 18368 3608 18420
rect 3660 18368 3666 18420
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18377 9827 18411
rect 9769 18371 9827 18377
rect 4154 18340 4160 18352
rect 3436 18312 4160 18340
rect 3436 18281 3464 18312
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 5626 18300 5632 18352
rect 5684 18340 5690 18352
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 5684 18312 7665 18340
rect 5684 18300 5690 18312
rect 7653 18309 7665 18312
rect 7699 18309 7711 18343
rect 9784 18340 9812 18371
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 9916 18380 10793 18408
rect 9916 18368 9922 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 10781 18371 10839 18377
rect 11790 18368 11796 18420
rect 11848 18408 11854 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 11848 18380 14289 18408
rect 11848 18368 11854 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 17957 18411 18015 18417
rect 17957 18408 17969 18411
rect 14277 18371 14335 18377
rect 15212 18380 17969 18408
rect 10042 18340 10048 18352
rect 9784 18312 10048 18340
rect 7653 18303 7711 18309
rect 10042 18300 10048 18312
rect 10100 18300 10106 18352
rect 11238 18340 11244 18352
rect 10796 18312 11244 18340
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18241 3019 18275
rect 2961 18235 3019 18241
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 1762 18164 1768 18216
rect 1820 18164 1826 18216
rect 2976 18136 3004 18235
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4120 18244 4445 18272
rect 4120 18232 4126 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18272 10011 18275
rect 10796 18272 10824 18312
rect 11238 18300 11244 18312
rect 11296 18300 11302 18352
rect 12434 18300 12440 18352
rect 12492 18300 12498 18352
rect 13170 18300 13176 18352
rect 13228 18300 13234 18352
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 15212 18340 15240 18380
rect 17957 18377 17969 18380
rect 18003 18377 18015 18411
rect 17957 18371 18015 18377
rect 19061 18411 19119 18417
rect 19061 18377 19073 18411
rect 19107 18408 19119 18411
rect 23290 18408 23296 18420
rect 19107 18380 23296 18408
rect 19107 18377 19119 18380
rect 19061 18371 19119 18377
rect 23290 18368 23296 18380
rect 23348 18368 23354 18420
rect 25774 18408 25780 18420
rect 24044 18380 25780 18408
rect 17221 18343 17279 18349
rect 17221 18340 17233 18343
rect 13320 18312 15240 18340
rect 15304 18312 17233 18340
rect 13320 18300 13326 18312
rect 9999 18244 10824 18272
rect 10873 18275 10931 18281
rect 9999 18241 10011 18244
rect 9953 18235 10011 18241
rect 10873 18241 10885 18275
rect 10919 18272 10931 18275
rect 11790 18272 11796 18284
rect 10919 18244 11796 18272
rect 10919 18241 10931 18244
rect 10873 18235 10931 18241
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4246 18204 4252 18216
rect 4203 18176 4252 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 6822 18136 6828 18148
rect 2976 18108 6828 18136
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 7852 18136 7880 18235
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 13446 18232 13452 18284
rect 13504 18232 13510 18284
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14182 18272 14188 18284
rect 13872 18244 14188 18272
rect 13872 18232 13878 18244
rect 14182 18232 14188 18244
rect 14240 18272 14246 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 14240 18244 15209 18272
rect 14240 18232 14246 18244
rect 15197 18241 15209 18244
rect 15243 18272 15255 18275
rect 15304 18272 15332 18312
rect 17221 18309 17233 18312
rect 17267 18309 17279 18343
rect 17221 18303 17279 18309
rect 17405 18343 17463 18349
rect 17405 18309 17417 18343
rect 17451 18340 17463 18343
rect 18506 18340 18512 18352
rect 17451 18312 18512 18340
rect 17451 18309 17463 18312
rect 17405 18303 17463 18309
rect 18506 18300 18512 18312
rect 18564 18300 18570 18352
rect 19150 18340 19156 18352
rect 18616 18312 19156 18340
rect 15243 18244 15332 18272
rect 16301 18275 16359 18281
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 16301 18241 16313 18275
rect 16347 18272 16359 18275
rect 18230 18272 18236 18284
rect 16347 18244 18236 18272
rect 16347 18241 16359 18244
rect 16301 18235 16359 18241
rect 18230 18232 18236 18244
rect 18288 18232 18294 18284
rect 18325 18275 18383 18281
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 18371 18244 18552 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10652 18176 10977 18204
rect 10652 18164 10658 18176
rect 10965 18173 10977 18176
rect 11011 18204 11023 18207
rect 11698 18204 11704 18216
rect 11011 18176 11704 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 14369 18207 14427 18213
rect 12584 18176 13952 18204
rect 12584 18164 12590 18176
rect 13924 18145 13952 18176
rect 14369 18173 14381 18207
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 13909 18139 13967 18145
rect 7852 18108 11836 18136
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 9824 18040 10425 18068
rect 9824 18028 9830 18040
rect 10413 18037 10425 18040
rect 10459 18037 10471 18071
rect 10413 18031 10471 18037
rect 11698 18028 11704 18080
rect 11756 18028 11762 18080
rect 11808 18068 11836 18108
rect 13909 18105 13921 18139
rect 13955 18105 13967 18139
rect 14384 18136 14412 18167
rect 14550 18164 14556 18216
rect 14608 18164 14614 18216
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16482 18204 16488 18216
rect 15703 18176 16488 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 16666 18164 16672 18216
rect 16724 18204 16730 18216
rect 17494 18204 17500 18216
rect 16724 18176 17500 18204
rect 16724 18164 16730 18176
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 18417 18207 18475 18213
rect 18417 18173 18429 18207
rect 18463 18173 18475 18207
rect 18417 18167 18475 18173
rect 14384 18108 15700 18136
rect 13909 18099 13967 18105
rect 13630 18068 13636 18080
rect 11808 18040 13636 18068
rect 13630 18028 13636 18040
rect 13688 18028 13694 18080
rect 15013 18071 15071 18077
rect 15013 18037 15025 18071
rect 15059 18068 15071 18071
rect 15102 18068 15108 18080
rect 15059 18040 15108 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15672 18068 15700 18108
rect 15746 18096 15752 18148
rect 15804 18136 15810 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15804 18108 16129 18136
rect 15804 18096 15810 18108
rect 16117 18105 16129 18108
rect 16163 18105 16175 18139
rect 16117 18099 16175 18105
rect 16298 18096 16304 18148
rect 16356 18136 16362 18148
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 16356 18108 16865 18136
rect 16356 18096 16362 18108
rect 16853 18105 16865 18108
rect 16899 18136 16911 18139
rect 18322 18136 18328 18148
rect 16899 18108 18328 18136
rect 16899 18105 16911 18108
rect 16853 18099 16911 18105
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 16574 18068 16580 18080
rect 15672 18040 16580 18068
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 18432 18068 18460 18167
rect 18524 18136 18552 18244
rect 18616 18213 18644 18312
rect 19150 18300 19156 18312
rect 19208 18340 19214 18352
rect 19889 18343 19947 18349
rect 19889 18340 19901 18343
rect 19208 18312 19901 18340
rect 19208 18300 19214 18312
rect 19889 18309 19901 18312
rect 19935 18309 19947 18343
rect 19889 18303 19947 18309
rect 19978 18300 19984 18352
rect 20036 18340 20042 18352
rect 20036 18312 20378 18340
rect 20036 18300 20042 18312
rect 21450 18300 21456 18352
rect 21508 18340 21514 18352
rect 21726 18340 21732 18352
rect 21508 18312 21732 18340
rect 21508 18300 21514 18312
rect 21726 18300 21732 18312
rect 21784 18300 21790 18352
rect 22465 18343 22523 18349
rect 22465 18309 22477 18343
rect 22511 18340 22523 18343
rect 24044 18340 24072 18380
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 27246 18408 27252 18420
rect 26283 18380 27252 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27522 18368 27528 18420
rect 27580 18368 27586 18420
rect 27617 18411 27675 18417
rect 27617 18377 27629 18411
rect 27663 18408 27675 18411
rect 27706 18408 27712 18420
rect 27663 18380 27712 18408
rect 27663 18377 27675 18380
rect 27617 18371 27675 18377
rect 27706 18368 27712 18380
rect 27764 18368 27770 18420
rect 28721 18411 28779 18417
rect 28721 18377 28733 18411
rect 28767 18408 28779 18411
rect 29730 18408 29736 18420
rect 28767 18380 29736 18408
rect 28767 18377 28779 18380
rect 28721 18371 28779 18377
rect 29730 18368 29736 18380
rect 29788 18368 29794 18420
rect 29822 18368 29828 18420
rect 29880 18408 29886 18420
rect 30377 18411 30435 18417
rect 30377 18408 30389 18411
rect 29880 18380 30389 18408
rect 29880 18368 29886 18380
rect 30377 18377 30389 18380
rect 30423 18377 30435 18411
rect 30377 18371 30435 18377
rect 30837 18411 30895 18417
rect 30837 18377 30849 18411
rect 30883 18408 30895 18411
rect 31202 18408 31208 18420
rect 30883 18380 31208 18408
rect 30883 18377 30895 18380
rect 30837 18371 30895 18377
rect 31202 18368 31208 18380
rect 31260 18368 31266 18420
rect 32306 18368 32312 18420
rect 32364 18408 32370 18420
rect 32677 18411 32735 18417
rect 32677 18408 32689 18411
rect 32364 18380 32689 18408
rect 32364 18368 32370 18380
rect 32677 18377 32689 18380
rect 32723 18408 32735 18411
rect 32950 18408 32956 18420
rect 32723 18380 32956 18408
rect 32723 18377 32735 18380
rect 32677 18371 32735 18377
rect 32950 18368 32956 18380
rect 33008 18368 33014 18420
rect 33045 18411 33103 18417
rect 33045 18377 33057 18411
rect 33091 18408 33103 18411
rect 33091 18380 35204 18408
rect 33091 18377 33103 18380
rect 33045 18371 33103 18377
rect 22511 18312 24072 18340
rect 22511 18309 22523 18312
rect 22465 18303 22523 18309
rect 24118 18300 24124 18352
rect 24176 18300 24182 18352
rect 28813 18343 28871 18349
rect 24964 18312 27568 18340
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 22603 18244 23244 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 19610 18204 19616 18216
rect 19383 18176 19616 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 22462 18204 22468 18216
rect 20404 18176 22468 18204
rect 20404 18164 20410 18176
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 22649 18207 22707 18213
rect 22649 18173 22661 18207
rect 22695 18173 22707 18207
rect 23216 18204 23244 18244
rect 23290 18232 23296 18284
rect 23348 18232 23354 18284
rect 24964 18204 24992 18312
rect 27540 18284 27568 18312
rect 28813 18309 28825 18343
rect 28859 18340 28871 18343
rect 32122 18340 32128 18352
rect 28859 18312 32128 18340
rect 28859 18309 28871 18312
rect 28813 18303 28871 18309
rect 32122 18300 32128 18312
rect 32180 18300 32186 18352
rect 35176 18340 35204 18380
rect 35342 18368 35348 18420
rect 35400 18368 35406 18420
rect 35526 18368 35532 18420
rect 35584 18408 35590 18420
rect 35897 18411 35955 18417
rect 35897 18408 35909 18411
rect 35584 18380 35909 18408
rect 35584 18368 35590 18380
rect 35897 18377 35909 18380
rect 35943 18377 35955 18411
rect 35897 18371 35955 18377
rect 36814 18368 36820 18420
rect 36872 18408 36878 18420
rect 36909 18411 36967 18417
rect 36909 18408 36921 18411
rect 36872 18380 36921 18408
rect 36872 18368 36878 18380
rect 36909 18377 36921 18380
rect 36955 18377 36967 18411
rect 36909 18371 36967 18377
rect 37277 18411 37335 18417
rect 37277 18377 37289 18411
rect 37323 18408 37335 18411
rect 37550 18408 37556 18420
rect 37323 18380 37556 18408
rect 37323 18377 37335 18380
rect 37277 18371 37335 18377
rect 37550 18368 37556 18380
rect 37608 18368 37614 18420
rect 37734 18368 37740 18420
rect 37792 18408 37798 18420
rect 40405 18411 40463 18417
rect 40405 18408 40417 18411
rect 37792 18380 40417 18408
rect 37792 18368 37798 18380
rect 40405 18377 40417 18380
rect 40451 18377 40463 18411
rect 40405 18371 40463 18377
rect 40862 18368 40868 18420
rect 40920 18368 40926 18420
rect 48774 18368 48780 18420
rect 48832 18368 48838 18420
rect 36170 18340 36176 18352
rect 35176 18312 36176 18340
rect 36170 18300 36176 18312
rect 36228 18300 36234 18352
rect 37458 18300 37464 18352
rect 37516 18340 37522 18352
rect 38010 18340 38016 18352
rect 37516 18312 38016 18340
rect 37516 18300 37522 18312
rect 38010 18300 38016 18312
rect 38068 18300 38074 18352
rect 40773 18343 40831 18349
rect 40773 18309 40785 18343
rect 40819 18340 40831 18343
rect 48406 18340 48412 18352
rect 40819 18312 48412 18340
rect 40819 18309 40831 18312
rect 40773 18303 40831 18309
rect 48406 18300 48412 18312
rect 48464 18300 48470 18352
rect 25038 18232 25044 18284
rect 25096 18232 25102 18284
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 26329 18275 26387 18281
rect 26329 18241 26341 18275
rect 26375 18272 26387 18275
rect 26375 18244 27476 18272
rect 26375 18241 26387 18244
rect 26329 18235 26387 18241
rect 23216 18176 24992 18204
rect 22649 18167 22707 18173
rect 19426 18136 19432 18148
rect 18524 18108 19432 18136
rect 19426 18096 19432 18108
rect 19484 18096 19490 18148
rect 22097 18139 22155 18145
rect 22097 18136 22109 18139
rect 20916 18108 22109 18136
rect 20916 18068 20944 18108
rect 22097 18105 22109 18108
rect 22143 18105 22155 18139
rect 22097 18099 22155 18105
rect 18432 18040 20944 18068
rect 21358 18028 21364 18080
rect 21416 18028 21422 18080
rect 21450 18028 21456 18080
rect 21508 18068 21514 18080
rect 22664 18068 22692 18167
rect 25222 18164 25228 18216
rect 25280 18164 25286 18216
rect 26418 18164 26424 18216
rect 26476 18164 26482 18216
rect 27448 18204 27476 18244
rect 27522 18232 27528 18284
rect 27580 18232 27586 18284
rect 30469 18275 30527 18281
rect 27632 18244 29868 18272
rect 27632 18204 27660 18244
rect 27448 18176 27660 18204
rect 27706 18164 27712 18216
rect 27764 18164 27770 18216
rect 28905 18207 28963 18213
rect 28905 18204 28917 18207
rect 28460 18176 28917 18204
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 24673 18139 24731 18145
rect 24673 18136 24685 18139
rect 23808 18108 24685 18136
rect 23808 18096 23814 18108
rect 24673 18105 24685 18108
rect 24719 18105 24731 18139
rect 24673 18099 24731 18105
rect 24964 18108 26004 18136
rect 21508 18040 22692 18068
rect 21508 18028 21514 18040
rect 22830 18028 22836 18080
rect 22888 18068 22894 18080
rect 24964 18068 24992 18108
rect 22888 18040 24992 18068
rect 22888 18028 22894 18040
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25869 18071 25927 18077
rect 25869 18068 25881 18071
rect 25096 18040 25881 18068
rect 25096 18028 25102 18040
rect 25869 18037 25881 18040
rect 25915 18037 25927 18071
rect 25976 18068 26004 18108
rect 26050 18096 26056 18148
rect 26108 18136 26114 18148
rect 28353 18139 28411 18145
rect 28353 18136 28365 18139
rect 26108 18108 28365 18136
rect 26108 18096 26114 18108
rect 28353 18105 28365 18108
rect 28399 18105 28411 18139
rect 28353 18099 28411 18105
rect 27062 18068 27068 18080
rect 25976 18040 27068 18068
rect 25869 18031 25927 18037
rect 27062 18028 27068 18040
rect 27120 18028 27126 18080
rect 27154 18028 27160 18080
rect 27212 18028 27218 18080
rect 27614 18028 27620 18080
rect 27672 18068 27678 18080
rect 28460 18068 28488 18176
rect 28905 18173 28917 18176
rect 28951 18173 28963 18207
rect 28905 18167 28963 18173
rect 27672 18040 28488 18068
rect 27672 18028 27678 18040
rect 29730 18028 29736 18080
rect 29788 18028 29794 18080
rect 29840 18068 29868 18244
rect 30469 18241 30481 18275
rect 30515 18272 30527 18275
rect 31297 18275 31355 18281
rect 31297 18272 31309 18275
rect 30515 18244 31309 18272
rect 30515 18241 30527 18244
rect 30469 18235 30527 18241
rect 31297 18241 31309 18244
rect 31343 18241 31355 18275
rect 33318 18272 33324 18284
rect 31297 18235 31355 18241
rect 32416 18244 33324 18272
rect 32416 18216 32444 18244
rect 33318 18232 33324 18244
rect 33376 18232 33382 18284
rect 30285 18207 30343 18213
rect 30285 18173 30297 18207
rect 30331 18173 30343 18207
rect 30285 18167 30343 18173
rect 30300 18136 30328 18167
rect 30558 18164 30564 18216
rect 30616 18204 30622 18216
rect 30926 18204 30932 18216
rect 30616 18176 30932 18204
rect 30616 18164 30622 18176
rect 30926 18164 30932 18176
rect 30984 18164 30990 18216
rect 32398 18164 32404 18216
rect 32456 18164 32462 18216
rect 32585 18207 32643 18213
rect 32585 18173 32597 18207
rect 32631 18173 32643 18207
rect 32585 18167 32643 18173
rect 30300 18108 30972 18136
rect 30742 18068 30748 18080
rect 29840 18040 30748 18068
rect 30742 18028 30748 18040
rect 30800 18028 30806 18080
rect 30944 18068 30972 18108
rect 31018 18096 31024 18148
rect 31076 18136 31082 18148
rect 32600 18136 32628 18167
rect 33594 18164 33600 18216
rect 33652 18164 33658 18216
rect 33873 18207 33931 18213
rect 33873 18173 33885 18207
rect 33919 18204 33931 18207
rect 34514 18204 34520 18216
rect 33919 18176 34520 18204
rect 33919 18173 33931 18176
rect 33873 18167 33931 18173
rect 34514 18164 34520 18176
rect 34572 18164 34578 18216
rect 31076 18108 32628 18136
rect 31076 18096 31082 18108
rect 34992 18080 35020 18258
rect 36262 18232 36268 18284
rect 36320 18232 36326 18284
rect 36357 18275 36415 18281
rect 36357 18241 36369 18275
rect 36403 18272 36415 18275
rect 37182 18272 37188 18284
rect 36403 18244 37188 18272
rect 36403 18241 36415 18244
rect 36357 18235 36415 18241
rect 37182 18232 37188 18244
rect 37240 18232 37246 18284
rect 37918 18232 37924 18284
rect 37976 18272 37982 18284
rect 37976 18244 38410 18272
rect 37976 18232 37982 18244
rect 39758 18232 39764 18284
rect 39816 18232 39822 18284
rect 48593 18275 48651 18281
rect 48593 18241 48605 18275
rect 48639 18272 48651 18275
rect 49326 18272 49332 18284
rect 48639 18244 49332 18272
rect 48639 18241 48651 18244
rect 48593 18235 48651 18241
rect 49326 18232 49332 18244
rect 49384 18232 49390 18284
rect 36541 18207 36599 18213
rect 36541 18173 36553 18207
rect 36587 18204 36599 18207
rect 37734 18204 37740 18216
rect 36587 18176 37740 18204
rect 36587 18173 36599 18176
rect 36541 18167 36599 18173
rect 37734 18164 37740 18176
rect 37792 18164 37798 18216
rect 37826 18164 37832 18216
rect 37884 18204 37890 18216
rect 39485 18207 39543 18213
rect 39485 18204 39497 18207
rect 37884 18176 39497 18204
rect 37884 18164 37890 18176
rect 39485 18173 39497 18176
rect 39531 18204 39543 18207
rect 40957 18207 41015 18213
rect 40957 18204 40969 18207
rect 39531 18176 40969 18204
rect 39531 18173 39543 18176
rect 39485 18167 39543 18173
rect 40957 18173 40969 18176
rect 41003 18173 41015 18207
rect 40957 18167 41015 18173
rect 35710 18096 35716 18148
rect 35768 18136 35774 18148
rect 36722 18136 36728 18148
rect 35768 18108 36728 18136
rect 35768 18096 35774 18108
rect 36722 18096 36728 18108
rect 36780 18096 36786 18148
rect 37090 18136 37096 18148
rect 36924 18108 37096 18136
rect 33686 18068 33692 18080
rect 30944 18040 33692 18068
rect 33686 18028 33692 18040
rect 33744 18028 33750 18080
rect 34974 18028 34980 18080
rect 35032 18068 35038 18080
rect 36538 18068 36544 18080
rect 35032 18040 36544 18068
rect 35032 18028 35038 18040
rect 36538 18028 36544 18040
rect 36596 18068 36602 18080
rect 36924 18068 36952 18108
rect 37090 18096 37096 18108
rect 37148 18136 37154 18148
rect 37553 18139 37611 18145
rect 37553 18136 37565 18139
rect 37148 18108 37565 18136
rect 37148 18096 37154 18108
rect 37553 18105 37565 18108
rect 37599 18136 37611 18139
rect 37918 18136 37924 18148
rect 37599 18108 37924 18136
rect 37599 18105 37611 18108
rect 37553 18099 37611 18105
rect 37918 18096 37924 18108
rect 37976 18096 37982 18148
rect 38010 18096 38016 18148
rect 38068 18096 38074 18148
rect 40218 18136 40224 18148
rect 39960 18108 40224 18136
rect 36596 18040 36952 18068
rect 36596 18028 36602 18040
rect 36998 18028 37004 18080
rect 37056 18068 37062 18080
rect 37274 18068 37280 18080
rect 37056 18040 37280 18068
rect 37056 18028 37062 18040
rect 37274 18028 37280 18040
rect 37332 18028 37338 18080
rect 37458 18028 37464 18080
rect 37516 18068 37522 18080
rect 37645 18071 37703 18077
rect 37645 18068 37657 18071
rect 37516 18040 37657 18068
rect 37516 18028 37522 18040
rect 37645 18037 37657 18040
rect 37691 18037 37703 18071
rect 38028 18068 38056 18096
rect 39960 18068 39988 18108
rect 40218 18096 40224 18108
rect 40276 18096 40282 18148
rect 38028 18040 39988 18068
rect 37645 18031 37703 18037
rect 40034 18028 40040 18080
rect 40092 18028 40098 18080
rect 49142 18028 49148 18080
rect 49200 18028 49206 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 10137 17867 10195 17873
rect 10137 17833 10149 17867
rect 10183 17864 10195 17867
rect 10226 17864 10232 17876
rect 10183 17836 10232 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 10594 17824 10600 17876
rect 10652 17824 10658 17876
rect 12897 17867 12955 17873
rect 12897 17833 12909 17867
rect 12943 17864 12955 17867
rect 13538 17864 13544 17876
rect 12943 17836 13544 17864
rect 12943 17833 12955 17836
rect 12897 17827 12955 17833
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 14277 17867 14335 17873
rect 14277 17833 14289 17867
rect 14323 17864 14335 17867
rect 14550 17864 14556 17876
rect 14323 17836 14556 17864
rect 14323 17833 14335 17836
rect 14277 17827 14335 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 16666 17864 16672 17876
rect 14752 17836 16672 17864
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17728 10379 17731
rect 11422 17728 11428 17740
rect 10367 17700 11428 17728
rect 10367 17697 10379 17700
rect 10321 17691 10379 17697
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 12345 17731 12403 17737
rect 12345 17697 12357 17731
rect 12391 17728 12403 17731
rect 12526 17728 12532 17740
rect 12391 17700 12532 17728
rect 12391 17697 12403 17700
rect 12345 17691 12403 17697
rect 12526 17688 12532 17700
rect 12584 17728 12590 17740
rect 13446 17728 13452 17740
rect 12584 17700 13452 17728
rect 12584 17688 12590 17700
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 14752 17728 14780 17836
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17276 17836 17509 17864
rect 17276 17824 17282 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17497 17827 17555 17833
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 19392 17836 19441 17864
rect 19392 17824 19398 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19429 17827 19487 17833
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 21082 17864 21088 17876
rect 19668 17836 21088 17864
rect 19668 17824 19674 17836
rect 19978 17796 19984 17808
rect 16776 17768 19984 17796
rect 13648 17700 14780 17728
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 10410 17660 10416 17672
rect 3007 17632 10416 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13648 17660 13676 17700
rect 15378 17688 15384 17740
rect 15436 17728 15442 17740
rect 15749 17731 15807 17737
rect 15749 17728 15761 17731
rect 15436 17700 15761 17728
rect 15436 17688 15442 17700
rect 15749 17697 15761 17700
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 16022 17688 16028 17740
rect 16080 17688 16086 17740
rect 16298 17688 16304 17740
rect 16356 17728 16362 17740
rect 16776 17728 16804 17768
rect 19978 17756 19984 17768
rect 20036 17756 20042 17808
rect 16356 17700 16804 17728
rect 16356 17688 16362 17700
rect 16850 17688 16856 17740
rect 16908 17688 16914 17740
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 18693 17731 18751 17737
rect 18693 17728 18705 17731
rect 18380 17700 18705 17728
rect 18380 17688 18386 17700
rect 18693 17697 18705 17700
rect 18739 17728 18751 17731
rect 20088 17728 20116 17836
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 21174 17824 21180 17876
rect 21232 17864 21238 17876
rect 22278 17864 22284 17876
rect 21232 17836 22284 17864
rect 21232 17824 21238 17836
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 22612 17836 23305 17864
rect 22612 17824 22618 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 23566 17824 23572 17876
rect 23624 17864 23630 17876
rect 25777 17867 25835 17873
rect 25777 17864 25789 17867
rect 23624 17836 25789 17864
rect 23624 17824 23630 17836
rect 25777 17833 25789 17836
rect 25823 17833 25835 17867
rect 25777 17827 25835 17833
rect 26234 17824 26240 17876
rect 26292 17824 26298 17876
rect 26344 17836 28764 17864
rect 22094 17756 22100 17808
rect 22152 17796 22158 17808
rect 24581 17799 24639 17805
rect 24581 17796 24593 17799
rect 22152 17768 24593 17796
rect 22152 17756 22158 17768
rect 24581 17765 24593 17768
rect 24627 17765 24639 17799
rect 24581 17759 24639 17765
rect 25222 17756 25228 17808
rect 25280 17796 25286 17808
rect 26344 17796 26372 17836
rect 25280 17768 26372 17796
rect 28736 17796 28764 17836
rect 28810 17824 28816 17876
rect 28868 17864 28874 17876
rect 29089 17867 29147 17873
rect 29089 17864 29101 17867
rect 28868 17836 29101 17864
rect 28868 17824 28874 17836
rect 29089 17833 29101 17836
rect 29135 17833 29147 17867
rect 29089 17827 29147 17833
rect 29638 17824 29644 17876
rect 29696 17824 29702 17876
rect 31478 17824 31484 17876
rect 31536 17864 31542 17876
rect 33873 17867 33931 17873
rect 33873 17864 33885 17867
rect 31536 17836 33885 17864
rect 31536 17824 31542 17836
rect 30006 17796 30012 17808
rect 28736 17768 30012 17796
rect 25280 17756 25286 17768
rect 30006 17756 30012 17768
rect 30064 17756 30070 17808
rect 18739 17700 20116 17728
rect 18739 17697 18751 17700
rect 18693 17691 18751 17697
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 21174 17728 21180 17740
rect 20312 17700 21180 17728
rect 20312 17688 20318 17700
rect 21174 17688 21180 17700
rect 21232 17688 21238 17740
rect 21634 17688 21640 17740
rect 21692 17728 21698 17740
rect 21729 17731 21787 17737
rect 21729 17728 21741 17731
rect 21692 17700 21741 17728
rect 21692 17688 21698 17700
rect 21729 17697 21741 17700
rect 21775 17697 21787 17731
rect 21729 17691 21787 17697
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22186 17728 22192 17740
rect 22051 17700 22192 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22186 17688 22192 17700
rect 22244 17688 22250 17740
rect 23937 17731 23995 17737
rect 23937 17697 23949 17731
rect 23983 17728 23995 17731
rect 24854 17728 24860 17740
rect 23983 17700 24860 17728
rect 23983 17697 23995 17700
rect 23937 17691 23995 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17697 25191 17731
rect 28442 17728 28448 17740
rect 25133 17691 25191 17697
rect 25976 17700 28448 17728
rect 13127 17632 13676 17660
rect 13725 17663 13783 17669
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13725 17629 13737 17663
rect 13771 17660 13783 17663
rect 13771 17632 14504 17660
rect 13771 17629 13783 17632
rect 13725 17623 13783 17629
rect 1026 17552 1032 17604
rect 1084 17592 1090 17604
rect 1765 17595 1823 17601
rect 1765 17592 1777 17595
rect 1084 17564 1777 17592
rect 1084 17552 1090 17564
rect 1765 17561 1777 17564
rect 1811 17561 1823 17595
rect 11974 17592 11980 17604
rect 11638 17564 11980 17592
rect 1765 17555 1823 17561
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 12066 17552 12072 17604
rect 12124 17552 12130 17604
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12084 17524 12112 17552
rect 11756 17496 12112 17524
rect 11756 17484 11762 17496
rect 13538 17484 13544 17536
rect 13596 17484 13602 17536
rect 14476 17524 14504 17632
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 16540 17632 17141 17660
rect 16540 17620 16546 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17660 18015 17663
rect 18874 17660 18880 17672
rect 18003 17632 18880 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19659 17632 20484 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 15286 17552 15292 17604
rect 15344 17592 15350 17604
rect 15654 17592 15660 17604
rect 15344 17564 15660 17592
rect 15344 17552 15350 17564
rect 15654 17552 15660 17564
rect 15712 17552 15718 17604
rect 20346 17592 20352 17604
rect 15856 17564 20352 17592
rect 15856 17524 15884 17564
rect 20346 17552 20352 17564
rect 20404 17552 20410 17604
rect 14476 17496 15884 17524
rect 15930 17484 15936 17536
rect 15988 17524 15994 17536
rect 16298 17524 16304 17536
rect 15988 17496 16304 17524
rect 15988 17484 15994 17496
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 16482 17484 16488 17536
rect 16540 17484 16546 17536
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17402 17524 17408 17536
rect 17083 17496 17408 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 20254 17524 20260 17536
rect 18656 17496 20260 17524
rect 18656 17484 18662 17496
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 20456 17524 20484 17632
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 25148 17660 25176 17691
rect 25976 17669 26004 17700
rect 28442 17688 28448 17700
rect 28500 17688 28506 17740
rect 28537 17731 28595 17737
rect 28537 17697 28549 17731
rect 28583 17728 28595 17731
rect 29086 17728 29092 17740
rect 28583 17700 29092 17728
rect 28583 17697 28595 17700
rect 28537 17691 28595 17697
rect 29086 17688 29092 17700
rect 29144 17688 29150 17740
rect 29914 17688 29920 17740
rect 29972 17728 29978 17740
rect 30282 17728 30288 17740
rect 29972 17700 30288 17728
rect 29972 17688 29978 17700
rect 30282 17688 30288 17700
rect 30340 17728 30346 17740
rect 31110 17728 31116 17740
rect 30340 17700 31116 17728
rect 30340 17688 30346 17700
rect 31110 17688 31116 17700
rect 31168 17688 31174 17740
rect 31478 17688 31484 17740
rect 31536 17688 31542 17740
rect 31588 17737 31616 17836
rect 33873 17833 33885 17836
rect 33919 17864 33931 17867
rect 38378 17864 38384 17876
rect 33919 17836 38384 17864
rect 33919 17833 33931 17836
rect 33873 17827 33931 17833
rect 38378 17824 38384 17836
rect 38436 17824 38442 17876
rect 39942 17824 39948 17876
rect 40000 17864 40006 17876
rect 40497 17867 40555 17873
rect 40497 17864 40509 17867
rect 40000 17836 40509 17864
rect 40000 17824 40006 17836
rect 40497 17833 40509 17836
rect 40543 17833 40555 17867
rect 40497 17827 40555 17833
rect 40586 17824 40592 17876
rect 40644 17864 40650 17876
rect 49142 17864 49148 17876
rect 40644 17836 49148 17864
rect 40644 17824 40650 17836
rect 49142 17824 49148 17836
rect 49200 17824 49206 17876
rect 33962 17796 33968 17808
rect 32968 17768 33968 17796
rect 32968 17737 32996 17768
rect 33962 17756 33968 17768
rect 34020 17796 34026 17808
rect 34057 17799 34115 17805
rect 34057 17796 34069 17799
rect 34020 17768 34069 17796
rect 34020 17756 34026 17768
rect 34057 17765 34069 17768
rect 34103 17796 34115 17799
rect 34238 17796 34244 17808
rect 34103 17768 34244 17796
rect 34103 17765 34115 17768
rect 34057 17759 34115 17765
rect 34238 17756 34244 17768
rect 34296 17756 34302 17808
rect 34333 17799 34391 17805
rect 34333 17765 34345 17799
rect 34379 17796 34391 17799
rect 34974 17796 34980 17808
rect 34379 17768 34980 17796
rect 34379 17765 34391 17768
rect 34333 17759 34391 17765
rect 34974 17756 34980 17768
rect 35032 17756 35038 17808
rect 38749 17799 38807 17805
rect 38749 17765 38761 17799
rect 38795 17796 38807 17799
rect 40862 17796 40868 17808
rect 38795 17768 40868 17796
rect 38795 17765 38807 17768
rect 38749 17759 38807 17765
rect 40862 17756 40868 17768
rect 40920 17756 40926 17808
rect 31573 17731 31631 17737
rect 31573 17697 31585 17731
rect 31619 17697 31631 17731
rect 31573 17691 31631 17697
rect 32953 17731 33011 17737
rect 32953 17697 32965 17731
rect 32999 17697 33011 17731
rect 32953 17691 33011 17697
rect 33045 17731 33103 17737
rect 33045 17697 33057 17731
rect 33091 17728 33103 17731
rect 33226 17728 33232 17740
rect 33091 17700 33232 17728
rect 33091 17697 33103 17700
rect 33045 17691 33103 17697
rect 33226 17688 33232 17700
rect 33284 17688 33290 17740
rect 34514 17688 34520 17740
rect 34572 17728 34578 17740
rect 35710 17728 35716 17740
rect 34572 17700 35716 17728
rect 34572 17688 34578 17700
rect 35710 17688 35716 17700
rect 35768 17728 35774 17740
rect 35805 17731 35863 17737
rect 35805 17728 35817 17731
rect 35768 17700 35817 17728
rect 35768 17688 35774 17700
rect 35805 17697 35817 17700
rect 35851 17697 35863 17731
rect 35805 17691 35863 17697
rect 37274 17688 37280 17740
rect 37332 17728 37338 17740
rect 38105 17731 38163 17737
rect 38105 17728 38117 17731
rect 37332 17700 38117 17728
rect 37332 17688 37338 17700
rect 38105 17697 38117 17700
rect 38151 17697 38163 17731
rect 39209 17731 39267 17737
rect 39209 17728 39221 17731
rect 38105 17691 38163 17697
rect 38672 17700 39221 17728
rect 38672 17672 38700 17700
rect 39209 17697 39221 17700
rect 39255 17728 39267 17731
rect 40034 17728 40040 17740
rect 39255 17700 40040 17728
rect 39255 17697 39267 17700
rect 39209 17691 39267 17697
rect 40034 17688 40040 17700
rect 40092 17688 40098 17740
rect 40678 17688 40684 17740
rect 40736 17728 40742 17740
rect 40957 17731 41015 17737
rect 40957 17728 40969 17731
rect 40736 17700 40969 17728
rect 40736 17688 40742 17700
rect 40957 17697 40969 17700
rect 41003 17697 41015 17731
rect 40957 17691 41015 17697
rect 41049 17731 41107 17737
rect 41049 17697 41061 17731
rect 41095 17697 41107 17731
rect 41049 17691 41107 17697
rect 23532 17632 25176 17660
rect 25961 17663 26019 17669
rect 23532 17620 23538 17632
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 27430 17620 27436 17672
rect 27488 17620 27494 17672
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17660 28871 17663
rect 28902 17660 28908 17672
rect 28859 17632 28908 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 28902 17620 28908 17632
rect 28960 17660 28966 17672
rect 31665 17663 31723 17669
rect 28960 17632 30788 17660
rect 28960 17620 28966 17632
rect 30760 17604 30788 17632
rect 31665 17629 31677 17663
rect 31711 17660 31723 17663
rect 31754 17660 31760 17672
rect 31711 17632 31760 17660
rect 31711 17629 31723 17632
rect 31665 17623 31723 17629
rect 31754 17620 31760 17632
rect 31812 17620 31818 17672
rect 34425 17663 34483 17669
rect 34425 17660 34437 17663
rect 33428 17632 34437 17660
rect 20990 17552 20996 17604
rect 21048 17552 21054 17604
rect 21726 17552 21732 17604
rect 21784 17592 21790 17604
rect 22281 17595 22339 17601
rect 22281 17592 22293 17595
rect 21784 17564 22293 17592
rect 21784 17552 21790 17564
rect 22281 17561 22293 17564
rect 22327 17561 22339 17595
rect 22281 17555 22339 17561
rect 22833 17595 22891 17601
rect 22833 17561 22845 17595
rect 22879 17592 22891 17595
rect 23661 17595 23719 17601
rect 23661 17592 23673 17595
rect 22879 17564 23673 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 23661 17561 23673 17564
rect 23707 17561 23719 17595
rect 23661 17555 23719 17561
rect 24762 17552 24768 17604
rect 24820 17592 24826 17604
rect 26421 17595 26479 17601
rect 26421 17592 26433 17595
rect 24820 17564 26433 17592
rect 24820 17552 24826 17564
rect 26421 17561 26433 17564
rect 26467 17592 26479 17595
rect 27246 17592 27252 17604
rect 26467 17564 27252 17592
rect 26467 17561 26479 17564
rect 26421 17555 26479 17561
rect 27246 17552 27252 17564
rect 27304 17552 27310 17604
rect 29365 17595 29423 17601
rect 29365 17592 29377 17595
rect 28966 17564 29377 17592
rect 22094 17524 22100 17536
rect 20456 17496 22100 17524
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 23750 17484 23756 17536
rect 23808 17484 23814 17536
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24912 17496 24961 17524
rect 24912 17484 24918 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 27065 17527 27123 17533
rect 27065 17493 27077 17527
rect 27111 17524 27123 17527
rect 27614 17524 27620 17536
rect 27111 17496 27620 17524
rect 27111 17493 27123 17496
rect 27065 17487 27123 17493
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 28810 17484 28816 17536
rect 28868 17524 28874 17536
rect 28966 17524 28994 17564
rect 29365 17561 29377 17564
rect 29411 17592 29423 17595
rect 29917 17595 29975 17601
rect 29917 17592 29929 17595
rect 29411 17564 29929 17592
rect 29411 17561 29423 17564
rect 29365 17555 29423 17561
rect 29917 17561 29929 17564
rect 29963 17592 29975 17595
rect 30006 17592 30012 17604
rect 29963 17564 30012 17592
rect 29963 17561 29975 17564
rect 29917 17555 29975 17561
rect 30006 17552 30012 17564
rect 30064 17552 30070 17604
rect 30742 17552 30748 17604
rect 30800 17552 30806 17604
rect 33428 17536 33456 17632
rect 34425 17629 34437 17632
rect 34471 17629 34483 17663
rect 34425 17623 34483 17629
rect 37550 17620 37556 17672
rect 37608 17620 37614 17672
rect 37918 17620 37924 17672
rect 37976 17660 37982 17672
rect 38654 17660 38660 17672
rect 37976 17632 38660 17660
rect 37976 17620 37982 17632
rect 38654 17620 38660 17632
rect 38712 17620 38718 17672
rect 38838 17620 38844 17672
rect 38896 17660 38902 17672
rect 41064 17660 41092 17691
rect 38896 17632 41092 17660
rect 48593 17663 48651 17669
rect 38896 17620 38902 17632
rect 48593 17629 48605 17663
rect 48639 17660 48651 17663
rect 49326 17660 49332 17672
rect 48639 17632 49332 17660
rect 48639 17629 48651 17632
rect 48593 17623 48651 17629
rect 49326 17620 49332 17632
rect 49384 17620 49390 17672
rect 35986 17592 35992 17604
rect 33520 17564 35992 17592
rect 28868 17496 28994 17524
rect 28868 17484 28874 17496
rect 31938 17484 31944 17536
rect 31996 17524 32002 17536
rect 32033 17527 32091 17533
rect 32033 17524 32045 17527
rect 31996 17496 32045 17524
rect 31996 17484 32002 17496
rect 32033 17493 32045 17496
rect 32079 17493 32091 17527
rect 32033 17487 32091 17493
rect 32306 17484 32312 17536
rect 32364 17484 32370 17536
rect 33137 17527 33195 17533
rect 33137 17493 33149 17527
rect 33183 17524 33195 17527
rect 33410 17524 33416 17536
rect 33183 17496 33416 17524
rect 33183 17493 33195 17496
rect 33137 17487 33195 17493
rect 33410 17484 33416 17496
rect 33468 17484 33474 17536
rect 33520 17533 33548 17564
rect 35986 17552 35992 17564
rect 36044 17552 36050 17604
rect 36538 17552 36544 17604
rect 36596 17552 36602 17604
rect 36998 17552 37004 17604
rect 37056 17592 37062 17604
rect 37277 17595 37335 17601
rect 37277 17592 37289 17595
rect 37056 17564 37289 17592
rect 37056 17552 37062 17564
rect 37277 17561 37289 17564
rect 37323 17561 37335 17595
rect 37277 17555 37335 17561
rect 37366 17552 37372 17604
rect 37424 17592 37430 17604
rect 38381 17595 38439 17601
rect 38381 17592 38393 17595
rect 37424 17564 38393 17592
rect 37424 17552 37430 17564
rect 38381 17561 38393 17564
rect 38427 17561 38439 17595
rect 38381 17555 38439 17561
rect 40865 17595 40923 17601
rect 40865 17561 40877 17595
rect 40911 17592 40923 17595
rect 48406 17592 48412 17604
rect 40911 17564 48412 17592
rect 40911 17561 40923 17564
rect 40865 17555 40923 17561
rect 48406 17552 48412 17564
rect 48464 17552 48470 17604
rect 48777 17595 48835 17601
rect 48777 17561 48789 17595
rect 48823 17592 48835 17595
rect 49234 17592 49240 17604
rect 48823 17564 49240 17592
rect 48823 17561 48835 17564
rect 48777 17555 48835 17561
rect 49234 17552 49240 17564
rect 49292 17552 49298 17604
rect 33505 17527 33563 17533
rect 33505 17493 33517 17527
rect 33551 17493 33563 17527
rect 33505 17487 33563 17493
rect 35066 17484 35072 17536
rect 35124 17484 35130 17536
rect 35437 17527 35495 17533
rect 35437 17493 35449 17527
rect 35483 17524 35495 17527
rect 35526 17524 35532 17536
rect 35483 17496 35532 17524
rect 35483 17493 35495 17496
rect 35437 17487 35495 17493
rect 35526 17484 35532 17496
rect 35584 17484 35590 17536
rect 36630 17484 36636 17536
rect 36688 17524 36694 17536
rect 38289 17527 38347 17533
rect 38289 17524 38301 17527
rect 36688 17496 38301 17524
rect 36688 17484 36694 17496
rect 38289 17493 38301 17496
rect 38335 17493 38347 17527
rect 38289 17487 38347 17493
rect 38930 17484 38936 17536
rect 38988 17524 38994 17536
rect 39025 17527 39083 17533
rect 39025 17524 39037 17527
rect 38988 17496 39037 17524
rect 38988 17484 38994 17496
rect 39025 17493 39037 17496
rect 39071 17493 39083 17527
rect 39025 17487 39083 17493
rect 49142 17484 49148 17536
rect 49200 17484 49206 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 11793 17323 11851 17329
rect 11793 17320 11805 17323
rect 7892 17292 11805 17320
rect 7892 17280 7898 17292
rect 11793 17289 11805 17292
rect 11839 17289 11851 17323
rect 11793 17283 11851 17289
rect 13081 17323 13139 17329
rect 13081 17289 13093 17323
rect 13127 17320 13139 17323
rect 13354 17320 13360 17332
rect 13127 17292 13360 17320
rect 13127 17289 13139 17292
rect 13081 17283 13139 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14056 17292 14933 17320
rect 14056 17280 14062 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 15562 17280 15568 17332
rect 15620 17280 15626 17332
rect 15672 17292 18092 17320
rect 3326 17212 3332 17264
rect 3384 17252 3390 17264
rect 3384 17224 10916 17252
rect 3384 17212 3390 17224
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 4338 17184 4344 17196
rect 3007 17156 4344 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 9490 17144 9496 17196
rect 9548 17184 9554 17196
rect 10502 17184 10508 17196
rect 9548 17156 10508 17184
rect 9548 17144 9554 17156
rect 10502 17144 10508 17156
rect 10560 17184 10566 17196
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10560 17156 10701 17184
rect 10560 17144 10566 17156
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 10778 17144 10784 17196
rect 10836 17144 10842 17196
rect 10888 17184 10916 17224
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11882 17252 11888 17264
rect 11480 17224 11888 17252
rect 11480 17212 11486 17224
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 12989 17255 13047 17261
rect 12989 17252 13001 17255
rect 12216 17224 13001 17252
rect 12216 17212 12222 17224
rect 12989 17221 13001 17224
rect 13035 17221 13047 17255
rect 12989 17215 13047 17221
rect 13906 17212 13912 17264
rect 13964 17252 13970 17264
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 13964 17224 14289 17252
rect 13964 17212 13970 17224
rect 14277 17221 14289 17224
rect 14323 17221 14335 17255
rect 14277 17215 14335 17221
rect 14734 17212 14740 17264
rect 14792 17252 14798 17264
rect 15672 17252 15700 17292
rect 14792 17224 15700 17252
rect 14792 17212 14798 17224
rect 15746 17212 15752 17264
rect 15804 17252 15810 17264
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15804 17224 15945 17252
rect 15804 17212 15810 17224
rect 15933 17221 15945 17224
rect 15979 17221 15991 17255
rect 15933 17215 15991 17221
rect 16022 17212 16028 17264
rect 16080 17252 16086 17264
rect 17954 17252 17960 17264
rect 16080 17224 17960 17252
rect 16080 17212 16086 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 18064 17252 18092 17292
rect 19150 17280 19156 17332
rect 19208 17280 19214 17332
rect 19702 17320 19708 17332
rect 19260 17292 19708 17320
rect 19260 17252 19288 17292
rect 19702 17280 19708 17292
rect 19760 17280 19766 17332
rect 20898 17320 20904 17332
rect 20548 17292 20904 17320
rect 20548 17252 20576 17292
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 22649 17323 22707 17329
rect 22649 17289 22661 17323
rect 22695 17320 22707 17323
rect 23474 17320 23480 17332
rect 22695 17292 23480 17320
rect 22695 17289 22707 17292
rect 22649 17283 22707 17289
rect 23474 17280 23480 17292
rect 23532 17280 23538 17332
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 24946 17320 24952 17332
rect 24903 17292 24952 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 24946 17280 24952 17292
rect 25004 17280 25010 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 27341 17323 27399 17329
rect 27341 17320 27353 17323
rect 25363 17292 27353 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 27341 17289 27353 17292
rect 27387 17289 27399 17323
rect 27341 17283 27399 17289
rect 27706 17280 27712 17332
rect 27764 17280 27770 17332
rect 27798 17280 27804 17332
rect 27856 17320 27862 17332
rect 28997 17323 29055 17329
rect 28997 17320 29009 17323
rect 27856 17292 29009 17320
rect 27856 17280 27862 17292
rect 28997 17289 29009 17292
rect 29043 17289 29055 17323
rect 28997 17283 29055 17289
rect 29270 17280 29276 17332
rect 29328 17320 29334 17332
rect 30101 17323 30159 17329
rect 30101 17320 30113 17323
rect 29328 17292 30113 17320
rect 29328 17280 29334 17292
rect 30101 17289 30113 17292
rect 30147 17289 30159 17323
rect 30101 17283 30159 17289
rect 30561 17323 30619 17329
rect 30561 17289 30573 17323
rect 30607 17289 30619 17323
rect 30561 17283 30619 17289
rect 18064 17224 19288 17252
rect 20194 17224 20576 17252
rect 20625 17255 20683 17261
rect 20625 17221 20637 17255
rect 20671 17252 20683 17255
rect 20990 17252 20996 17264
rect 20671 17224 20996 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 20990 17212 20996 17224
rect 21048 17252 21054 17264
rect 21450 17252 21456 17264
rect 21048 17224 21456 17252
rect 21048 17212 21054 17224
rect 21450 17212 21456 17224
rect 21508 17212 21514 17264
rect 21542 17212 21548 17264
rect 21600 17252 21606 17264
rect 22097 17255 22155 17261
rect 22097 17252 22109 17255
rect 21600 17224 22109 17252
rect 21600 17212 21606 17224
rect 22097 17221 22109 17224
rect 22143 17252 22155 17255
rect 22830 17252 22836 17264
rect 22143 17224 22836 17252
rect 22143 17221 22155 17224
rect 22097 17215 22155 17221
rect 22830 17212 22836 17224
rect 22888 17252 22894 17264
rect 22888 17224 22954 17252
rect 22888 17212 22894 17224
rect 24118 17212 24124 17264
rect 24176 17252 24182 17264
rect 24176 17224 24440 17252
rect 24176 17212 24182 17224
rect 10888 17156 13032 17184
rect 934 17076 940 17128
rect 992 17116 998 17128
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 992 17088 1777 17116
rect 992 17076 998 17088
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 5868 17088 9873 17116
rect 5868 17076 5874 17088
rect 9490 16940 9496 16992
rect 9548 16940 9554 16992
rect 9692 16980 9720 17088
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17085 10655 17119
rect 12802 17116 12808 17128
rect 10597 17079 10655 17085
rect 10796 17088 12808 17116
rect 9769 17051 9827 17057
rect 9769 17017 9781 17051
rect 9815 17048 9827 17051
rect 10137 17051 10195 17057
rect 10137 17048 10149 17051
rect 9815 17020 10149 17048
rect 9815 17017 9827 17020
rect 9769 17011 9827 17017
rect 10137 17017 10149 17020
rect 10183 17048 10195 17051
rect 10612 17048 10640 17079
rect 10796 17048 10824 17088
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 13004 17116 13032 17156
rect 15102 17144 15108 17196
rect 15160 17144 15166 17196
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 15764 17184 15792 17212
rect 16942 17184 16948 17196
rect 15252 17156 15792 17184
rect 15948 17156 16948 17184
rect 15252 17144 15258 17156
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13004 17088 14105 17116
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 14642 17076 14648 17128
rect 14700 17116 14706 17128
rect 15948 17116 15976 17156
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 18693 17187 18751 17193
rect 18693 17153 18705 17187
rect 18739 17184 18751 17187
rect 18874 17184 18880 17196
rect 18739 17156 18880 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 14700 17088 15976 17116
rect 16025 17119 16083 17125
rect 14700 17076 14706 17088
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 10183 17020 10824 17048
rect 11149 17051 11207 17057
rect 10183 17017 10195 17020
rect 10137 17011 10195 17017
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 12618 17048 12624 17060
rect 11195 17020 12624 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 16040 17048 16068 17079
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 17052 17116 17080 17147
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 22186 17184 22192 17196
rect 20947 17156 22192 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 22186 17144 22192 17156
rect 22244 17184 22250 17196
rect 22738 17184 22744 17196
rect 22244 17156 22744 17184
rect 22244 17144 22250 17156
rect 22738 17144 22744 17156
rect 22796 17144 22802 17196
rect 24412 17193 24440 17224
rect 25958 17212 25964 17264
rect 26016 17212 26022 17264
rect 28905 17255 28963 17261
rect 28905 17221 28917 17255
rect 28951 17252 28963 17255
rect 29638 17252 29644 17264
rect 28951 17224 29644 17252
rect 28951 17221 28963 17224
rect 28905 17215 28963 17221
rect 29638 17212 29644 17224
rect 29696 17212 29702 17264
rect 30576 17252 30604 17283
rect 30926 17280 30932 17332
rect 30984 17320 30990 17332
rect 31297 17323 31355 17329
rect 31297 17320 31309 17323
rect 30984 17292 31309 17320
rect 30984 17280 30990 17292
rect 31297 17289 31309 17292
rect 31343 17289 31355 17323
rect 31297 17283 31355 17289
rect 31389 17323 31447 17329
rect 31389 17289 31401 17323
rect 31435 17320 31447 17323
rect 31570 17320 31576 17332
rect 31435 17292 31576 17320
rect 31435 17289 31447 17292
rect 31389 17283 31447 17289
rect 31570 17280 31576 17292
rect 31628 17280 31634 17332
rect 33594 17320 33600 17332
rect 32324 17292 33600 17320
rect 30650 17252 30656 17264
rect 30576 17224 30656 17252
rect 30650 17212 30656 17224
rect 30708 17212 30714 17264
rect 30742 17212 30748 17264
rect 30800 17252 30806 17264
rect 32324 17252 32352 17292
rect 33594 17280 33600 17292
rect 33652 17280 33658 17332
rect 34054 17280 34060 17332
rect 34112 17280 34118 17332
rect 35066 17280 35072 17332
rect 35124 17320 35130 17332
rect 37829 17323 37887 17329
rect 37829 17320 37841 17323
rect 35124 17292 37841 17320
rect 35124 17280 35130 17292
rect 37829 17289 37841 17292
rect 37875 17289 37887 17323
rect 40586 17320 40592 17332
rect 37829 17283 37887 17289
rect 37936 17292 40592 17320
rect 33870 17252 33876 17264
rect 30800 17224 32352 17252
rect 33810 17224 33876 17252
rect 30800 17212 30806 17224
rect 24397 17187 24455 17193
rect 24397 17153 24409 17187
rect 24443 17153 24455 17187
rect 24397 17147 24455 17153
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17184 25283 17187
rect 25590 17184 25596 17196
rect 25271 17156 25596 17184
rect 25271 17153 25283 17156
rect 25225 17147 25283 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 26418 17184 26424 17196
rect 25700 17156 26424 17184
rect 19886 17116 19892 17128
rect 17052 17088 19892 17116
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 19978 17076 19984 17128
rect 20036 17116 20042 17128
rect 21818 17116 21824 17128
rect 20036 17088 21824 17116
rect 20036 17076 20042 17088
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 22002 17076 22008 17128
rect 22060 17076 22066 17128
rect 24121 17119 24179 17125
rect 24121 17085 24133 17119
rect 24167 17116 24179 17119
rect 24167 17088 24624 17116
rect 24167 17085 24179 17088
rect 24121 17079 24179 17085
rect 24596 17060 24624 17088
rect 25498 17076 25504 17128
rect 25556 17076 25562 17128
rect 16482 17048 16488 17060
rect 16040 17020 16488 17048
rect 16482 17008 16488 17020
rect 16540 17048 16546 17060
rect 16540 17020 17540 17048
rect 16540 17008 16546 17020
rect 12158 16980 12164 16992
rect 9692 16952 12164 16980
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12434 16940 12440 16992
rect 12492 16940 12498 16992
rect 13446 16940 13452 16992
rect 13504 16940 13510 16992
rect 13817 16983 13875 16989
rect 13817 16949 13829 16983
rect 13863 16980 13875 16983
rect 14090 16980 14096 16992
rect 13863 16952 14096 16980
rect 13863 16949 13875 16952
rect 13817 16943 13875 16949
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 16758 16940 16764 16992
rect 16816 16980 16822 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16816 16952 16957 16980
rect 16816 16940 16822 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 17402 16940 17408 16992
rect 17460 16940 17466 16992
rect 17512 16980 17540 17020
rect 20824 17020 22094 17048
rect 20824 16980 20852 17020
rect 17512 16952 20852 16980
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21177 16983 21235 16989
rect 21177 16980 21189 16983
rect 20956 16952 21189 16980
rect 20956 16940 20962 16952
rect 21177 16949 21189 16952
rect 21223 16980 21235 16983
rect 21542 16980 21548 16992
rect 21223 16952 21548 16980
rect 21223 16949 21235 16952
rect 21177 16943 21235 16949
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 22066 16980 22094 17020
rect 24578 17008 24584 17060
rect 24636 17048 24642 17060
rect 25700 17048 25728 17156
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 27062 17144 27068 17196
rect 27120 17184 27126 17196
rect 27120 17156 27936 17184
rect 27120 17144 27126 17156
rect 27798 17116 27804 17128
rect 24636 17020 25728 17048
rect 25792 17088 27804 17116
rect 24636 17008 24642 17020
rect 25792 16980 25820 17088
rect 27798 17076 27804 17088
rect 27856 17076 27862 17128
rect 27908 17125 27936 17156
rect 28258 17144 28264 17196
rect 28316 17184 28322 17196
rect 29178 17184 29184 17196
rect 28316 17156 29184 17184
rect 28316 17144 28322 17156
rect 29178 17144 29184 17156
rect 29236 17144 29242 17196
rect 30193 17187 30251 17193
rect 30193 17153 30205 17187
rect 30239 17184 30251 17187
rect 30239 17156 31432 17184
rect 30239 17153 30251 17156
rect 30193 17147 30251 17153
rect 27893 17119 27951 17125
rect 27893 17085 27905 17119
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 28721 17119 28779 17125
rect 28721 17085 28733 17119
rect 28767 17085 28779 17119
rect 28721 17079 28779 17085
rect 26878 17008 26884 17060
rect 26936 17048 26942 17060
rect 28736 17048 28764 17079
rect 29914 17076 29920 17128
rect 29972 17076 29978 17128
rect 30742 17076 30748 17128
rect 30800 17116 30806 17128
rect 31113 17119 31171 17125
rect 31113 17116 31125 17119
rect 30800 17088 31125 17116
rect 30800 17076 30806 17088
rect 31113 17085 31125 17088
rect 31159 17085 31171 17119
rect 31404 17116 31432 17156
rect 32214 17144 32220 17196
rect 32272 17184 32278 17196
rect 32324 17193 32352 17224
rect 33870 17212 33876 17224
rect 33928 17252 33934 17264
rect 34974 17252 34980 17264
rect 33928 17224 34980 17252
rect 33928 17212 33934 17224
rect 34974 17212 34980 17224
rect 35032 17212 35038 17264
rect 35526 17212 35532 17264
rect 35584 17252 35590 17264
rect 37001 17255 37059 17261
rect 37001 17252 37013 17255
rect 35584 17224 37013 17252
rect 35584 17212 35590 17224
rect 37001 17221 37013 17224
rect 37047 17221 37059 17255
rect 37936 17252 37964 17292
rect 40586 17280 40592 17292
rect 40644 17280 40650 17332
rect 48406 17280 48412 17332
rect 48464 17280 48470 17332
rect 37001 17215 37059 17221
rect 37108 17224 37964 17252
rect 38565 17255 38623 17261
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 32272 17156 32321 17184
rect 32272 17144 32278 17156
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 35618 17144 35624 17196
rect 35676 17184 35682 17196
rect 36265 17187 36323 17193
rect 36265 17184 36277 17187
rect 35676 17156 36277 17184
rect 35676 17144 35682 17156
rect 36265 17153 36277 17156
rect 36311 17153 36323 17187
rect 36265 17147 36323 17153
rect 36354 17144 36360 17196
rect 36412 17144 36418 17196
rect 31404 17088 32352 17116
rect 31113 17079 31171 17085
rect 32324 17060 32352 17088
rect 32582 17076 32588 17128
rect 32640 17076 32646 17128
rect 34790 17076 34796 17128
rect 34848 17076 34854 17128
rect 36170 17076 36176 17128
rect 36228 17076 36234 17128
rect 37108 17116 37136 17224
rect 38565 17221 38577 17255
rect 38611 17252 38623 17255
rect 38654 17252 38660 17264
rect 38611 17224 38660 17252
rect 38611 17221 38623 17224
rect 38565 17215 38623 17221
rect 38654 17212 38660 17224
rect 38712 17252 38718 17264
rect 38712 17224 39238 17252
rect 38712 17212 38718 17224
rect 40126 17212 40132 17264
rect 40184 17252 40190 17264
rect 40405 17255 40463 17261
rect 40405 17252 40417 17255
rect 40184 17224 40417 17252
rect 40184 17212 40190 17224
rect 40405 17221 40417 17224
rect 40451 17221 40463 17255
rect 40405 17215 40463 17221
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17184 37979 17187
rect 38930 17184 38936 17196
rect 37967 17156 38936 17184
rect 37967 17153 37979 17156
rect 37921 17147 37979 17153
rect 38930 17144 38936 17156
rect 38988 17144 38994 17196
rect 48593 17187 48651 17193
rect 48593 17153 48605 17187
rect 48639 17184 48651 17187
rect 48774 17184 48780 17196
rect 48639 17156 48780 17184
rect 48639 17153 48651 17156
rect 48593 17147 48651 17153
rect 48774 17144 48780 17156
rect 48832 17144 48838 17196
rect 49237 17187 49295 17193
rect 49237 17153 49249 17187
rect 49283 17184 49295 17187
rect 49326 17184 49332 17196
rect 49283 17156 49332 17184
rect 49283 17153 49295 17156
rect 49237 17147 49295 17153
rect 49326 17144 49332 17156
rect 49384 17144 49390 17196
rect 36280 17088 37136 17116
rect 26936 17020 28764 17048
rect 29365 17051 29423 17057
rect 26936 17008 26942 17020
rect 29365 17017 29377 17051
rect 29411 17048 29423 17051
rect 32122 17048 32128 17060
rect 29411 17020 32128 17048
rect 29411 17017 29423 17020
rect 29365 17011 29423 17017
rect 32122 17008 32128 17020
rect 32180 17008 32186 17060
rect 32306 17008 32312 17060
rect 32364 17008 32370 17060
rect 35434 17008 35440 17060
rect 35492 17048 35498 17060
rect 36280 17048 36308 17088
rect 37826 17076 37832 17128
rect 37884 17116 37890 17128
rect 38013 17119 38071 17125
rect 38013 17116 38025 17119
rect 37884 17088 38025 17116
rect 37884 17076 37890 17088
rect 38013 17085 38025 17088
rect 38059 17085 38071 17119
rect 38013 17079 38071 17085
rect 38378 17076 38384 17128
rect 38436 17116 38442 17128
rect 38436 17088 40632 17116
rect 38436 17076 38442 17088
rect 35492 17020 36308 17048
rect 35492 17008 35498 17020
rect 36446 17008 36452 17060
rect 36504 17048 36510 17060
rect 37461 17051 37519 17057
rect 37461 17048 37473 17051
rect 36504 17020 37473 17048
rect 36504 17008 36510 17020
rect 37461 17017 37473 17020
rect 37507 17017 37519 17051
rect 40604 17048 40632 17088
rect 40678 17076 40684 17128
rect 40736 17076 40742 17128
rect 49050 17076 49056 17128
rect 49108 17076 49114 17128
rect 43898 17048 43904 17060
rect 40604 17020 43904 17048
rect 37461 17011 37519 17017
rect 43898 17008 43904 17020
rect 43956 17008 43962 17060
rect 22066 16952 25820 16980
rect 26234 16940 26240 16992
rect 26292 16980 26298 16992
rect 27982 16980 27988 16992
rect 26292 16952 27988 16980
rect 26292 16940 26298 16952
rect 27982 16940 27988 16952
rect 28040 16940 28046 16992
rect 28626 16940 28632 16992
rect 28684 16980 28690 16992
rect 31294 16980 31300 16992
rect 28684 16952 31300 16980
rect 28684 16940 28690 16952
rect 31294 16940 31300 16952
rect 31352 16940 31358 16992
rect 31754 16940 31760 16992
rect 31812 16940 31818 16992
rect 31846 16940 31852 16992
rect 31904 16980 31910 16992
rect 35342 16980 35348 16992
rect 31904 16952 35348 16980
rect 31904 16940 31910 16952
rect 35342 16940 35348 16952
rect 35400 16940 35406 16992
rect 36722 16940 36728 16992
rect 36780 16940 36786 16992
rect 38838 16940 38844 16992
rect 38896 16980 38902 16992
rect 38933 16983 38991 16989
rect 38933 16980 38945 16983
rect 38896 16952 38945 16980
rect 38896 16940 38902 16952
rect 38933 16949 38945 16952
rect 38979 16949 38991 16983
rect 38933 16943 38991 16949
rect 40034 16940 40040 16992
rect 40092 16980 40098 16992
rect 40957 16983 41015 16989
rect 40957 16980 40969 16983
rect 40092 16952 40969 16980
rect 40092 16940 40098 16952
rect 40957 16949 40969 16952
rect 41003 16980 41015 16983
rect 41046 16980 41052 16992
rect 41003 16952 41052 16980
rect 41003 16949 41015 16952
rect 40957 16943 41015 16949
rect 41046 16940 41052 16952
rect 41104 16940 41110 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 10410 16736 10416 16788
rect 10468 16736 10474 16788
rect 14826 16776 14832 16788
rect 13280 16748 14832 16776
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 13280 16708 13308 16748
rect 14826 16736 14832 16748
rect 14884 16776 14890 16788
rect 14884 16748 16252 16776
rect 14884 16736 14890 16748
rect 10376 16680 12434 16708
rect 10376 16668 10382 16680
rect 12406 16652 12434 16680
rect 13188 16680 13308 16708
rect 14185 16711 14243 16717
rect 4430 16600 4436 16652
rect 4488 16640 4494 16652
rect 5442 16640 5448 16652
rect 4488 16612 5448 16640
rect 4488 16600 4494 16612
rect 5442 16600 5448 16612
rect 5500 16640 5506 16652
rect 7929 16643 7987 16649
rect 5500 16612 7696 16640
rect 5500 16600 5506 16612
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3326 16572 3332 16584
rect 3007 16544 3332 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 1026 16464 1032 16516
rect 1084 16504 1090 16516
rect 1765 16507 1823 16513
rect 1765 16504 1777 16507
rect 1084 16476 1777 16504
rect 1084 16464 1090 16476
rect 1765 16473 1777 16476
rect 1811 16473 1823 16507
rect 7668 16504 7696 16612
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 9030 16640 9036 16652
rect 7975 16612 9036 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 10962 16600 10968 16652
rect 11020 16640 11026 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11020 16612 11161 16640
rect 11020 16600 11026 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 12406 16612 12440 16652
rect 11149 16603 11207 16609
rect 12434 16600 12440 16612
rect 12492 16640 12498 16652
rect 13188 16649 13216 16680
rect 14185 16677 14197 16711
rect 14231 16708 14243 16711
rect 14274 16708 14280 16720
rect 14231 16680 14280 16708
rect 14231 16677 14243 16680
rect 14185 16671 14243 16677
rect 14274 16668 14280 16680
rect 14332 16668 14338 16720
rect 15562 16708 15568 16720
rect 14568 16680 15568 16708
rect 13173 16643 13231 16649
rect 12492 16612 13124 16640
rect 12492 16600 12498 16612
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 7800 16544 8125 16572
rect 7800 16532 7806 16544
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12308 16544 12357 16572
rect 12308 16532 12314 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 13096 16572 13124 16612
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13311 16612 14044 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13280 16572 13308 16603
rect 13096 16544 13308 16572
rect 13357 16575 13415 16581
rect 12345 16535 12403 16541
rect 13357 16541 13369 16575
rect 13403 16572 13415 16575
rect 13814 16572 13820 16584
rect 13403 16544 13820 16572
rect 13403 16541 13415 16544
rect 13357 16535 13415 16541
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 8021 16507 8079 16513
rect 8021 16504 8033 16507
rect 7668 16476 8033 16504
rect 1765 16467 1823 16473
rect 8021 16473 8033 16476
rect 8067 16473 8079 16507
rect 9674 16504 9680 16516
rect 8021 16467 8079 16473
rect 8496 16476 9680 16504
rect 8496 16445 8524 16476
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 10045 16507 10103 16513
rect 10045 16473 10057 16507
rect 10091 16504 10103 16507
rect 10502 16504 10508 16516
rect 10091 16476 10508 16504
rect 10091 16473 10103 16476
rect 10045 16467 10103 16473
rect 10502 16464 10508 16476
rect 10560 16464 10566 16516
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 12802 16504 12808 16516
rect 11471 16476 12808 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 8481 16439 8539 16445
rect 8481 16405 8493 16439
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 9030 16396 9036 16448
rect 9088 16396 9094 16448
rect 11330 16396 11336 16448
rect 11388 16396 11394 16448
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16436 11851 16439
rect 12434 16436 12440 16448
rect 11839 16408 12440 16436
rect 11839 16405 11851 16408
rect 11793 16399 11851 16405
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 12529 16439 12587 16445
rect 12529 16405 12541 16439
rect 12575 16436 12587 16439
rect 12710 16436 12716 16448
rect 12575 16408 12716 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 13262 16396 13268 16448
rect 13320 16436 13326 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 13320 16408 13737 16436
rect 13320 16396 13326 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13832 16436 13860 16532
rect 14016 16504 14044 16612
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 14568 16649 14596 16680
rect 15562 16668 15568 16680
rect 15620 16668 15626 16720
rect 16224 16649 16252 16748
rect 17402 16736 17408 16788
rect 17460 16776 17466 16788
rect 17460 16748 18828 16776
rect 17460 16736 17466 16748
rect 18800 16708 18828 16748
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 20990 16776 20996 16788
rect 20772 16748 20996 16776
rect 20772 16736 20778 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21726 16776 21732 16788
rect 21100 16748 21732 16776
rect 21100 16708 21128 16748
rect 21726 16736 21732 16748
rect 21784 16736 21790 16788
rect 21818 16736 21824 16788
rect 21876 16776 21882 16788
rect 21876 16748 23244 16776
rect 21876 16736 21882 16748
rect 18800 16680 21128 16708
rect 23216 16708 23244 16748
rect 23290 16736 23296 16788
rect 23348 16776 23354 16788
rect 24765 16779 24823 16785
rect 24765 16776 24777 16779
rect 23348 16748 24777 16776
rect 23348 16736 23354 16748
rect 24765 16745 24777 16748
rect 24811 16776 24823 16779
rect 28810 16776 28816 16788
rect 24811 16748 28816 16776
rect 24811 16745 24823 16748
rect 24765 16739 24823 16745
rect 28810 16736 28816 16748
rect 28868 16736 28874 16788
rect 29181 16779 29239 16785
rect 29181 16745 29193 16779
rect 29227 16776 29239 16779
rect 30098 16776 30104 16788
rect 29227 16748 30104 16776
rect 29227 16745 29239 16748
rect 29181 16739 29239 16745
rect 30098 16736 30104 16748
rect 30156 16736 30162 16788
rect 34514 16776 34520 16788
rect 31128 16748 34520 16776
rect 26050 16708 26056 16720
rect 23216 16680 23704 16708
rect 14553 16643 14611 16649
rect 14148 16612 14504 16640
rect 14148 16600 14154 16612
rect 14476 16572 14504 16612
rect 14553 16609 14565 16643
rect 14599 16609 14611 16643
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 14553 16603 14611 16609
rect 14660 16612 16129 16640
rect 14660 16572 14688 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16609 16267 16643
rect 16850 16640 16856 16652
rect 16209 16603 16267 16609
rect 16316 16612 16856 16640
rect 14476 16544 14688 16572
rect 14734 16532 14740 16584
rect 14792 16532 14798 16584
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16025 16575 16083 16581
rect 16025 16572 16037 16575
rect 15896 16544 16037 16572
rect 15896 16532 15902 16544
rect 16025 16541 16037 16544
rect 16071 16541 16083 16575
rect 16132 16572 16160 16603
rect 16316 16572 16344 16612
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 17954 16600 17960 16652
rect 18012 16640 18018 16652
rect 18877 16643 18935 16649
rect 18877 16640 18889 16643
rect 18012 16612 18889 16640
rect 18012 16600 18018 16612
rect 18877 16609 18889 16612
rect 18923 16640 18935 16643
rect 19150 16640 19156 16652
rect 18923 16612 19156 16640
rect 18923 16609 18935 16612
rect 18877 16603 18935 16609
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 22462 16600 22468 16652
rect 22520 16600 22526 16652
rect 22738 16600 22744 16652
rect 22796 16600 22802 16652
rect 16132 16544 16344 16572
rect 16025 16535 16083 16541
rect 14752 16504 14780 16532
rect 14016 16476 14780 16504
rect 16040 16504 16068 16535
rect 17494 16532 17500 16584
rect 17552 16532 17558 16584
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 16669 16507 16727 16513
rect 16669 16504 16681 16507
rect 16040 16476 16681 16504
rect 16669 16473 16681 16476
rect 16715 16473 16727 16507
rect 16669 16467 16727 16473
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 17000 16476 17356 16504
rect 17000 16464 17006 16476
rect 14182 16436 14188 16448
rect 13832 16408 14188 16436
rect 13725 16399 13783 16405
rect 14182 16396 14188 16408
rect 14240 16436 14246 16448
rect 14829 16439 14887 16445
rect 14829 16436 14841 16439
rect 14240 16408 14841 16436
rect 14240 16396 14246 16408
rect 14829 16405 14841 16408
rect 14875 16405 14887 16439
rect 14829 16399 14887 16405
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16436 15255 16439
rect 15470 16436 15476 16448
rect 15243 16408 15476 16436
rect 15243 16405 15255 16408
rect 15197 16399 15255 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15654 16396 15660 16448
rect 15712 16396 15718 16448
rect 17126 16396 17132 16448
rect 17184 16396 17190 16448
rect 17328 16436 17356 16476
rect 18598 16464 18604 16516
rect 18656 16464 18662 16516
rect 20272 16504 20300 16535
rect 20898 16532 20904 16584
rect 20956 16572 20962 16584
rect 23676 16572 23704 16680
rect 23768 16680 26056 16708
rect 23768 16649 23796 16680
rect 26050 16668 26056 16680
rect 26108 16668 26114 16720
rect 27338 16668 27344 16720
rect 27396 16708 27402 16720
rect 27396 16680 27752 16708
rect 27396 16668 27402 16680
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23937 16643 23995 16649
rect 23937 16609 23949 16643
rect 23983 16640 23995 16643
rect 23983 16612 25544 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 25222 16572 25228 16584
rect 20956 16544 21390 16572
rect 23676 16544 25228 16572
rect 20956 16532 20962 16544
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 18708 16476 20116 16504
rect 20272 16476 21220 16504
rect 18708 16436 18736 16476
rect 17328 16408 18736 16436
rect 19058 16396 19064 16448
rect 19116 16436 19122 16448
rect 20088 16445 20116 16476
rect 19429 16439 19487 16445
rect 19429 16436 19441 16439
rect 19116 16408 19441 16436
rect 19116 16396 19122 16408
rect 19429 16405 19441 16408
rect 19475 16405 19487 16439
rect 19429 16399 19487 16405
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16405 20131 16439
rect 20073 16399 20131 16405
rect 20625 16439 20683 16445
rect 20625 16405 20637 16439
rect 20671 16436 20683 16439
rect 20898 16436 20904 16448
rect 20671 16408 20904 16436
rect 20671 16405 20683 16408
rect 20625 16399 20683 16405
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 21192 16436 21220 16476
rect 22554 16464 22560 16516
rect 22612 16504 22618 16516
rect 24581 16507 24639 16513
rect 22612 16476 23796 16504
rect 22612 16464 22618 16476
rect 22830 16436 22836 16448
rect 21192 16408 22836 16436
rect 22830 16396 22836 16408
rect 22888 16396 22894 16448
rect 23290 16396 23296 16448
rect 23348 16396 23354 16448
rect 23658 16396 23664 16448
rect 23716 16396 23722 16448
rect 23768 16436 23796 16476
rect 24581 16473 24593 16507
rect 24627 16504 24639 16507
rect 24946 16504 24952 16516
rect 24627 16476 24952 16504
rect 24627 16473 24639 16476
rect 24581 16467 24639 16473
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 25314 16436 25320 16448
rect 23768 16408 25320 16436
rect 25314 16396 25320 16408
rect 25372 16396 25378 16448
rect 25516 16436 25544 16612
rect 25682 16600 25688 16652
rect 25740 16640 25746 16652
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 25740 16612 27077 16640
rect 25740 16600 25746 16612
rect 27065 16609 27077 16612
rect 27111 16640 27123 16643
rect 27614 16640 27620 16652
rect 27111 16612 27620 16640
rect 27111 16609 27123 16612
rect 27065 16603 27123 16609
rect 27614 16600 27620 16612
rect 27672 16600 27678 16652
rect 27724 16640 27752 16680
rect 27798 16668 27804 16720
rect 27856 16708 27862 16720
rect 28721 16711 28779 16717
rect 28721 16708 28733 16711
rect 27856 16680 28733 16708
rect 27856 16668 27862 16680
rect 28721 16677 28733 16680
rect 28767 16708 28779 16711
rect 31018 16708 31024 16720
rect 28767 16680 31024 16708
rect 28767 16677 28779 16680
rect 28721 16671 28779 16677
rect 31018 16668 31024 16680
rect 31076 16668 31082 16720
rect 27985 16643 28043 16649
rect 27985 16640 27997 16643
rect 27724 16612 27997 16640
rect 27985 16609 27997 16612
rect 28031 16640 28043 16643
rect 28074 16640 28080 16652
rect 28031 16612 28080 16640
rect 28031 16609 28043 16612
rect 27985 16603 28043 16609
rect 28074 16600 28080 16612
rect 28132 16600 28138 16652
rect 28258 16600 28264 16652
rect 28316 16600 28322 16652
rect 28353 16643 28411 16649
rect 28353 16609 28365 16643
rect 28399 16640 28411 16643
rect 28534 16640 28540 16652
rect 28399 16612 28540 16640
rect 28399 16609 28411 16612
rect 28353 16603 28411 16609
rect 28534 16600 28540 16612
rect 28592 16600 28598 16652
rect 28626 16600 28632 16652
rect 28684 16600 28690 16652
rect 29270 16600 29276 16652
rect 29328 16600 29334 16652
rect 29454 16600 29460 16652
rect 29512 16640 29518 16652
rect 29825 16643 29883 16649
rect 29825 16640 29837 16643
rect 29512 16612 29837 16640
rect 29512 16600 29518 16612
rect 29825 16609 29837 16612
rect 29871 16609 29883 16643
rect 29825 16603 29883 16609
rect 30009 16643 30067 16649
rect 30009 16609 30021 16643
rect 30055 16640 30067 16643
rect 30098 16640 30104 16652
rect 30055 16612 30104 16640
rect 30055 16609 30067 16612
rect 30009 16603 30067 16609
rect 30098 16600 30104 16612
rect 30156 16600 30162 16652
rect 31128 16649 31156 16748
rect 34514 16736 34520 16748
rect 34572 16736 34578 16788
rect 36265 16779 36323 16785
rect 36265 16745 36277 16779
rect 36311 16776 36323 16779
rect 36354 16776 36360 16788
rect 36311 16748 36360 16776
rect 36311 16745 36323 16748
rect 36265 16739 36323 16745
rect 36354 16736 36360 16748
rect 36412 16736 36418 16788
rect 40218 16736 40224 16788
rect 40276 16736 40282 16788
rect 41046 16736 41052 16788
rect 41104 16736 41110 16788
rect 41230 16736 41236 16788
rect 41288 16736 41294 16788
rect 48774 16736 48780 16788
rect 48832 16736 48838 16788
rect 31294 16668 31300 16720
rect 31352 16708 31358 16720
rect 34425 16711 34483 16717
rect 31352 16680 32352 16708
rect 31352 16668 31358 16680
rect 31113 16643 31171 16649
rect 31113 16609 31125 16643
rect 31159 16609 31171 16643
rect 31113 16603 31171 16609
rect 31205 16643 31263 16649
rect 31205 16609 31217 16643
rect 31251 16640 31263 16643
rect 31251 16612 31754 16640
rect 31251 16609 31263 16612
rect 31205 16603 31263 16609
rect 27341 16575 27399 16581
rect 27341 16541 27353 16575
rect 27387 16572 27399 16575
rect 28902 16572 28908 16584
rect 27387 16544 28908 16572
rect 27387 16541 27399 16544
rect 27341 16535 27399 16541
rect 28902 16532 28908 16544
rect 28960 16532 28966 16584
rect 31018 16572 31024 16584
rect 29288 16544 31024 16572
rect 26634 16476 26740 16504
rect 26712 16448 26740 16476
rect 26970 16464 26976 16516
rect 27028 16504 27034 16516
rect 29288 16504 29316 16544
rect 31018 16532 31024 16544
rect 31076 16532 31082 16584
rect 31726 16572 31754 16612
rect 32214 16600 32220 16652
rect 32272 16600 32278 16652
rect 32324 16640 32352 16680
rect 34425 16677 34437 16711
rect 34471 16708 34483 16711
rect 34974 16708 34980 16720
rect 34471 16680 34980 16708
rect 34471 16677 34483 16680
rect 34425 16671 34483 16677
rect 34974 16668 34980 16680
rect 35032 16668 35038 16720
rect 37550 16708 37556 16720
rect 35084 16680 37556 16708
rect 35084 16649 35112 16680
rect 37550 16668 37556 16680
rect 37608 16668 37614 16720
rect 40236 16708 40264 16736
rect 41509 16711 41567 16717
rect 41509 16708 41521 16711
rect 40236 16680 41521 16708
rect 41509 16677 41521 16680
rect 41555 16708 41567 16711
rect 41966 16708 41972 16720
rect 41555 16680 41972 16708
rect 41555 16677 41567 16680
rect 41509 16671 41567 16677
rect 41966 16668 41972 16680
rect 42024 16668 42030 16720
rect 35069 16643 35127 16649
rect 32324 16612 35020 16640
rect 31846 16572 31852 16584
rect 31726 16544 31852 16572
rect 31846 16532 31852 16544
rect 31904 16532 31910 16584
rect 34992 16572 35020 16612
rect 35069 16609 35081 16643
rect 35115 16609 35127 16643
rect 36725 16643 36783 16649
rect 36725 16640 36737 16643
rect 35069 16603 35127 16609
rect 35176 16612 36737 16640
rect 35176 16572 35204 16612
rect 36725 16609 36737 16612
rect 36771 16609 36783 16643
rect 36725 16603 36783 16609
rect 34992 16544 35204 16572
rect 35526 16532 35532 16584
rect 35584 16572 35590 16584
rect 35805 16575 35863 16581
rect 35805 16572 35817 16575
rect 35584 16544 35817 16572
rect 35584 16532 35590 16544
rect 35805 16541 35817 16544
rect 35851 16541 35863 16575
rect 36740 16572 36768 16603
rect 36814 16600 36820 16652
rect 36872 16600 36878 16652
rect 37277 16643 37335 16649
rect 37277 16640 37289 16643
rect 36924 16612 37289 16640
rect 36924 16572 36952 16612
rect 37277 16609 37289 16612
rect 37323 16609 37335 16643
rect 37277 16603 37335 16609
rect 37826 16600 37832 16652
rect 37884 16640 37890 16652
rect 38838 16640 38844 16652
rect 37884 16612 38844 16640
rect 37884 16600 37890 16612
rect 38838 16600 38844 16612
rect 38896 16640 38902 16652
rect 39209 16643 39267 16649
rect 39209 16640 39221 16643
rect 38896 16612 39221 16640
rect 38896 16600 38902 16612
rect 39209 16609 39221 16612
rect 39255 16609 39267 16643
rect 39209 16603 39267 16609
rect 40221 16643 40279 16649
rect 40221 16609 40233 16643
rect 40267 16640 40279 16643
rect 40310 16640 40316 16652
rect 40267 16612 40316 16640
rect 40267 16609 40279 16612
rect 40221 16603 40279 16609
rect 40310 16600 40316 16612
rect 40368 16600 40374 16652
rect 41046 16600 41052 16652
rect 41104 16640 41110 16652
rect 41104 16612 41414 16640
rect 41104 16600 41110 16612
rect 36740 16544 36952 16572
rect 35805 16535 35863 16541
rect 39482 16532 39488 16584
rect 39540 16572 39546 16584
rect 40678 16572 40684 16584
rect 39540 16544 40684 16572
rect 39540 16532 39546 16544
rect 40678 16532 40684 16544
rect 40736 16532 40742 16584
rect 41386 16572 41414 16612
rect 41598 16572 41604 16584
rect 41386 16544 41604 16572
rect 41598 16532 41604 16544
rect 41656 16532 41662 16584
rect 48593 16575 48651 16581
rect 48593 16541 48605 16575
rect 48639 16572 48651 16575
rect 49329 16575 49387 16581
rect 49329 16572 49341 16575
rect 48639 16544 49341 16572
rect 48639 16541 48651 16544
rect 48593 16535 48651 16541
rect 49329 16541 49341 16544
rect 49375 16572 49387 16575
rect 49418 16572 49424 16584
rect 49375 16544 49424 16572
rect 49375 16541 49387 16544
rect 49329 16535 49387 16541
rect 49418 16532 49424 16544
rect 49476 16532 49482 16584
rect 27028 16476 29316 16504
rect 27028 16464 27034 16476
rect 29362 16464 29368 16516
rect 29420 16504 29426 16516
rect 30101 16507 30159 16513
rect 30101 16504 30113 16507
rect 29420 16476 30113 16504
rect 29420 16464 29426 16476
rect 30101 16473 30113 16476
rect 30147 16473 30159 16507
rect 32214 16504 32220 16516
rect 30101 16467 30159 16473
rect 30484 16476 32220 16504
rect 25593 16439 25651 16445
rect 25593 16436 25605 16439
rect 25516 16408 25605 16436
rect 25593 16405 25605 16408
rect 25639 16436 25651 16439
rect 26142 16436 26148 16448
rect 25639 16408 26148 16436
rect 25639 16405 25651 16408
rect 25593 16399 25651 16405
rect 26142 16396 26148 16408
rect 26200 16396 26206 16448
rect 26234 16396 26240 16448
rect 26292 16436 26298 16448
rect 26694 16436 26700 16448
rect 26292 16408 26700 16436
rect 26292 16396 26298 16408
rect 26694 16396 26700 16408
rect 26752 16436 26758 16448
rect 27430 16436 27436 16448
rect 26752 16408 27436 16436
rect 26752 16396 26758 16408
rect 27430 16396 27436 16408
rect 27488 16436 27494 16448
rect 27617 16439 27675 16445
rect 27617 16436 27629 16439
rect 27488 16408 27629 16436
rect 27488 16396 27494 16408
rect 27617 16405 27629 16408
rect 27663 16405 27675 16439
rect 27617 16399 27675 16405
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 28626 16436 28632 16448
rect 28316 16408 28632 16436
rect 28316 16396 28322 16408
rect 28626 16396 28632 16408
rect 28684 16396 28690 16448
rect 30484 16445 30512 16476
rect 32214 16464 32220 16476
rect 32272 16464 32278 16516
rect 32398 16464 32404 16516
rect 32456 16504 32462 16516
rect 32493 16507 32551 16513
rect 32493 16504 32505 16507
rect 32456 16476 32505 16504
rect 32456 16464 32462 16476
rect 32493 16473 32505 16476
rect 32539 16473 32551 16507
rect 33870 16504 33876 16516
rect 33718 16476 33876 16504
rect 32493 16467 32551 16473
rect 33870 16464 33876 16476
rect 33928 16464 33934 16516
rect 35894 16504 35900 16516
rect 33980 16476 35900 16504
rect 33980 16448 34008 16476
rect 35894 16464 35900 16476
rect 35952 16464 35958 16516
rect 38654 16464 38660 16516
rect 38712 16464 38718 16516
rect 40218 16464 40224 16516
rect 40276 16504 40282 16516
rect 40313 16507 40371 16513
rect 40313 16504 40325 16507
rect 40276 16476 40325 16504
rect 40276 16464 40282 16476
rect 40313 16473 40325 16476
rect 40359 16473 40371 16507
rect 40313 16467 40371 16473
rect 40405 16507 40463 16513
rect 40405 16473 40417 16507
rect 40451 16504 40463 16507
rect 41230 16504 41236 16516
rect 40451 16476 41236 16504
rect 40451 16473 40463 16476
rect 40405 16467 40463 16473
rect 41230 16464 41236 16476
rect 41288 16464 41294 16516
rect 30469 16439 30527 16445
rect 30469 16405 30481 16439
rect 30515 16405 30527 16439
rect 30469 16399 30527 16405
rect 31294 16396 31300 16448
rect 31352 16396 31358 16448
rect 31662 16396 31668 16448
rect 31720 16396 31726 16448
rect 33962 16396 33968 16448
rect 34020 16396 34026 16448
rect 34054 16396 34060 16448
rect 34112 16436 34118 16448
rect 34330 16436 34336 16448
rect 34112 16408 34336 16436
rect 34112 16396 34118 16408
rect 34330 16396 34336 16408
rect 34388 16436 34394 16448
rect 36538 16436 36544 16448
rect 34388 16408 36544 16436
rect 34388 16396 34394 16408
rect 36538 16396 36544 16408
rect 36596 16396 36602 16448
rect 36633 16439 36691 16445
rect 36633 16405 36645 16439
rect 36679 16436 36691 16439
rect 36998 16436 37004 16448
rect 36679 16408 37004 16436
rect 36679 16405 36691 16408
rect 36633 16399 36691 16405
rect 36998 16396 37004 16408
rect 37056 16436 37062 16448
rect 37458 16436 37464 16448
rect 37056 16408 37464 16436
rect 37056 16396 37062 16408
rect 37458 16396 37464 16408
rect 37516 16396 37522 16448
rect 37737 16439 37795 16445
rect 37737 16405 37749 16439
rect 37783 16436 37795 16439
rect 38562 16436 38568 16448
rect 37783 16408 38568 16436
rect 37783 16405 37795 16408
rect 37737 16399 37795 16405
rect 38562 16396 38568 16408
rect 38620 16396 38626 16448
rect 40773 16439 40831 16445
rect 40773 16405 40785 16439
rect 40819 16436 40831 16439
rect 40954 16436 40960 16448
rect 40819 16408 40960 16436
rect 40819 16405 40831 16408
rect 40773 16399 40831 16405
rect 40954 16396 40960 16408
rect 41012 16396 41018 16448
rect 49142 16396 49148 16448
rect 49200 16396 49206 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 8294 16192 8300 16244
rect 8352 16192 8358 16244
rect 9214 16192 9220 16244
rect 9272 16192 9278 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11977 16235 12035 16241
rect 11977 16232 11989 16235
rect 11388 16204 11989 16232
rect 11388 16192 11394 16204
rect 11977 16201 11989 16204
rect 12023 16201 12035 16235
rect 11977 16195 12035 16201
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 13173 16235 13231 16241
rect 13173 16232 13185 16235
rect 12483 16204 13185 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 13173 16201 13185 16204
rect 13219 16201 13231 16235
rect 13173 16195 13231 16201
rect 13372 16204 14872 16232
rect 10870 16164 10876 16176
rect 2976 16136 10876 16164
rect 2976 16105 3004 16136
rect 10870 16124 10876 16136
rect 10928 16124 10934 16176
rect 11422 16124 11428 16176
rect 11480 16164 11486 16176
rect 13372 16164 13400 16204
rect 11480 16136 13400 16164
rect 13541 16167 13599 16173
rect 11480 16124 11486 16136
rect 13541 16133 13553 16167
rect 13587 16164 13599 16167
rect 13998 16164 14004 16176
rect 13587 16136 14004 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 14844 16173 14872 16204
rect 15102 16192 15108 16244
rect 15160 16232 15166 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15160 16204 15945 16232
rect 15160 16192 15166 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 15933 16195 15991 16201
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 16448 16204 17417 16232
rect 16448 16192 16454 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 17773 16235 17831 16241
rect 17773 16201 17785 16235
rect 17819 16232 17831 16235
rect 18322 16232 18328 16244
rect 17819 16204 18328 16232
rect 17819 16201 17831 16204
rect 17773 16195 17831 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 19392 16204 30604 16232
rect 19392 16192 19398 16204
rect 14829 16167 14887 16173
rect 14829 16133 14841 16167
rect 14875 16164 14887 16167
rect 16298 16164 16304 16176
rect 14875 16136 16304 16164
rect 14875 16133 14887 16136
rect 14829 16127 14887 16133
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 16850 16124 16856 16176
rect 16908 16164 16914 16176
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 16908 16136 17049 16164
rect 16908 16124 16914 16136
rect 17037 16133 17049 16136
rect 17083 16133 17095 16167
rect 17037 16127 17095 16133
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 17184 16136 19441 16164
rect 17184 16124 17190 16136
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 4304 16068 8217 16096
rect 4304 16056 4310 16068
rect 8205 16065 8217 16068
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10459 16068 11069 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 11698 16096 11704 16108
rect 11103 16068 11704 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 1026 15988 1032 16040
rect 1084 16028 1090 16040
rect 1765 16031 1823 16037
rect 1765 16028 1777 16031
rect 1084 16000 1777 16028
rect 1084 15988 1090 16000
rect 1765 15997 1777 16000
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 9030 16028 9036 16040
rect 8159 16000 9036 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 9324 16028 9352 16059
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16096 12403 16099
rect 13170 16096 13176 16108
rect 12391 16068 13176 16096
rect 12391 16065 12403 16068
rect 12345 16059 12403 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 14737 16099 14795 16105
rect 13320 16068 13492 16096
rect 13320 16056 13326 16068
rect 10778 16028 10784 16040
rect 9324 16000 10784 16028
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 12621 16031 12679 16037
rect 12621 16028 12633 16031
rect 11020 16000 12633 16028
rect 11020 15988 11026 16000
rect 12621 15997 12633 16000
rect 12667 16028 12679 16031
rect 13354 16028 13360 16040
rect 12667 16000 13360 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 13464 16028 13492 16068
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 13464 16000 13645 16028
rect 13633 15997 13645 16000
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 13725 16031 13783 16037
rect 13725 15997 13737 16031
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 8665 15963 8723 15969
rect 8665 15929 8677 15963
rect 8711 15960 8723 15963
rect 9766 15960 9772 15972
rect 8711 15932 9772 15960
rect 8711 15929 8723 15932
rect 8665 15923 8723 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 13740 15960 13768 15991
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14752 16028 14780 16059
rect 15010 16056 15016 16108
rect 15068 16096 15074 16108
rect 17770 16096 17776 16108
rect 15068 16068 17776 16096
rect 15068 16056 15074 16068
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 13872 16000 14780 16028
rect 13872 15988 13878 16000
rect 14826 15988 14832 16040
rect 14884 16028 14890 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14884 16000 14933 16028
rect 14884 15988 14890 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15562 15988 15568 16040
rect 15620 16028 15626 16040
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 15620 16000 15669 16028
rect 15620 15988 15626 16000
rect 15657 15997 15669 16000
rect 15703 15997 15715 16031
rect 15657 15991 15715 15997
rect 15838 15988 15844 16040
rect 15896 15988 15902 16040
rect 16761 16031 16819 16037
rect 16761 15997 16773 16031
rect 16807 16028 16819 16031
rect 17126 16028 17132 16040
rect 16807 16000 17132 16028
rect 16807 15997 16819 16000
rect 16761 15991 16819 15997
rect 17126 15988 17132 16000
rect 17184 15988 17190 16040
rect 17972 16037 18000 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 20898 16164 20904 16176
rect 20654 16136 20904 16164
rect 19429 16127 19487 16133
rect 20898 16124 20904 16136
rect 20956 16164 20962 16176
rect 21542 16164 21548 16176
rect 20956 16136 21548 16164
rect 20956 16124 20962 16136
rect 21542 16124 21548 16136
rect 21600 16124 21606 16176
rect 24762 16164 24768 16176
rect 23400 16136 24768 16164
rect 19150 16056 19156 16108
rect 19208 16056 19214 16108
rect 23400 16096 23428 16136
rect 24762 16124 24768 16136
rect 24820 16124 24826 16176
rect 25774 16164 25780 16176
rect 25622 16136 25780 16164
rect 25774 16124 25780 16136
rect 25832 16164 25838 16176
rect 26142 16164 26148 16176
rect 25832 16136 26148 16164
rect 25832 16124 25838 16136
rect 26142 16124 26148 16136
rect 26200 16124 26206 16176
rect 27798 16164 27804 16176
rect 26344 16136 27804 16164
rect 20732 16068 23428 16096
rect 17865 16031 17923 16037
rect 17865 15997 17877 16031
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 15997 18015 16031
rect 20622 16028 20628 16040
rect 17957 15991 18015 15997
rect 18064 16000 20628 16028
rect 13906 15960 13912 15972
rect 9876 15932 10640 15960
rect 13740 15932 13912 15960
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 9876 15892 9904 15932
rect 6880 15864 9904 15892
rect 6880 15852 6886 15864
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 10376 15864 10517 15892
rect 10376 15852 10382 15864
rect 10505 15861 10517 15864
rect 10551 15861 10563 15895
rect 10612 15892 10640 15932
rect 13906 15920 13912 15932
rect 13964 15920 13970 15972
rect 14274 15920 14280 15972
rect 14332 15960 14338 15972
rect 15286 15960 15292 15972
rect 14332 15932 15292 15960
rect 14332 15920 14338 15932
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 17586 15960 17592 15972
rect 16347 15932 17592 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 17586 15920 17592 15932
rect 17644 15920 17650 15972
rect 17880 15960 17908 15991
rect 18064 15960 18092 16000
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 17880 15932 18092 15960
rect 18156 15932 19012 15960
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10612 15864 10977 15892
rect 10505 15855 10563 15861
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11480 15864 11621 15892
rect 11480 15852 11486 15864
rect 11609 15861 11621 15864
rect 11655 15861 11667 15895
rect 11609 15855 11667 15861
rect 12710 15852 12716 15904
rect 12768 15892 12774 15904
rect 12894 15892 12900 15904
rect 12768 15864 12900 15892
rect 12768 15852 12774 15864
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 14369 15895 14427 15901
rect 14369 15892 14381 15895
rect 14056 15864 14381 15892
rect 14056 15852 14062 15864
rect 14369 15861 14381 15864
rect 14415 15861 14427 15895
rect 14369 15855 14427 15861
rect 16942 15852 16948 15904
rect 17000 15852 17006 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 18156 15892 18184 15932
rect 17368 15864 18184 15892
rect 17368 15852 17374 15864
rect 18874 15852 18880 15904
rect 18932 15852 18938 15904
rect 18984 15892 19012 15932
rect 20732 15892 20760 16068
rect 23474 16056 23480 16108
rect 23532 16056 23538 16108
rect 26344 16105 26372 16136
rect 27798 16124 27804 16136
rect 27856 16164 27862 16176
rect 28902 16164 28908 16176
rect 27856 16136 28908 16164
rect 27856 16124 27862 16136
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 26694 16056 26700 16108
rect 26752 16056 26758 16108
rect 27338 16056 27344 16108
rect 27396 16096 27402 16108
rect 28368 16105 28396 16136
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 30576 16164 30604 16204
rect 30650 16192 30656 16244
rect 30708 16232 30714 16244
rect 30929 16235 30987 16241
rect 30929 16232 30941 16235
rect 30708 16204 30941 16232
rect 30708 16192 30714 16204
rect 30929 16201 30941 16204
rect 30975 16201 30987 16235
rect 30929 16195 30987 16201
rect 31754 16192 31760 16244
rect 31812 16232 31818 16244
rect 33781 16235 33839 16241
rect 33781 16232 33793 16235
rect 31812 16204 33793 16232
rect 31812 16192 31818 16204
rect 33781 16201 33793 16204
rect 33827 16201 33839 16235
rect 33781 16195 33839 16201
rect 34790 16192 34796 16244
rect 34848 16232 34854 16244
rect 34848 16204 36952 16232
rect 34848 16192 34854 16204
rect 31662 16164 31668 16176
rect 30576 16136 31668 16164
rect 31662 16124 31668 16136
rect 31720 16164 31726 16176
rect 32030 16164 32036 16176
rect 31720 16136 32036 16164
rect 31720 16124 31726 16136
rect 32030 16124 32036 16136
rect 32088 16124 32094 16176
rect 34517 16167 34575 16173
rect 34517 16164 34529 16167
rect 32600 16136 34529 16164
rect 27525 16099 27583 16105
rect 27525 16096 27537 16099
rect 27396 16068 27537 16096
rect 27396 16056 27402 16068
rect 27525 16065 27537 16068
rect 27571 16065 27583 16099
rect 27525 16059 27583 16065
rect 27617 16099 27675 16105
rect 27617 16065 27629 16099
rect 27663 16096 27675 16099
rect 28353 16099 28411 16105
rect 27663 16068 27844 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 23293 16031 23351 16037
rect 23293 15997 23305 16031
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 20898 15920 20904 15972
rect 20956 15960 20962 15972
rect 21358 15960 21364 15972
rect 20956 15932 21364 15960
rect 20956 15920 20962 15932
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 22741 15963 22799 15969
rect 22741 15960 22753 15963
rect 21560 15932 22753 15960
rect 21560 15904 21588 15932
rect 22741 15929 22753 15932
rect 22787 15929 22799 15963
rect 23308 15960 23336 15991
rect 23382 15988 23388 16040
rect 23440 15988 23446 16040
rect 24578 16028 24584 16040
rect 23492 16000 24584 16028
rect 23492 15960 23520 16000
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 26050 15988 26056 16040
rect 26108 15988 26114 16040
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 23308 15932 23520 15960
rect 23845 15963 23903 15969
rect 22741 15923 22799 15929
rect 23845 15929 23857 15963
rect 23891 15960 23903 15963
rect 24854 15960 24860 15972
rect 23891 15932 24860 15960
rect 23891 15929 23903 15932
rect 23845 15923 23903 15929
rect 24854 15920 24860 15932
rect 24912 15920 24918 15972
rect 27338 15920 27344 15972
rect 27396 15960 27402 15972
rect 27724 15960 27752 15991
rect 27396 15932 27752 15960
rect 27396 15920 27402 15932
rect 18984 15864 20760 15892
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21542 15892 21548 15904
rect 21315 15864 21548 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 21818 15852 21824 15904
rect 21876 15892 21882 15904
rect 22462 15892 22468 15904
rect 21876 15864 22468 15892
rect 21876 15852 21882 15864
rect 22462 15852 22468 15864
rect 22520 15852 22526 15904
rect 26694 15852 26700 15904
rect 26752 15892 26758 15904
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 26752 15864 27169 15892
rect 26752 15852 26758 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27816 15892 27844 16068
rect 28353 16065 28365 16099
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 28626 15988 28632 16040
rect 28684 15988 28690 16040
rect 28994 15988 29000 16040
rect 29052 16028 29058 16040
rect 29362 16028 29368 16040
rect 29052 16000 29368 16028
rect 29052 15988 29058 16000
rect 29362 15988 29368 16000
rect 29420 16028 29426 16040
rect 29748 16028 29776 16082
rect 30098 16056 30104 16108
rect 30156 16096 30162 16108
rect 30156 16068 30788 16096
rect 30156 16056 30162 16068
rect 29420 16000 29776 16028
rect 29420 15988 29426 16000
rect 29748 15960 29776 16000
rect 29822 15988 29828 16040
rect 29880 16028 29886 16040
rect 30653 16031 30711 16037
rect 30653 16028 30665 16031
rect 29880 16000 30665 16028
rect 29880 15988 29886 16000
rect 30653 15997 30665 16000
rect 30699 15997 30711 16031
rect 30760 16028 30788 16068
rect 30834 16056 30840 16108
rect 30892 16056 30898 16108
rect 31018 16056 31024 16108
rect 31076 16096 31082 16108
rect 32600 16105 32628 16136
rect 34517 16133 34529 16136
rect 34563 16133 34575 16167
rect 34517 16127 34575 16133
rect 34974 16124 34980 16176
rect 35032 16164 35038 16176
rect 35032 16136 35466 16164
rect 35032 16124 35038 16136
rect 32585 16099 32643 16105
rect 32585 16096 32597 16099
rect 31076 16068 32597 16096
rect 31076 16056 31082 16068
rect 32585 16065 32597 16068
rect 32631 16065 32643 16099
rect 32585 16059 32643 16065
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16065 32735 16099
rect 32677 16059 32735 16065
rect 31386 16028 31392 16040
rect 30760 16000 31392 16028
rect 30653 15991 30711 15997
rect 31386 15988 31392 16000
rect 31444 15988 31450 16040
rect 32490 15988 32496 16040
rect 32548 15988 32554 16040
rect 32692 15960 32720 16059
rect 33318 16056 33324 16108
rect 33376 16096 33382 16108
rect 36924 16105 36952 16204
rect 37182 16192 37188 16244
rect 37240 16232 37246 16244
rect 40497 16235 40555 16241
rect 40497 16232 40509 16235
rect 37240 16204 40509 16232
rect 37240 16192 37246 16204
rect 40497 16201 40509 16204
rect 40543 16201 40555 16235
rect 40497 16195 40555 16201
rect 40954 16192 40960 16244
rect 41012 16192 41018 16244
rect 38473 16167 38531 16173
rect 38473 16133 38485 16167
rect 38519 16164 38531 16167
rect 38562 16164 38568 16176
rect 38519 16136 38568 16164
rect 38519 16133 38531 16136
rect 38473 16127 38531 16133
rect 38562 16124 38568 16136
rect 38620 16124 38626 16176
rect 39942 16164 39948 16176
rect 39698 16136 39948 16164
rect 39942 16124 39948 16136
rect 40000 16124 40006 16176
rect 33873 16099 33931 16105
rect 33873 16096 33885 16099
rect 33376 16068 33885 16096
rect 33376 16056 33382 16068
rect 33873 16065 33885 16068
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 36909 16099 36967 16105
rect 36909 16065 36921 16099
rect 36955 16096 36967 16099
rect 37366 16096 37372 16108
rect 36955 16068 37372 16096
rect 36955 16065 36967 16068
rect 36909 16059 36967 16065
rect 37366 16056 37372 16068
rect 37424 16096 37430 16108
rect 38197 16099 38255 16105
rect 38197 16096 38209 16099
rect 37424 16068 38209 16096
rect 37424 16056 37430 16068
rect 38197 16065 38209 16068
rect 38243 16065 38255 16099
rect 38197 16059 38255 16065
rect 40865 16099 40923 16105
rect 40865 16065 40877 16099
rect 40911 16096 40923 16099
rect 48682 16096 48688 16108
rect 40911 16068 48688 16096
rect 40911 16065 40923 16068
rect 40865 16059 40923 16065
rect 48682 16056 48688 16068
rect 48740 16056 48746 16108
rect 48777 16099 48835 16105
rect 48777 16065 48789 16099
rect 48823 16096 48835 16099
rect 49326 16096 49332 16108
rect 48823 16068 49332 16096
rect 48823 16065 48835 16068
rect 48777 16059 48835 16065
rect 49326 16056 49332 16068
rect 49384 16056 49390 16108
rect 32766 15988 32772 16040
rect 32824 16028 32830 16040
rect 33597 16031 33655 16037
rect 33597 16028 33609 16031
rect 32824 16000 33609 16028
rect 32824 15988 32830 16000
rect 33597 15997 33609 16000
rect 33643 15997 33655 16031
rect 36262 16028 36268 16040
rect 33597 15991 33655 15997
rect 35544 16000 36268 16028
rect 35544 15972 35572 16000
rect 36262 15988 36268 16000
rect 36320 15988 36326 16040
rect 36633 16031 36691 16037
rect 36633 15997 36645 16031
rect 36679 16028 36691 16031
rect 37274 16028 37280 16040
rect 36679 16000 37280 16028
rect 36679 15997 36691 16000
rect 36633 15991 36691 15997
rect 37274 15988 37280 16000
rect 37332 15988 37338 16040
rect 37458 15988 37464 16040
rect 37516 15988 37522 16040
rect 39206 15988 39212 16040
rect 39264 16028 39270 16040
rect 41049 16031 41107 16037
rect 41049 16028 41061 16031
rect 39264 16000 41061 16028
rect 39264 15988 39270 16000
rect 41049 15997 41061 16000
rect 41095 16028 41107 16031
rect 41782 16028 41788 16040
rect 41095 16000 41788 16028
rect 41095 15997 41107 16000
rect 41049 15991 41107 15997
rect 41782 15988 41788 16000
rect 41840 15988 41846 16040
rect 33410 15960 33416 15972
rect 29748 15932 31708 15960
rect 32692 15932 33416 15960
rect 28626 15892 28632 15904
rect 27816 15864 28632 15892
rect 27157 15855 27215 15861
rect 28626 15852 28632 15864
rect 28684 15852 28690 15904
rect 30101 15895 30159 15901
rect 30101 15861 30113 15895
rect 30147 15892 30159 15895
rect 30742 15892 30748 15904
rect 30147 15864 30748 15892
rect 30147 15861 30159 15864
rect 30101 15855 30159 15861
rect 30742 15852 30748 15864
rect 30800 15852 30806 15904
rect 31297 15895 31355 15901
rect 31297 15861 31309 15895
rect 31343 15892 31355 15895
rect 31386 15892 31392 15904
rect 31343 15864 31392 15892
rect 31343 15861 31355 15864
rect 31297 15855 31355 15861
rect 31386 15852 31392 15864
rect 31444 15852 31450 15904
rect 31680 15901 31708 15932
rect 33410 15920 33416 15932
rect 33468 15960 33474 15972
rect 34330 15960 34336 15972
rect 33468 15932 34336 15960
rect 33468 15920 33474 15932
rect 34330 15920 34336 15932
rect 34388 15960 34394 15972
rect 34701 15963 34759 15969
rect 34701 15960 34713 15963
rect 34388 15932 34713 15960
rect 34388 15920 34394 15932
rect 34701 15929 34713 15932
rect 34747 15929 34759 15963
rect 34701 15923 34759 15929
rect 35526 15920 35532 15972
rect 35584 15920 35590 15972
rect 49142 15920 49148 15972
rect 49200 15920 49206 15972
rect 31665 15895 31723 15901
rect 31665 15861 31677 15895
rect 31711 15892 31723 15895
rect 31754 15892 31760 15904
rect 31711 15864 31760 15892
rect 31711 15861 31723 15864
rect 31665 15855 31723 15861
rect 31754 15852 31760 15864
rect 31812 15852 31818 15904
rect 31846 15852 31852 15904
rect 31904 15892 31910 15904
rect 32674 15892 32680 15904
rect 31904 15864 32680 15892
rect 31904 15852 31910 15864
rect 32674 15852 32680 15864
rect 32732 15852 32738 15904
rect 33045 15895 33103 15901
rect 33045 15861 33057 15895
rect 33091 15892 33103 15895
rect 33686 15892 33692 15904
rect 33091 15864 33692 15892
rect 33091 15861 33103 15864
rect 33045 15855 33103 15861
rect 33686 15852 33692 15864
rect 33744 15852 33750 15904
rect 34241 15895 34299 15901
rect 34241 15861 34253 15895
rect 34287 15892 34299 15895
rect 34606 15892 34612 15904
rect 34287 15864 34612 15892
rect 34287 15861 34299 15864
rect 34241 15855 34299 15861
rect 34606 15852 34612 15864
rect 34664 15852 34670 15904
rect 35158 15852 35164 15904
rect 35216 15892 35222 15904
rect 36814 15892 36820 15904
rect 35216 15864 36820 15892
rect 35216 15852 35222 15864
rect 36814 15852 36820 15864
rect 36872 15852 36878 15904
rect 39945 15895 40003 15901
rect 39945 15861 39957 15895
rect 39991 15892 40003 15895
rect 40310 15892 40316 15904
rect 39991 15864 40316 15892
rect 39991 15861 40003 15864
rect 39945 15855 40003 15861
rect 40310 15852 40316 15864
rect 40368 15852 40374 15904
rect 41598 15852 41604 15904
rect 41656 15892 41662 15904
rect 42058 15892 42064 15904
rect 41656 15864 42064 15892
rect 41656 15852 41662 15864
rect 42058 15852 42064 15864
rect 42116 15852 42122 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10744 15660 10793 15688
rect 10744 15648 10750 15660
rect 10781 15657 10793 15660
rect 10827 15688 10839 15691
rect 10962 15688 10968 15700
rect 10827 15660 10968 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 12158 15648 12164 15700
rect 12216 15688 12222 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 12216 15660 14289 15688
rect 12216 15648 12222 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 16574 15648 16580 15700
rect 16632 15688 16638 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 16632 15660 16773 15688
rect 16632 15648 16638 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 16761 15651 16819 15657
rect 17862 15648 17868 15700
rect 17920 15648 17926 15700
rect 18049 15691 18107 15697
rect 18049 15657 18061 15691
rect 18095 15688 18107 15691
rect 18782 15688 18788 15700
rect 18095 15660 18788 15688
rect 18095 15657 18107 15660
rect 18049 15651 18107 15657
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 18966 15648 18972 15700
rect 19024 15648 19030 15700
rect 19337 15691 19395 15697
rect 19337 15657 19349 15691
rect 19383 15688 19395 15691
rect 19518 15688 19524 15700
rect 19383 15660 19524 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 19886 15648 19892 15700
rect 19944 15648 19950 15700
rect 20806 15648 20812 15700
rect 20864 15688 20870 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20864 15660 21189 15688
rect 20864 15648 20870 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 21177 15651 21235 15657
rect 21358 15648 21364 15700
rect 21416 15688 21422 15700
rect 21416 15660 24072 15688
rect 21416 15648 21422 15660
rect 12894 15620 12900 15632
rect 12452 15592 12900 15620
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12452 15552 12480 15592
rect 12894 15580 12900 15592
rect 12952 15580 12958 15632
rect 15102 15620 15108 15632
rect 13188 15592 15108 15620
rect 12299 15524 12480 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12526 15512 12532 15564
rect 12584 15512 12590 15564
rect 13188 15561 13216 15592
rect 15102 15580 15108 15592
rect 15160 15580 15166 15632
rect 15378 15580 15384 15632
rect 15436 15620 15442 15632
rect 15838 15620 15844 15632
rect 15436 15592 15844 15620
rect 15436 15580 15442 15592
rect 15838 15580 15844 15592
rect 15896 15620 15902 15632
rect 15896 15592 17356 15620
rect 15896 15580 15902 15592
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 14918 15512 14924 15564
rect 14976 15512 14982 15564
rect 15562 15512 15568 15564
rect 15620 15552 15626 15564
rect 16114 15552 16120 15564
rect 15620 15524 16120 15552
rect 15620 15512 15626 15524
rect 16114 15512 16120 15524
rect 16172 15552 16178 15564
rect 16390 15552 16396 15564
rect 16172 15524 16396 15552
rect 16172 15512 16178 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 17328 15561 17356 15592
rect 18414 15580 18420 15632
rect 18472 15580 18478 15632
rect 21910 15620 21916 15632
rect 20364 15592 21916 15620
rect 20364 15561 20392 15592
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 22462 15580 22468 15632
rect 22520 15620 22526 15632
rect 23842 15620 23848 15632
rect 22520 15592 23848 15620
rect 22520 15580 22526 15592
rect 23842 15580 23848 15592
rect 23900 15580 23906 15632
rect 24044 15564 24072 15660
rect 26050 15648 26056 15700
rect 26108 15688 26114 15700
rect 26786 15688 26792 15700
rect 26108 15660 26792 15688
rect 26108 15648 26114 15660
rect 26786 15648 26792 15660
rect 26844 15688 26850 15700
rect 27065 15691 27123 15697
rect 27065 15688 27077 15691
rect 26844 15660 27077 15688
rect 26844 15648 26850 15660
rect 27065 15657 27077 15660
rect 27111 15657 27123 15691
rect 27065 15651 27123 15657
rect 30190 15648 30196 15700
rect 30248 15688 30254 15700
rect 34333 15691 34391 15697
rect 30248 15660 32996 15688
rect 30248 15648 30254 15660
rect 27522 15620 27528 15632
rect 25240 15592 27528 15620
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 20349 15555 20407 15561
rect 20349 15521 20361 15555
rect 20395 15521 20407 15555
rect 20349 15515 20407 15521
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 21358 15552 21364 15564
rect 20579 15524 21364 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 21729 15555 21787 15561
rect 21729 15552 21741 15555
rect 21508 15524 21741 15552
rect 21508 15512 21514 15524
rect 21729 15521 21741 15524
rect 21775 15521 21787 15555
rect 23290 15552 23296 15564
rect 21729 15515 21787 15521
rect 21836 15524 23296 15552
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 10226 15484 10232 15496
rect 3007 15456 10232 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 13265 15487 13323 15493
rect 13265 15484 13277 15487
rect 12676 15456 13277 15484
rect 12676 15444 12682 15456
rect 13265 15453 13277 15456
rect 13311 15453 13323 15487
rect 13265 15447 13323 15453
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13446 15484 13452 15496
rect 13403 15456 13452 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 13722 15444 13728 15496
rect 13780 15444 13786 15496
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 18414 15484 18420 15496
rect 14783 15456 18420 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 21836 15484 21864 15524
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 23753 15555 23811 15561
rect 23753 15521 23765 15555
rect 23799 15552 23811 15555
rect 23934 15552 23940 15564
rect 23799 15524 23940 15552
rect 23799 15521 23811 15524
rect 23753 15515 23811 15521
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 24026 15512 24032 15564
rect 24084 15552 24090 15564
rect 25240 15561 25268 15592
rect 27522 15580 27528 15592
rect 27580 15580 27586 15632
rect 32217 15623 32275 15629
rect 32217 15589 32229 15623
rect 32263 15620 32275 15623
rect 32582 15620 32588 15632
rect 32263 15592 32588 15620
rect 32263 15589 32275 15592
rect 32217 15583 32275 15589
rect 32582 15580 32588 15592
rect 32640 15580 32646 15632
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 24084 15524 25237 15552
rect 24084 15512 24090 15524
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25225 15515 25283 15521
rect 25314 15512 25320 15564
rect 25372 15552 25378 15564
rect 26421 15555 26479 15561
rect 26421 15552 26433 15555
rect 25372 15524 26433 15552
rect 25372 15512 25378 15524
rect 26421 15521 26433 15524
rect 26467 15521 26479 15555
rect 26421 15515 26479 15521
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 26660 15524 27997 15552
rect 26660 15512 26666 15524
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 30469 15555 30527 15561
rect 30469 15521 30481 15555
rect 30515 15552 30527 15555
rect 31110 15552 31116 15564
rect 30515 15524 31116 15552
rect 30515 15521 30527 15524
rect 30469 15515 30527 15521
rect 31110 15512 31116 15524
rect 31168 15512 31174 15564
rect 31478 15512 31484 15564
rect 31536 15552 31542 15564
rect 32398 15552 32404 15564
rect 31536 15524 32404 15552
rect 31536 15512 31542 15524
rect 32398 15512 32404 15524
rect 32456 15512 32462 15564
rect 32968 15561 32996 15660
rect 34333 15657 34345 15691
rect 34379 15688 34391 15691
rect 34974 15688 34980 15700
rect 34379 15660 34980 15688
rect 34379 15657 34391 15660
rect 34333 15651 34391 15657
rect 34974 15648 34980 15660
rect 35032 15648 35038 15700
rect 35618 15648 35624 15700
rect 35676 15688 35682 15700
rect 36633 15691 36691 15697
rect 35676 15660 36308 15688
rect 35676 15648 35682 15660
rect 33413 15623 33471 15629
rect 33413 15589 33425 15623
rect 33459 15620 33471 15623
rect 34422 15620 34428 15632
rect 33459 15592 34428 15620
rect 33459 15589 33471 15592
rect 33413 15583 33471 15589
rect 34422 15580 34428 15592
rect 34480 15580 34486 15632
rect 36280 15620 36308 15660
rect 36633 15657 36645 15691
rect 36679 15688 36691 15691
rect 37274 15688 37280 15700
rect 36679 15660 37280 15688
rect 36679 15657 36691 15660
rect 36633 15651 36691 15657
rect 37274 15648 37280 15660
rect 37332 15648 37338 15700
rect 37734 15648 37740 15700
rect 37792 15648 37798 15700
rect 41782 15648 41788 15700
rect 41840 15648 41846 15700
rect 42058 15648 42064 15700
rect 42116 15648 42122 15700
rect 48682 15648 48688 15700
rect 48740 15688 48746 15700
rect 49145 15691 49203 15697
rect 49145 15688 49157 15691
rect 48740 15660 49157 15688
rect 48740 15648 48746 15660
rect 49145 15657 49157 15660
rect 49191 15657 49203 15691
rect 49145 15651 49203 15657
rect 37458 15620 37464 15632
rect 36280 15592 37464 15620
rect 37458 15580 37464 15592
rect 37516 15580 37522 15632
rect 32861 15555 32919 15561
rect 32861 15521 32873 15555
rect 32907 15521 32919 15555
rect 32861 15515 32919 15521
rect 32953 15555 33011 15561
rect 32953 15521 32965 15555
rect 32999 15521 33011 15555
rect 32953 15515 33011 15521
rect 18647 15456 21864 15484
rect 23569 15487 23627 15493
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 27154 15484 27160 15496
rect 23615 15456 27160 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27706 15444 27712 15496
rect 27764 15484 27770 15496
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27764 15456 27813 15484
rect 27764 15444 27770 15456
rect 27801 15453 27813 15456
rect 27847 15484 27859 15487
rect 28445 15487 28503 15493
rect 28445 15484 28457 15487
rect 27847 15456 28457 15484
rect 27847 15453 27859 15456
rect 27801 15447 27859 15453
rect 28445 15453 28457 15456
rect 28491 15453 28503 15487
rect 28445 15447 28503 15453
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15484 29055 15487
rect 29043 15456 30512 15484
rect 29043 15453 29055 15456
rect 28997 15447 29055 15453
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 1765 15419 1823 15425
rect 1765 15416 1777 15419
rect 992 15388 1777 15416
rect 992 15376 998 15388
rect 1765 15385 1777 15388
rect 1811 15385 1823 15419
rect 1765 15379 1823 15385
rect 4706 15376 4712 15428
rect 4764 15416 4770 15428
rect 6365 15419 6423 15425
rect 6365 15416 6377 15419
rect 4764 15388 6377 15416
rect 4764 15376 4770 15388
rect 6365 15385 6377 15388
rect 6411 15385 6423 15419
rect 6365 15379 6423 15385
rect 6549 15419 6607 15425
rect 6549 15385 6561 15419
rect 6595 15416 6607 15419
rect 10505 15419 10563 15425
rect 6595 15388 10364 15416
rect 6595 15385 6607 15388
rect 6549 15379 6607 15385
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 10336 15348 10364 15388
rect 10505 15385 10517 15419
rect 10551 15416 10563 15419
rect 10962 15416 10968 15428
rect 10551 15388 10968 15416
rect 10551 15385 10563 15388
rect 10505 15379 10563 15385
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 11974 15416 11980 15428
rect 11822 15388 11980 15416
rect 11974 15376 11980 15388
rect 12032 15416 12038 15428
rect 12526 15416 12532 15428
rect 12032 15388 12532 15416
rect 12032 15376 12038 15388
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 13740 15416 13768 15444
rect 15933 15419 15991 15425
rect 15933 15416 15945 15419
rect 13740 15388 15945 15416
rect 15933 15385 15945 15388
rect 15979 15416 15991 15419
rect 16758 15416 16764 15428
rect 15979 15388 16764 15416
rect 15979 15385 15991 15388
rect 15933 15379 15991 15385
rect 16758 15376 16764 15388
rect 16816 15376 16822 15428
rect 17126 15376 17132 15428
rect 17184 15376 17190 15428
rect 17221 15419 17279 15425
rect 17221 15385 17233 15419
rect 17267 15416 17279 15419
rect 17862 15416 17868 15428
rect 17267 15388 17868 15416
rect 17267 15385 17279 15388
rect 17221 15379 17279 15385
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 21266 15416 21272 15428
rect 18708 15388 21272 15416
rect 18708 15360 18736 15388
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 21545 15419 21603 15425
rect 21545 15385 21557 15419
rect 21591 15416 21603 15419
rect 21591 15388 21864 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 11882 15348 11888 15360
rect 10336 15320 11888 15348
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 13538 15308 13544 15360
rect 13596 15348 13602 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13596 15320 13737 15348
rect 13596 15308 13602 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 14642 15308 14648 15360
rect 14700 15308 14706 15360
rect 15562 15308 15568 15360
rect 15620 15308 15626 15360
rect 16025 15351 16083 15357
rect 16025 15317 16037 15351
rect 16071 15348 16083 15351
rect 16298 15348 16304 15360
rect 16071 15320 16304 15348
rect 16071 15317 16083 15320
rect 16025 15311 16083 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 18690 15348 18696 15360
rect 16448 15320 18696 15348
rect 16448 15308 16454 15320
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 19978 15348 19984 15360
rect 19567 15320 19984 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20254 15308 20260 15360
rect 20312 15308 20318 15360
rect 20346 15308 20352 15360
rect 20404 15348 20410 15360
rect 20898 15348 20904 15360
rect 20404 15320 20904 15348
rect 20404 15308 20410 15320
rect 20898 15308 20904 15320
rect 20956 15308 20962 15360
rect 21450 15308 21456 15360
rect 21508 15348 21514 15360
rect 21637 15351 21695 15357
rect 21637 15348 21649 15351
rect 21508 15320 21649 15348
rect 21508 15308 21514 15320
rect 21637 15317 21649 15320
rect 21683 15317 21695 15351
rect 21836 15348 21864 15388
rect 21910 15376 21916 15428
rect 21968 15416 21974 15428
rect 23477 15419 23535 15425
rect 21968 15388 23152 15416
rect 21968 15376 21974 15388
rect 22186 15348 22192 15360
rect 21836 15320 22192 15348
rect 21637 15311 21695 15317
rect 22186 15308 22192 15320
rect 22244 15308 22250 15360
rect 23124 15357 23152 15388
rect 23477 15385 23489 15419
rect 23523 15416 23535 15419
rect 25041 15419 25099 15425
rect 23523 15388 24716 15416
rect 23523 15385 23535 15388
rect 23477 15379 23535 15385
rect 24688 15357 24716 15388
rect 25041 15385 25053 15419
rect 25087 15416 25099 15419
rect 25958 15416 25964 15428
rect 25087 15388 25964 15416
rect 25087 15385 25099 15388
rect 25041 15379 25099 15385
rect 25958 15376 25964 15388
rect 26016 15376 26022 15428
rect 26326 15376 26332 15428
rect 26384 15416 26390 15428
rect 27246 15416 27252 15428
rect 26384 15388 27252 15416
rect 26384 15376 26390 15388
rect 27246 15376 27252 15388
rect 27304 15376 27310 15428
rect 27893 15419 27951 15425
rect 27893 15385 27905 15419
rect 27939 15416 27951 15419
rect 28350 15416 28356 15428
rect 27939 15388 28356 15416
rect 27939 15385 27951 15388
rect 27893 15379 27951 15385
rect 28350 15376 28356 15388
rect 28408 15416 28414 15428
rect 28629 15419 28687 15425
rect 28629 15416 28641 15419
rect 28408 15388 28641 15416
rect 28408 15376 28414 15388
rect 28629 15385 28641 15388
rect 28675 15385 28687 15419
rect 28629 15379 28687 15385
rect 29181 15419 29239 15425
rect 29181 15385 29193 15419
rect 29227 15416 29239 15419
rect 30098 15416 30104 15428
rect 29227 15388 30104 15416
rect 29227 15385 29239 15388
rect 29181 15379 29239 15385
rect 30098 15376 30104 15388
rect 30156 15376 30162 15428
rect 30484 15416 30512 15456
rect 31846 15444 31852 15496
rect 31904 15444 31910 15496
rect 32876 15484 32904 15515
rect 34790 15512 34796 15564
rect 34848 15552 34854 15564
rect 34885 15555 34943 15561
rect 34885 15552 34897 15555
rect 34848 15524 34897 15552
rect 34848 15512 34854 15524
rect 34885 15521 34897 15524
rect 34931 15521 34943 15555
rect 34885 15515 34943 15521
rect 35161 15555 35219 15561
rect 35161 15521 35173 15555
rect 35207 15552 35219 15555
rect 35894 15552 35900 15564
rect 35207 15524 35900 15552
rect 35207 15521 35219 15524
rect 35161 15515 35219 15521
rect 35894 15512 35900 15524
rect 35952 15512 35958 15564
rect 37366 15512 37372 15564
rect 37424 15552 37430 15564
rect 39482 15552 39488 15564
rect 37424 15524 39488 15552
rect 37424 15512 37430 15524
rect 39482 15512 39488 15524
rect 39540 15552 39546 15564
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 39540 15524 40049 15552
rect 39540 15512 39546 15524
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 40310 15512 40316 15564
rect 40368 15512 40374 15564
rect 34054 15484 34060 15496
rect 32876 15456 34060 15484
rect 34054 15444 34060 15456
rect 34112 15444 34118 15496
rect 48869 15487 48927 15493
rect 48869 15453 48881 15487
rect 48915 15484 48927 15487
rect 49326 15484 49332 15496
rect 48915 15456 49332 15484
rect 48915 15453 48927 15456
rect 48869 15447 48927 15453
rect 49326 15444 49332 15456
rect 49384 15444 49390 15496
rect 30650 15416 30656 15428
rect 30484 15388 30656 15416
rect 30650 15376 30656 15388
rect 30708 15376 30714 15428
rect 30742 15376 30748 15428
rect 30800 15376 30806 15428
rect 35066 15376 35072 15428
rect 35124 15416 35130 15428
rect 35124 15388 35650 15416
rect 35124 15376 35130 15388
rect 35360 15360 35388 15388
rect 38654 15376 38660 15428
rect 38712 15376 38718 15428
rect 39206 15376 39212 15428
rect 39264 15376 39270 15428
rect 39942 15376 39948 15428
rect 40000 15416 40006 15428
rect 40000 15388 40802 15416
rect 40000 15376 40006 15388
rect 23109 15351 23167 15357
rect 23109 15317 23121 15351
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 24673 15351 24731 15357
rect 24673 15317 24685 15351
rect 24719 15317 24731 15351
rect 24673 15311 24731 15317
rect 25133 15351 25191 15357
rect 25133 15317 25145 15351
rect 25179 15348 25191 15351
rect 25222 15348 25228 15360
rect 25179 15320 25228 15348
rect 25179 15317 25191 15320
rect 25133 15311 25191 15317
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 25866 15308 25872 15360
rect 25924 15308 25930 15360
rect 26237 15351 26295 15357
rect 26237 15317 26249 15351
rect 26283 15348 26295 15351
rect 26418 15348 26424 15360
rect 26283 15320 26424 15348
rect 26283 15317 26295 15320
rect 26237 15311 26295 15317
rect 26418 15308 26424 15320
rect 26476 15348 26482 15360
rect 26970 15348 26976 15360
rect 26476 15320 26976 15348
rect 26476 15308 26482 15320
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 27430 15308 27436 15360
rect 27488 15308 27494 15360
rect 29362 15308 29368 15360
rect 29420 15308 29426 15360
rect 30009 15351 30067 15357
rect 30009 15317 30021 15351
rect 30055 15348 30067 15351
rect 30834 15348 30840 15360
rect 30055 15320 30840 15348
rect 30055 15317 30067 15320
rect 30009 15311 30067 15317
rect 30834 15308 30840 15320
rect 30892 15308 30898 15360
rect 32306 15308 32312 15360
rect 32364 15348 32370 15360
rect 33045 15351 33103 15357
rect 33045 15348 33057 15351
rect 32364 15320 33057 15348
rect 32364 15308 32370 15320
rect 33045 15317 33057 15320
rect 33091 15348 33103 15351
rect 33502 15348 33508 15360
rect 33091 15320 33508 15348
rect 33091 15317 33103 15320
rect 33045 15311 33103 15317
rect 33502 15308 33508 15320
rect 33560 15308 33566 15360
rect 33870 15308 33876 15360
rect 33928 15308 33934 15360
rect 35342 15308 35348 15360
rect 35400 15308 35406 15360
rect 36446 15308 36452 15360
rect 36504 15348 36510 15360
rect 37093 15351 37151 15357
rect 37093 15348 37105 15351
rect 36504 15320 37105 15348
rect 36504 15308 36510 15320
rect 37093 15317 37105 15320
rect 37139 15317 37151 15351
rect 37093 15311 37151 15317
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 9674 15104 9680 15156
rect 9732 15104 9738 15156
rect 9766 15104 9772 15156
rect 9824 15104 9830 15156
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11848 15116 11897 15144
rect 11848 15104 11854 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12342 15144 12348 15156
rect 12032 15116 12348 15144
rect 12032 15104 12038 15116
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 12952 15116 13369 15144
rect 12952 15104 12958 15116
rect 13357 15113 13369 15116
rect 13403 15144 13415 15147
rect 13906 15144 13912 15156
rect 13403 15116 13912 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 13906 15104 13912 15116
rect 13964 15144 13970 15156
rect 13964 15116 14504 15144
rect 13964 15104 13970 15116
rect 10870 15036 10876 15088
rect 10928 15036 10934 15088
rect 10962 15036 10968 15088
rect 11020 15076 11026 15088
rect 11057 15079 11115 15085
rect 11057 15076 11069 15079
rect 11020 15048 11069 15076
rect 11020 15036 11026 15048
rect 11057 15045 11069 15048
rect 11103 15076 11115 15079
rect 11606 15076 11612 15088
rect 11103 15048 11612 15076
rect 11103 15045 11115 15048
rect 11057 15039 11115 15045
rect 11606 15036 11612 15048
rect 11664 15036 11670 15088
rect 13446 15076 13452 15088
rect 12360 15048 13452 15076
rect 934 14968 940 15020
rect 992 15008 998 15020
rect 1765 15011 1823 15017
rect 1765 15008 1777 15011
rect 992 14980 1777 15008
rect 992 14968 998 14980
rect 1765 14977 1777 14980
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 4706 15008 4712 15020
rect 3007 14980 4712 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 10594 14968 10600 15020
rect 10652 15008 10658 15020
rect 12360 15017 12388 15048
rect 13446 15036 13452 15048
rect 13504 15036 13510 15088
rect 14274 15036 14280 15088
rect 14332 15036 14338 15088
rect 14476 15076 14504 15116
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 14608 15116 15577 15144
rect 14608 15104 14614 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 15933 15147 15991 15153
rect 15933 15113 15945 15147
rect 15979 15144 15991 15147
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 15979 15116 18337 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15144 18751 15147
rect 18739 15116 19334 15144
rect 18739 15113 18751 15116
rect 18693 15107 18751 15113
rect 14734 15076 14740 15088
rect 14476 15048 14740 15076
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 16022 15076 16028 15088
rect 15120 15048 16028 15076
rect 15120 15017 15148 15048
rect 16022 15036 16028 15048
rect 16080 15036 16086 15088
rect 19306 15076 19334 15116
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 19484 15116 19533 15144
rect 19484 15104 19490 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 19521 15107 19579 15113
rect 21450 15104 21456 15156
rect 21508 15144 21514 15156
rect 22005 15147 22063 15153
rect 22005 15144 22017 15147
rect 21508 15116 22017 15144
rect 21508 15104 21514 15116
rect 22005 15113 22017 15116
rect 22051 15113 22063 15147
rect 22005 15107 22063 15113
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23808 15116 24133 15144
rect 23808 15104 23814 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 24121 15107 24179 15113
rect 24762 15104 24768 15156
rect 24820 15144 24826 15156
rect 27065 15147 27123 15153
rect 24820 15116 26464 15144
rect 24820 15104 24826 15116
rect 19889 15079 19947 15085
rect 17144 15048 18828 15076
rect 19306 15048 19564 15076
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 10652 14980 12265 15008
rect 10652 14968 10658 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 14977 15163 15011
rect 17144 15008 17172 15048
rect 15105 14971 15163 14977
rect 15580 14980 17172 15008
rect 17221 15011 17279 15017
rect 9585 14943 9643 14949
rect 9585 14909 9597 14943
rect 9631 14940 9643 14943
rect 9766 14940 9772 14952
rect 9631 14912 9772 14940
rect 9631 14909 9643 14912
rect 9585 14903 9643 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12360 14940 12388 14971
rect 11655 14912 12388 14940
rect 12437 14943 12495 14949
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 10137 14875 10195 14881
rect 10137 14841 10149 14875
rect 10183 14872 10195 14875
rect 11974 14872 11980 14884
rect 10183 14844 11980 14872
rect 10183 14841 10195 14844
rect 10137 14835 10195 14841
rect 11974 14832 11980 14844
rect 12032 14832 12038 14884
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 12452 14872 12480 14903
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 14826 14940 14832 14952
rect 14516 14912 14832 14940
rect 14516 14900 14522 14912
rect 14826 14900 14832 14912
rect 14884 14940 14890 14952
rect 15580 14940 15608 14980
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 18690 15008 18696 15020
rect 17267 14980 18696 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 18800 15008 18828 15048
rect 19536 15020 19564 15048
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20806 15076 20812 15088
rect 19935 15048 20812 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 21085 15079 21143 15085
rect 21085 15045 21097 15079
rect 21131 15076 21143 15079
rect 21174 15076 21180 15088
rect 21131 15048 21180 15076
rect 21131 15045 21143 15048
rect 21085 15039 21143 15045
rect 21174 15036 21180 15048
rect 21232 15076 21238 15088
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 21232 15048 21833 15076
rect 21232 15036 21238 15048
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 21821 15039 21879 15045
rect 23385 15079 23443 15085
rect 23385 15045 23397 15079
rect 23431 15076 23443 15079
rect 25866 15076 25872 15088
rect 23431 15048 25872 15076
rect 23431 15045 23443 15048
rect 23385 15039 23443 15045
rect 25866 15036 25872 15048
rect 25924 15036 25930 15088
rect 18800 14980 18920 15008
rect 14884 14912 15608 14940
rect 14884 14900 14890 14912
rect 15654 14900 15660 14952
rect 15712 14940 15718 14952
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15712 14912 16037 14940
rect 15712 14900 15718 14912
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 12124 14844 12480 14872
rect 12124 14832 12130 14844
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 16132 14872 16160 14903
rect 16942 14900 16948 14952
rect 17000 14940 17006 14952
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 17000 14912 17325 14940
rect 17000 14900 17006 14912
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14909 17463 14943
rect 17405 14903 17463 14909
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 18782 14940 18788 14952
rect 18095 14912 18788 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 15436 14844 16160 14872
rect 15436 14832 15442 14844
rect 16298 14832 16304 14884
rect 16356 14872 16362 14884
rect 16356 14844 16988 14872
rect 16356 14832 16362 14844
rect 10594 14764 10600 14816
rect 10652 14764 10658 14816
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 12989 14807 13047 14813
rect 12989 14804 13001 14807
rect 12584 14776 13001 14804
rect 12584 14764 12590 14776
rect 12989 14773 13001 14776
rect 13035 14804 13047 14807
rect 14274 14804 14280 14816
rect 13035 14776 14280 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15396 14804 15424 14832
rect 14792 14776 15424 14804
rect 14792 14764 14798 14776
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 15988 14776 16865 14804
rect 15988 14764 15994 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16960 14804 16988 14844
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 17420 14872 17448 14903
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 18892 14949 18920 14980
rect 19518 14968 19524 15020
rect 19576 14968 19582 15020
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20898 15008 20904 15020
rect 20027 14980 20904 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 23290 14968 23296 15020
rect 23348 14968 23354 15020
rect 23934 15008 23940 15020
rect 23400 14980 23940 15008
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 20530 14940 20536 14952
rect 20211 14912 20536 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 20680 14912 21189 14940
rect 20680 14900 20686 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21266 14900 21272 14952
rect 21324 14900 21330 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 23400 14940 23428 14980
rect 23934 14968 23940 14980
rect 23992 14968 23998 15020
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 15008 24547 15011
rect 24946 15008 24952 15020
rect 24535 14980 24952 15008
rect 24535 14977 24547 14980
rect 24489 14971 24547 14977
rect 24946 14968 24952 14980
rect 25004 14968 25010 15020
rect 25222 14968 25228 15020
rect 25280 15008 25286 15020
rect 25317 15011 25375 15017
rect 25317 15008 25329 15011
rect 25280 14980 25329 15008
rect 25280 14968 25286 14980
rect 25317 14977 25329 14980
rect 25363 14977 25375 15011
rect 25317 14971 25375 14977
rect 25593 15011 25651 15017
rect 25593 14977 25605 15011
rect 25639 15008 25651 15011
rect 25958 15008 25964 15020
rect 25639 14980 25964 15008
rect 25639 14977 25651 14980
rect 25593 14971 25651 14977
rect 25958 14968 25964 14980
rect 26016 14968 26022 15020
rect 26234 14968 26240 15020
rect 26292 14968 26298 15020
rect 21968 14912 23428 14940
rect 21968 14900 21974 14912
rect 23566 14900 23572 14952
rect 23624 14900 23630 14952
rect 24578 14900 24584 14952
rect 24636 14900 24642 14952
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 24854 14900 24860 14952
rect 24912 14940 24918 14952
rect 26252 14940 26280 14968
rect 26436 14949 26464 15116
rect 27065 15113 27077 15147
rect 27111 15144 27123 15147
rect 27246 15144 27252 15156
rect 27111 15116 27252 15144
rect 27111 15113 27123 15116
rect 27065 15107 27123 15113
rect 27246 15104 27252 15116
rect 27304 15104 27310 15156
rect 27522 15104 27528 15156
rect 27580 15104 27586 15156
rect 28442 15104 28448 15156
rect 28500 15144 28506 15156
rect 29733 15147 29791 15153
rect 28500 15116 29684 15144
rect 28500 15104 28506 15116
rect 29656 15076 29684 15116
rect 29733 15113 29745 15147
rect 29779 15144 29791 15147
rect 29822 15144 29828 15156
rect 29779 15116 29828 15144
rect 29779 15113 29791 15116
rect 29733 15107 29791 15113
rect 29822 15104 29828 15116
rect 29880 15104 29886 15156
rect 30561 15147 30619 15153
rect 30561 15113 30573 15147
rect 30607 15144 30619 15147
rect 30650 15144 30656 15156
rect 30607 15116 30656 15144
rect 30607 15113 30619 15116
rect 30561 15107 30619 15113
rect 30650 15104 30656 15116
rect 30708 15104 30714 15156
rect 31294 15104 31300 15156
rect 31352 15144 31358 15156
rect 31389 15147 31447 15153
rect 31389 15144 31401 15147
rect 31352 15116 31401 15144
rect 31352 15104 31358 15116
rect 31389 15113 31401 15116
rect 31435 15113 31447 15147
rect 31389 15107 31447 15113
rect 32030 15104 32036 15156
rect 32088 15144 32094 15156
rect 33778 15144 33784 15156
rect 32088 15116 33784 15144
rect 32088 15104 32094 15116
rect 33778 15104 33784 15116
rect 33836 15104 33842 15156
rect 33870 15104 33876 15156
rect 33928 15104 33934 15156
rect 35069 15147 35127 15153
rect 35069 15113 35081 15147
rect 35115 15144 35127 15147
rect 35618 15144 35624 15156
rect 35115 15116 35624 15144
rect 35115 15113 35127 15116
rect 35069 15107 35127 15113
rect 35618 15104 35624 15116
rect 35676 15104 35682 15156
rect 36078 15104 36084 15156
rect 36136 15144 36142 15156
rect 36265 15147 36323 15153
rect 36265 15144 36277 15147
rect 36136 15116 36277 15144
rect 36136 15104 36142 15116
rect 36265 15113 36277 15116
rect 36311 15113 36323 15147
rect 36265 15107 36323 15113
rect 38654 15104 38660 15156
rect 38712 15144 38718 15156
rect 40129 15147 40187 15153
rect 40129 15144 40141 15147
rect 38712 15116 40141 15144
rect 38712 15104 38718 15116
rect 40129 15113 40141 15116
rect 40175 15113 40187 15147
rect 40129 15107 40187 15113
rect 29656 15048 31432 15076
rect 27246 14968 27252 15020
rect 27304 14968 27310 15020
rect 27798 14968 27804 15020
rect 27856 15008 27862 15020
rect 27985 15011 28043 15017
rect 27985 15008 27997 15011
rect 27856 14980 27997 15008
rect 27856 14968 27862 14980
rect 27985 14977 27997 14980
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 29362 14968 29368 15020
rect 29420 14968 29426 15020
rect 29546 14968 29552 15020
rect 29604 15008 29610 15020
rect 29604 14980 30788 15008
rect 29604 14968 29610 14980
rect 24912 14912 26280 14940
rect 26329 14943 26387 14949
rect 24912 14900 24918 14912
rect 26329 14909 26341 14943
rect 26375 14909 26387 14943
rect 26329 14903 26387 14909
rect 26421 14943 26479 14949
rect 26421 14909 26433 14943
rect 26467 14909 26479 14943
rect 26421 14903 26479 14909
rect 17276 14844 17448 14872
rect 17276 14832 17282 14844
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 17552 14844 20729 14872
rect 17552 14832 17558 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 20717 14835 20775 14841
rect 21082 14832 21088 14884
rect 21140 14872 21146 14884
rect 21450 14872 21456 14884
rect 21140 14844 21456 14872
rect 21140 14832 21146 14844
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 22830 14832 22836 14884
rect 22888 14872 22894 14884
rect 22925 14875 22983 14881
rect 22925 14872 22937 14875
rect 22888 14844 22937 14872
rect 22888 14832 22894 14844
rect 22925 14841 22937 14844
rect 22971 14841 22983 14875
rect 25869 14875 25927 14881
rect 25869 14872 25881 14875
rect 22925 14835 22983 14841
rect 24780 14844 25881 14872
rect 22370 14804 22376 14816
rect 16960 14776 22376 14804
rect 16853 14767 16911 14773
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 22646 14764 22652 14816
rect 22704 14804 22710 14816
rect 24780 14804 24808 14844
rect 25869 14841 25881 14844
rect 25915 14841 25927 14875
rect 26344 14872 26372 14903
rect 27154 14900 27160 14952
rect 27212 14940 27218 14952
rect 28261 14943 28319 14949
rect 28261 14940 28273 14943
rect 27212 14912 28273 14940
rect 27212 14900 27218 14912
rect 28261 14909 28273 14912
rect 28307 14940 28319 14943
rect 30282 14940 30288 14952
rect 28307 14912 30288 14940
rect 28307 14909 28319 14912
rect 28261 14903 28319 14909
rect 30282 14900 30288 14912
rect 30340 14900 30346 14952
rect 30374 14900 30380 14952
rect 30432 14940 30438 14952
rect 30760 14949 30788 14980
rect 30653 14943 30711 14949
rect 30653 14940 30665 14943
rect 30432 14912 30665 14940
rect 30432 14900 30438 14912
rect 30653 14909 30665 14912
rect 30699 14909 30711 14943
rect 30653 14903 30711 14909
rect 30745 14943 30803 14949
rect 30745 14909 30757 14943
rect 30791 14909 30803 14943
rect 31404 14940 31432 15048
rect 32306 15036 32312 15088
rect 32364 15076 32370 15088
rect 32364 15048 32904 15076
rect 32364 15036 32370 15048
rect 31754 14968 31760 15020
rect 31812 15008 31818 15020
rect 32677 15011 32735 15017
rect 32677 15008 32689 15011
rect 31812 14980 32689 15008
rect 31812 14968 31818 14980
rect 32677 14977 32689 14980
rect 32723 14977 32735 15011
rect 32677 14971 32735 14977
rect 32876 14949 32904 15048
rect 34238 15036 34244 15088
rect 34296 15076 34302 15088
rect 34882 15076 34888 15088
rect 34296 15048 34888 15076
rect 34296 15036 34302 15048
rect 34882 15036 34888 15048
rect 34940 15036 34946 15088
rect 35802 15036 35808 15088
rect 35860 15076 35866 15088
rect 36173 15079 36231 15085
rect 36173 15076 36185 15079
rect 35860 15048 36185 15076
rect 35860 15036 35866 15048
rect 36173 15045 36185 15048
rect 36219 15045 36231 15079
rect 36173 15039 36231 15045
rect 36354 15036 36360 15088
rect 36412 15076 36418 15088
rect 37642 15076 37648 15088
rect 36412 15048 37648 15076
rect 36412 15036 36418 15048
rect 37642 15036 37648 15048
rect 37700 15036 37706 15088
rect 37734 15036 37740 15088
rect 37792 15036 37798 15088
rect 38746 15036 38752 15088
rect 38804 15036 38810 15088
rect 40037 15079 40095 15085
rect 40037 15045 40049 15079
rect 40083 15076 40095 15079
rect 48406 15076 48412 15088
rect 40083 15048 48412 15076
rect 40083 15045 40095 15048
rect 40037 15039 40095 15045
rect 48406 15036 48412 15048
rect 48464 15036 48470 15088
rect 33962 15008 33968 15020
rect 33704 14980 33968 15008
rect 33704 14949 33732 14980
rect 33962 14968 33968 14980
rect 34020 14968 34026 15020
rect 34900 14980 37320 15008
rect 32769 14943 32827 14949
rect 31404 14912 31754 14940
rect 30745 14903 30803 14909
rect 27433 14875 27491 14881
rect 27433 14872 27445 14875
rect 26344 14844 27445 14872
rect 25869 14835 25927 14841
rect 27433 14841 27445 14844
rect 27479 14872 27491 14875
rect 31478 14872 31484 14884
rect 27479 14844 28120 14872
rect 27479 14841 27491 14844
rect 27433 14835 27491 14841
rect 22704 14776 24808 14804
rect 22704 14764 22710 14776
rect 24946 14764 24952 14816
rect 25004 14804 25010 14816
rect 25133 14807 25191 14813
rect 25133 14804 25145 14807
rect 25004 14776 25145 14804
rect 25004 14764 25010 14776
rect 25133 14773 25145 14776
rect 25179 14773 25191 14807
rect 25133 14767 25191 14773
rect 25406 14764 25412 14816
rect 25464 14804 25470 14816
rect 27982 14804 27988 14816
rect 25464 14776 27988 14804
rect 25464 14764 25470 14776
rect 27982 14764 27988 14776
rect 28040 14764 28046 14816
rect 28092 14804 28120 14844
rect 29288 14844 31484 14872
rect 29288 14804 29316 14844
rect 31478 14832 31484 14844
rect 31536 14832 31542 14884
rect 31726 14872 31754 14912
rect 32769 14909 32781 14943
rect 32815 14909 32827 14943
rect 32769 14903 32827 14909
rect 32861 14943 32919 14949
rect 32861 14909 32873 14943
rect 32907 14909 32919 14943
rect 32861 14903 32919 14909
rect 33689 14943 33747 14949
rect 33689 14909 33701 14943
rect 33735 14909 33747 14943
rect 33689 14903 33747 14909
rect 32309 14875 32367 14881
rect 32309 14872 32321 14875
rect 31726 14844 32321 14872
rect 32309 14841 32321 14844
rect 32355 14841 32367 14875
rect 32784 14872 32812 14903
rect 33778 14900 33784 14952
rect 33836 14900 33842 14952
rect 34900 14949 34928 14980
rect 34885 14943 34943 14949
rect 34885 14909 34897 14943
rect 34931 14909 34943 14943
rect 34885 14903 34943 14909
rect 34977 14943 35035 14949
rect 34977 14909 34989 14943
rect 35023 14940 35035 14943
rect 35894 14940 35900 14952
rect 35023 14912 35900 14940
rect 35023 14909 35035 14912
rect 34977 14903 35035 14909
rect 35894 14900 35900 14912
rect 35952 14900 35958 14952
rect 35986 14900 35992 14952
rect 36044 14900 36050 14952
rect 36078 14900 36084 14952
rect 36136 14940 36142 14952
rect 37001 14943 37059 14949
rect 37001 14940 37013 14943
rect 36136 14912 37013 14940
rect 36136 14900 36142 14912
rect 37001 14909 37013 14912
rect 37047 14940 37059 14943
rect 37090 14940 37096 14952
rect 37047 14912 37096 14940
rect 37047 14909 37059 14912
rect 37001 14903 37059 14909
rect 37090 14900 37096 14912
rect 37148 14900 37154 14952
rect 37292 14940 37320 14980
rect 37366 14968 37372 15020
rect 37424 15008 37430 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 37424 14980 37473 15008
rect 37424 14968 37430 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 40862 14968 40868 15020
rect 40920 14968 40926 15020
rect 48777 15011 48835 15017
rect 48777 14977 48789 15011
rect 48823 15008 48835 15011
rect 49326 15008 49332 15020
rect 48823 14980 49332 15008
rect 48823 14977 48835 14980
rect 48777 14971 48835 14977
rect 49326 14968 49332 14980
rect 49384 14968 49390 15020
rect 37826 14940 37832 14952
rect 37292 14912 37832 14940
rect 37826 14900 37832 14912
rect 37884 14900 37890 14952
rect 38286 14900 38292 14952
rect 38344 14940 38350 14952
rect 39209 14943 39267 14949
rect 39209 14940 39221 14943
rect 38344 14912 39221 14940
rect 38344 14900 38350 14912
rect 39209 14909 39221 14912
rect 39255 14909 39267 14943
rect 39209 14903 39267 14909
rect 39390 14900 39396 14952
rect 39448 14940 39454 14952
rect 40221 14943 40279 14949
rect 40221 14940 40233 14943
rect 39448 14912 40233 14940
rect 39448 14900 39454 14912
rect 40221 14909 40233 14912
rect 40267 14909 40279 14943
rect 40221 14903 40279 14909
rect 39669 14875 39727 14881
rect 39669 14872 39681 14875
rect 32784 14844 37044 14872
rect 32309 14835 32367 14841
rect 28092 14776 29316 14804
rect 30190 14764 30196 14816
rect 30248 14764 30254 14816
rect 30374 14764 30380 14816
rect 30432 14804 30438 14816
rect 31849 14807 31907 14813
rect 31849 14804 31861 14807
rect 30432 14776 31861 14804
rect 30432 14764 30438 14776
rect 31849 14773 31861 14776
rect 31895 14773 31907 14807
rect 31849 14767 31907 14773
rect 34238 14764 34244 14816
rect 34296 14764 34302 14816
rect 35437 14807 35495 14813
rect 35437 14773 35449 14807
rect 35483 14804 35495 14807
rect 36354 14804 36360 14816
rect 35483 14776 36360 14804
rect 35483 14773 35495 14776
rect 35437 14767 35495 14773
rect 36354 14764 36360 14776
rect 36412 14764 36418 14816
rect 36633 14807 36691 14813
rect 36633 14773 36645 14807
rect 36679 14804 36691 14807
rect 36814 14804 36820 14816
rect 36679 14776 36820 14804
rect 36679 14773 36691 14776
rect 36633 14767 36691 14773
rect 36814 14764 36820 14776
rect 36872 14764 36878 14816
rect 37016 14804 37044 14844
rect 38764 14844 39681 14872
rect 38764 14804 38792 14844
rect 39669 14841 39681 14844
rect 39715 14841 39727 14875
rect 39669 14835 39727 14841
rect 49142 14832 49148 14884
rect 49200 14832 49206 14884
rect 37016 14776 38792 14804
rect 41049 14807 41107 14813
rect 41049 14773 41061 14807
rect 41095 14804 41107 14807
rect 45646 14804 45652 14816
rect 41095 14776 45652 14804
rect 41095 14773 41107 14776
rect 41049 14767 41107 14773
rect 45646 14764 45652 14776
rect 45704 14764 45710 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11296 14572 11805 14600
rect 11296 14560 11302 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12860 14572 13001 14600
rect 12860 14560 12866 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 13998 14600 14004 14612
rect 12989 14563 13047 14569
rect 13372 14572 14004 14600
rect 10226 14492 10232 14544
rect 10284 14492 10290 14544
rect 13372 14532 13400 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14182 14560 14188 14612
rect 14240 14560 14246 14612
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 14642 14600 14648 14612
rect 14507 14572 14648 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 18141 14603 18199 14609
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18414 14600 18420 14612
rect 18187 14572 18420 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 19306 14572 23060 14600
rect 10612 14504 13400 14532
rect 934 14424 940 14476
rect 992 14464 998 14476
rect 1765 14467 1823 14473
rect 1765 14464 1777 14467
rect 992 14436 1777 14464
rect 992 14424 998 14436
rect 1765 14433 1777 14436
rect 1811 14433 1823 14467
rect 1765 14427 1823 14433
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 3007 14368 9505 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 9950 14396 9956 14408
rect 9723 14368 9956 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 9950 14356 9956 14368
rect 10008 14396 10014 14408
rect 10612 14396 10640 14504
rect 13446 14492 13452 14544
rect 13504 14532 13510 14544
rect 19306 14532 19334 14572
rect 13504 14504 19334 14532
rect 22388 14504 22692 14532
rect 13504 14492 13510 14504
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 13262 14464 13268 14476
rect 12483 14436 13268 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 13412 14436 13553 14464
rect 13412 14424 13418 14436
rect 13541 14433 13553 14436
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 13630 14424 13636 14476
rect 13688 14464 13694 14476
rect 14826 14464 14832 14476
rect 13688 14436 14832 14464
rect 13688 14424 13694 14436
rect 14826 14424 14832 14436
rect 14884 14424 14890 14476
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 10008 14368 10640 14396
rect 10008 14356 10014 14368
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14921 14399 14979 14405
rect 14921 14396 14933 14399
rect 13872 14368 14933 14396
rect 13872 14356 13878 14368
rect 14921 14365 14933 14368
rect 14967 14365 14979 14399
rect 14921 14359 14979 14365
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15120 14396 15148 14427
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 15436 14436 16957 14464
rect 15436 14424 15442 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17497 14467 17555 14473
rect 17497 14433 17509 14467
rect 17543 14464 17555 14467
rect 18693 14467 18751 14473
rect 18693 14464 18705 14467
rect 17543 14436 18705 14464
rect 17543 14433 17555 14436
rect 17497 14427 17555 14433
rect 18693 14433 18705 14436
rect 18739 14433 18751 14467
rect 18693 14427 18751 14433
rect 17402 14396 17408 14408
rect 15068 14368 17408 14396
rect 15068 14356 15074 14368
rect 17402 14356 17408 14368
rect 17460 14396 17466 14408
rect 17512 14396 17540 14427
rect 20070 14424 20076 14476
rect 20128 14424 20134 14476
rect 21082 14424 21088 14476
rect 21140 14424 21146 14476
rect 21358 14424 21364 14476
rect 21416 14424 21422 14476
rect 21450 14424 21456 14476
rect 21508 14464 21514 14476
rect 22388 14464 22416 14504
rect 21508 14436 22416 14464
rect 22664 14464 22692 14504
rect 22738 14492 22744 14544
rect 22796 14532 22802 14544
rect 22833 14535 22891 14541
rect 22833 14532 22845 14535
rect 22796 14504 22845 14532
rect 22796 14492 22802 14504
rect 22833 14501 22845 14504
rect 22879 14501 22891 14535
rect 23032 14532 23060 14572
rect 23106 14560 23112 14612
rect 23164 14600 23170 14612
rect 24578 14600 24584 14612
rect 23164 14572 24584 14600
rect 23164 14560 23170 14572
rect 24578 14560 24584 14572
rect 24636 14600 24642 14612
rect 24854 14600 24860 14612
rect 24636 14572 24860 14600
rect 24636 14560 24642 14572
rect 24854 14560 24860 14572
rect 24912 14560 24918 14612
rect 25498 14560 25504 14612
rect 25556 14600 25562 14612
rect 25593 14603 25651 14609
rect 25593 14600 25605 14603
rect 25556 14572 25605 14600
rect 25556 14560 25562 14572
rect 25593 14569 25605 14572
rect 25639 14569 25651 14603
rect 26326 14600 26332 14612
rect 25593 14563 25651 14569
rect 25700 14572 26332 14600
rect 25700 14532 25728 14572
rect 26326 14560 26332 14572
rect 26384 14560 26390 14612
rect 26510 14560 26516 14612
rect 26568 14600 26574 14612
rect 30374 14600 30380 14612
rect 26568 14572 30380 14600
rect 26568 14560 26574 14572
rect 30374 14560 30380 14572
rect 30432 14560 30438 14612
rect 30469 14603 30527 14609
rect 30469 14569 30481 14603
rect 30515 14600 30527 14603
rect 33778 14600 33784 14612
rect 30515 14572 33784 14600
rect 30515 14569 30527 14572
rect 30469 14563 30527 14569
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 34238 14560 34244 14612
rect 34296 14600 34302 14612
rect 34296 14572 36216 14600
rect 34296 14560 34302 14572
rect 29270 14532 29276 14544
rect 23032 14504 25728 14532
rect 27264 14504 29276 14532
rect 22833 14495 22891 14501
rect 27264 14464 27292 14504
rect 29270 14492 29276 14504
rect 29328 14532 29334 14544
rect 29730 14532 29736 14544
rect 29328 14504 29736 14532
rect 29328 14492 29334 14504
rect 29730 14492 29736 14504
rect 29788 14492 29794 14544
rect 31665 14535 31723 14541
rect 31665 14501 31677 14535
rect 31711 14532 31723 14535
rect 33318 14532 33324 14544
rect 31711 14504 33324 14532
rect 31711 14501 31723 14504
rect 31665 14495 31723 14501
rect 33318 14492 33324 14504
rect 33376 14492 33382 14544
rect 33502 14492 33508 14544
rect 33560 14492 33566 14544
rect 34057 14535 34115 14541
rect 34057 14501 34069 14535
rect 34103 14532 34115 14535
rect 36188 14532 36216 14572
rect 36354 14560 36360 14612
rect 36412 14600 36418 14612
rect 36633 14603 36691 14609
rect 36633 14600 36645 14603
rect 36412 14572 36645 14600
rect 36412 14560 36418 14572
rect 36633 14569 36645 14572
rect 36679 14569 36691 14603
rect 36633 14563 36691 14569
rect 36814 14560 36820 14612
rect 36872 14600 36878 14612
rect 38746 14600 38752 14612
rect 36872 14572 38752 14600
rect 36872 14560 36878 14572
rect 38746 14560 38752 14572
rect 38804 14560 38810 14612
rect 39942 14560 39948 14612
rect 40000 14600 40006 14612
rect 40037 14603 40095 14609
rect 40037 14600 40049 14603
rect 40000 14572 40049 14600
rect 40000 14560 40006 14572
rect 40037 14569 40049 14572
rect 40083 14569 40095 14603
rect 40037 14563 40095 14569
rect 37550 14532 37556 14544
rect 34103 14504 35020 14532
rect 36188 14504 37556 14532
rect 34103 14501 34115 14504
rect 34057 14495 34115 14501
rect 22664 14436 27292 14464
rect 21508 14424 21514 14436
rect 27890 14424 27896 14476
rect 27948 14464 27954 14476
rect 27985 14467 28043 14473
rect 27985 14464 27997 14467
rect 27948 14436 27997 14464
rect 27948 14424 27954 14436
rect 27985 14433 27997 14436
rect 28031 14464 28043 14467
rect 28718 14464 28724 14476
rect 28031 14436 28724 14464
rect 28031 14433 28043 14436
rect 27985 14427 28043 14433
rect 28718 14424 28724 14436
rect 28776 14424 28782 14476
rect 29917 14467 29975 14473
rect 29917 14433 29929 14467
rect 29963 14464 29975 14467
rect 30558 14464 30564 14476
rect 29963 14436 30564 14464
rect 29963 14433 29975 14436
rect 29917 14427 29975 14433
rect 30558 14424 30564 14436
rect 30616 14424 30622 14476
rect 30742 14424 30748 14476
rect 30800 14464 30806 14476
rect 31021 14467 31079 14473
rect 31021 14464 31033 14467
rect 30800 14436 31033 14464
rect 30800 14424 30806 14436
rect 31021 14433 31033 14436
rect 31067 14433 31079 14467
rect 31021 14427 31079 14433
rect 32309 14467 32367 14473
rect 32309 14433 32321 14467
rect 32355 14464 32367 14467
rect 32398 14464 32404 14476
rect 32355 14436 32404 14464
rect 32355 14433 32367 14436
rect 32309 14427 32367 14433
rect 32398 14424 32404 14436
rect 32456 14424 32462 14476
rect 32582 14424 32588 14476
rect 32640 14464 32646 14476
rect 33413 14467 33471 14473
rect 33413 14464 33425 14467
rect 32640 14436 33425 14464
rect 32640 14424 32646 14436
rect 33413 14433 33425 14436
rect 33459 14433 33471 14467
rect 33520 14464 33548 14492
rect 34333 14467 34391 14473
rect 34333 14464 34345 14467
rect 33520 14436 34345 14464
rect 33413 14427 33471 14433
rect 34333 14433 34345 14436
rect 34379 14433 34391 14467
rect 34333 14427 34391 14433
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 34885 14467 34943 14473
rect 34885 14464 34897 14467
rect 34848 14436 34897 14464
rect 34848 14424 34854 14436
rect 34885 14433 34897 14436
rect 34931 14433 34943 14467
rect 34992 14464 35020 14504
rect 37550 14492 37556 14504
rect 37608 14492 37614 14544
rect 49050 14492 49056 14544
rect 49108 14492 49114 14544
rect 37274 14464 37280 14476
rect 34992 14436 37280 14464
rect 34885 14427 34943 14433
rect 37274 14424 37280 14436
rect 37332 14424 37338 14476
rect 37366 14424 37372 14476
rect 37424 14464 37430 14476
rect 38841 14467 38899 14473
rect 38841 14464 38853 14467
rect 37424 14436 38853 14464
rect 37424 14424 37430 14436
rect 38841 14433 38853 14436
rect 38887 14433 38899 14467
rect 38841 14427 38899 14433
rect 17460 14368 17540 14396
rect 17460 14356 17466 14368
rect 17678 14356 17684 14408
rect 17736 14396 17742 14408
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 17736 14368 18613 14396
rect 17736 14356 17742 14368
rect 18601 14365 18613 14368
rect 18647 14396 18659 14399
rect 19334 14396 19340 14408
rect 18647 14368 19340 14396
rect 18647 14365 18659 14368
rect 18601 14359 18659 14365
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19886 14356 19892 14408
rect 19944 14356 19950 14408
rect 27341 14399 27399 14405
rect 27341 14365 27353 14399
rect 27387 14396 27399 14399
rect 27614 14396 27620 14408
rect 27387 14368 27620 14396
rect 27387 14365 27399 14368
rect 27341 14359 27399 14365
rect 27614 14356 27620 14368
rect 27672 14396 27678 14408
rect 30006 14396 30012 14408
rect 27672 14368 30012 14396
rect 27672 14356 27678 14368
rect 30006 14356 30012 14368
rect 30064 14356 30070 14408
rect 30098 14356 30104 14408
rect 30156 14356 30162 14408
rect 30834 14356 30840 14408
rect 30892 14396 30898 14408
rect 31297 14399 31355 14405
rect 31297 14396 31309 14399
rect 30892 14368 31309 14396
rect 30892 14356 30898 14368
rect 31297 14365 31309 14368
rect 31343 14365 31355 14399
rect 31297 14359 31355 14365
rect 32858 14356 32864 14408
rect 32916 14396 32922 14408
rect 33597 14399 33655 14405
rect 33597 14396 33609 14399
rect 32916 14368 33609 14396
rect 32916 14356 32922 14368
rect 33597 14365 33609 14368
rect 33643 14365 33655 14399
rect 33597 14359 33655 14365
rect 33686 14356 33692 14408
rect 33744 14356 33750 14408
rect 39298 14356 39304 14408
rect 39356 14356 39362 14408
rect 48593 14399 48651 14405
rect 48593 14365 48605 14399
rect 48639 14396 48651 14399
rect 49234 14396 49240 14408
rect 48639 14368 49240 14396
rect 48639 14365 48651 14368
rect 48593 14359 48651 14365
rect 49234 14356 49240 14368
rect 49292 14356 49298 14408
rect 10410 14288 10416 14340
rect 10468 14288 10474 14340
rect 11238 14288 11244 14340
rect 11296 14288 11302 14340
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12802 14328 12808 14340
rect 12207 14300 12808 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 12802 14288 12808 14300
rect 12860 14288 12866 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 15933 14331 15991 14337
rect 13403 14300 15056 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10560 14232 11161 14260
rect 10560 14220 10566 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 12618 14260 12624 14272
rect 12299 14232 12624 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 13906 14260 13912 14272
rect 13495 14232 13912 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13906 14220 13912 14232
rect 13964 14220 13970 14272
rect 14826 14220 14832 14272
rect 14884 14220 14890 14272
rect 15028 14260 15056 14300
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16761 14331 16819 14337
rect 16761 14328 16773 14331
rect 15979 14300 16773 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16761 14297 16773 14300
rect 16807 14297 16819 14331
rect 17865 14331 17923 14337
rect 16761 14291 16819 14297
rect 16868 14300 17816 14328
rect 16868 14272 16896 14300
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15028 14232 16405 14260
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 16850 14260 16856 14272
rect 16632 14232 16856 14260
rect 16632 14220 16638 14232
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 17218 14220 17224 14272
rect 17276 14260 17282 14272
rect 17589 14263 17647 14269
rect 17589 14260 17601 14263
rect 17276 14232 17601 14260
rect 17276 14220 17282 14232
rect 17589 14229 17601 14232
rect 17635 14229 17647 14263
rect 17788 14260 17816 14300
rect 17865 14297 17877 14331
rect 17911 14328 17923 14331
rect 19426 14328 19432 14340
rect 17911 14300 19432 14328
rect 17911 14297 17923 14300
rect 17865 14291 17923 14297
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 19978 14288 19984 14340
rect 20036 14328 20042 14340
rect 21450 14328 21456 14340
rect 20036 14300 21456 14328
rect 20036 14288 20042 14300
rect 21450 14288 21456 14300
rect 21508 14288 21514 14340
rect 21818 14328 21824 14340
rect 21560 14300 21824 14328
rect 21560 14272 21588 14300
rect 21818 14288 21824 14300
rect 21876 14288 21882 14340
rect 25774 14288 25780 14340
rect 25832 14328 25838 14340
rect 25832 14300 25898 14328
rect 25832 14288 25838 14300
rect 27062 14288 27068 14340
rect 27120 14288 27126 14340
rect 27706 14288 27712 14340
rect 27764 14328 27770 14340
rect 28169 14331 28227 14337
rect 28169 14328 28181 14331
rect 27764 14300 28181 14328
rect 27764 14288 27770 14300
rect 28169 14297 28181 14300
rect 28215 14297 28227 14331
rect 31205 14331 31263 14337
rect 31205 14328 31217 14331
rect 28169 14291 28227 14297
rect 28552 14300 31217 14328
rect 18414 14260 18420 14272
rect 17788 14232 18420 14260
rect 17589 14223 17647 14229
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 18966 14260 18972 14272
rect 18555 14232 18972 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 19518 14220 19524 14272
rect 19576 14220 19582 14272
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21542 14260 21548 14272
rect 20772 14232 21548 14260
rect 20772 14220 20778 14232
rect 21542 14220 21548 14232
rect 21600 14260 21606 14272
rect 23201 14263 23259 14269
rect 23201 14260 23213 14263
rect 21600 14232 23213 14260
rect 21600 14220 21606 14232
rect 23201 14229 23213 14232
rect 23247 14260 23259 14263
rect 23477 14263 23535 14269
rect 23477 14260 23489 14263
rect 23247 14232 23489 14260
rect 23247 14229 23259 14232
rect 23201 14223 23259 14229
rect 23477 14229 23489 14232
rect 23523 14229 23535 14263
rect 23477 14223 23535 14229
rect 23842 14220 23848 14272
rect 23900 14220 23906 14272
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 25130 14220 25136 14272
rect 25188 14220 25194 14272
rect 27522 14220 27528 14272
rect 27580 14260 27586 14272
rect 28077 14263 28135 14269
rect 28077 14260 28089 14263
rect 27580 14232 28089 14260
rect 27580 14220 27586 14232
rect 28077 14229 28089 14232
rect 28123 14260 28135 14263
rect 28442 14260 28448 14272
rect 28123 14232 28448 14260
rect 28123 14229 28135 14232
rect 28077 14223 28135 14229
rect 28442 14220 28448 14232
rect 28500 14220 28506 14272
rect 28552 14269 28580 14300
rect 31205 14297 31217 14300
rect 31251 14297 31263 14331
rect 31205 14291 31263 14297
rect 31478 14288 31484 14340
rect 31536 14328 31542 14340
rect 32030 14328 32036 14340
rect 31536 14300 32036 14328
rect 31536 14288 31542 14300
rect 32030 14288 32036 14300
rect 32088 14288 32094 14340
rect 32493 14331 32551 14337
rect 32493 14297 32505 14331
rect 32539 14328 32551 14331
rect 32539 14300 33732 14328
rect 32539 14297 32551 14300
rect 32493 14291 32551 14297
rect 33704 14272 33732 14300
rect 35158 14288 35164 14340
rect 35216 14288 35222 14340
rect 35434 14288 35440 14340
rect 35492 14328 35498 14340
rect 35492 14300 35650 14328
rect 35492 14288 35498 14300
rect 36630 14288 36636 14340
rect 36688 14328 36694 14340
rect 36688 14300 37398 14328
rect 36688 14288 36694 14300
rect 38286 14288 38292 14340
rect 38344 14328 38350 14340
rect 38565 14331 38623 14337
rect 38565 14328 38577 14331
rect 38344 14300 38577 14328
rect 38344 14288 38350 14300
rect 38565 14297 38577 14300
rect 38611 14297 38623 14331
rect 38565 14291 38623 14297
rect 28537 14263 28595 14269
rect 28537 14229 28549 14263
rect 28583 14229 28595 14263
rect 28537 14223 28595 14229
rect 28994 14220 29000 14272
rect 29052 14220 29058 14272
rect 29638 14220 29644 14272
rect 29696 14260 29702 14272
rect 30009 14263 30067 14269
rect 30009 14260 30021 14263
rect 29696 14232 30021 14260
rect 29696 14220 29702 14232
rect 30009 14229 30021 14232
rect 30055 14229 30067 14263
rect 30009 14223 30067 14229
rect 30374 14220 30380 14272
rect 30432 14260 30438 14272
rect 32401 14263 32459 14269
rect 32401 14260 32413 14263
rect 30432 14232 32413 14260
rect 30432 14220 30438 14232
rect 32401 14229 32413 14232
rect 32447 14229 32459 14263
rect 32401 14223 32459 14229
rect 32766 14220 32772 14272
rect 32824 14260 32830 14272
rect 32861 14263 32919 14269
rect 32861 14260 32873 14263
rect 32824 14232 32873 14260
rect 32824 14220 32830 14232
rect 32861 14229 32873 14232
rect 32907 14229 32919 14263
rect 32861 14223 32919 14229
rect 33686 14220 33692 14272
rect 33744 14220 33750 14272
rect 35176 14260 35204 14288
rect 35342 14260 35348 14272
rect 35176 14232 35348 14260
rect 35342 14220 35348 14232
rect 35400 14260 35406 14272
rect 35802 14260 35808 14272
rect 35400 14232 35808 14260
rect 35400 14220 35406 14232
rect 35802 14220 35808 14232
rect 35860 14220 35866 14272
rect 35894 14220 35900 14272
rect 35952 14260 35958 14272
rect 37093 14263 37151 14269
rect 37093 14260 37105 14263
rect 35952 14232 37105 14260
rect 35952 14220 35958 14232
rect 37093 14229 37105 14232
rect 37139 14260 37151 14263
rect 39390 14260 39396 14272
rect 37139 14232 39396 14260
rect 37139 14229 37151 14232
rect 37093 14223 37151 14229
rect 39390 14220 39396 14232
rect 39448 14220 39454 14272
rect 39482 14220 39488 14272
rect 39540 14220 39546 14272
rect 48314 14220 48320 14272
rect 48372 14260 48378 14272
rect 48685 14263 48743 14269
rect 48685 14260 48697 14263
rect 48372 14232 48697 14260
rect 48372 14220 48378 14232
rect 48685 14229 48697 14232
rect 48731 14229 48743 14263
rect 48685 14223 48743 14229
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 9950 14016 9956 14068
rect 10008 14016 10014 14068
rect 10410 14016 10416 14068
rect 10468 14016 10474 14068
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12342 14056 12348 14068
rect 12023 14028 12348 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 15013 14059 15071 14065
rect 15013 14056 15025 14059
rect 14332 14028 15025 14056
rect 14332 14016 14338 14028
rect 1026 13948 1032 14000
rect 1084 13988 1090 14000
rect 1765 13991 1823 13997
rect 1765 13988 1777 13991
rect 1084 13960 1777 13988
rect 1084 13948 1090 13960
rect 1765 13957 1777 13960
rect 1811 13957 1823 13991
rect 10502 13988 10508 14000
rect 1765 13951 1823 13957
rect 2976 13960 10508 13988
rect 2976 13929 3004 13960
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 10689 13991 10747 13997
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 11238 13988 11244 14000
rect 10735 13960 11244 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 13262 13948 13268 14000
rect 13320 13948 13326 14000
rect 14568 13988 14596 14028
rect 15013 14025 15025 14028
rect 15059 14025 15071 14059
rect 15013 14019 15071 14025
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 15252 14028 15577 14056
rect 15252 14016 15258 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 15930 14016 15936 14068
rect 15988 14016 15994 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 16632 14028 17141 14056
rect 16632 14016 16638 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17129 14019 17187 14025
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19058 14056 19064 14068
rect 18739 14028 19064 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 19886 14056 19892 14068
rect 19475 14028 19892 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21416 14028 21465 14056
rect 21416 14016 21422 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 24857 14059 24915 14065
rect 24857 14025 24869 14059
rect 24903 14056 24915 14059
rect 25314 14056 25320 14068
rect 24903 14028 25320 14056
rect 24903 14025 24915 14028
rect 24857 14019 24915 14025
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 27522 14056 27528 14068
rect 25556 14028 26004 14056
rect 25556 14016 25562 14028
rect 14734 13988 14740 14000
rect 14490 13960 14740 13988
rect 14734 13948 14740 13960
rect 14792 13948 14798 14000
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3568 13892 3985 13920
rect 3568 13880 3574 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11195 13892 12081 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 15838 13920 15844 13932
rect 12069 13883 12127 13889
rect 14752 13892 15844 13920
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13852 3755 13855
rect 10318 13852 10324 13864
rect 3743 13824 10324 13852
rect 3743 13821 3755 13824
rect 3697 13815 3755 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13821 11943 13855
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 11885 13815 11943 13821
rect 12406 13824 13001 13852
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 11900 13716 11928 13815
rect 12066 13744 12072 13796
rect 12124 13784 12130 13796
rect 12406 13784 12434 13824
rect 12989 13821 13001 13824
rect 13035 13852 13047 13855
rect 13630 13852 13636 13864
rect 13035 13824 13636 13852
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 14752 13861 14780 13892
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 15948 13929 15976 14016
rect 16025 13991 16083 13997
rect 16025 13957 16037 13991
rect 16071 13988 16083 13991
rect 19518 13988 19524 14000
rect 16071 13960 19524 13988
rect 16071 13957 16083 13960
rect 16025 13951 16083 13957
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 20622 13948 20628 14000
rect 20680 13948 20686 14000
rect 21818 13948 21824 14000
rect 21876 13988 21882 14000
rect 23477 13991 23535 13997
rect 21876 13960 22310 13988
rect 21876 13948 21882 13960
rect 23477 13957 23489 13991
rect 23523 13988 23535 13991
rect 24026 13988 24032 14000
rect 23523 13960 24032 13988
rect 23523 13957 23535 13960
rect 23477 13951 23535 13957
rect 24026 13948 24032 13960
rect 24084 13948 24090 14000
rect 25774 13948 25780 14000
rect 25832 13948 25838 14000
rect 25976 13988 26004 14028
rect 26620 14028 27528 14056
rect 26329 13991 26387 13997
rect 26329 13988 26341 13991
rect 25976 13960 26341 13988
rect 26329 13957 26341 13960
rect 26375 13957 26387 13991
rect 26329 13951 26387 13957
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16816 13892 16865 13920
rect 16816 13880 16822 13892
rect 16853 13889 16865 13892
rect 16899 13920 16911 13923
rect 17678 13920 17684 13932
rect 16899 13892 17684 13920
rect 16899 13889 16911 13892
rect 16853 13883 16911 13889
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18690 13920 18696 13932
rect 18472 13892 18696 13920
rect 18472 13880 18478 13892
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 19426 13920 19432 13932
rect 18831 13892 19432 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 26620 13929 26648 14028
rect 27522 14016 27528 14028
rect 27580 14016 27586 14068
rect 27617 14059 27675 14065
rect 27617 14025 27629 14059
rect 27663 14056 27675 14059
rect 28810 14056 28816 14068
rect 27663 14028 28816 14056
rect 27663 14025 27675 14028
rect 27617 14019 27675 14025
rect 28810 14016 28816 14028
rect 28868 14016 28874 14068
rect 30006 14016 30012 14068
rect 30064 14056 30070 14068
rect 31110 14056 31116 14068
rect 30064 14028 31116 14056
rect 30064 14016 30070 14028
rect 31110 14016 31116 14028
rect 31168 14016 31174 14068
rect 31757 14059 31815 14065
rect 31757 14025 31769 14059
rect 31803 14056 31815 14059
rect 31803 14028 33916 14056
rect 31803 14025 31815 14028
rect 31757 14019 31815 14025
rect 31846 13988 31852 14000
rect 30406 13960 31852 13988
rect 31846 13948 31852 13960
rect 31904 13948 31910 14000
rect 33318 13948 33324 14000
rect 33376 13948 33382 14000
rect 33888 13988 33916 14028
rect 34422 14016 34428 14068
rect 34480 14056 34486 14068
rect 34885 14059 34943 14065
rect 34885 14056 34897 14059
rect 34480 14028 34897 14056
rect 34480 14016 34486 14028
rect 34885 14025 34897 14028
rect 34931 14025 34943 14059
rect 34885 14019 34943 14025
rect 35253 14059 35311 14065
rect 35253 14025 35265 14059
rect 35299 14056 35311 14059
rect 35710 14056 35716 14068
rect 35299 14028 35716 14056
rect 35299 14025 35311 14028
rect 35253 14019 35311 14025
rect 35710 14016 35716 14028
rect 35768 14016 35774 14068
rect 35802 14016 35808 14068
rect 35860 14056 35866 14068
rect 36449 14059 36507 14065
rect 35860 14028 36216 14056
rect 35860 14016 35866 14028
rect 36081 13991 36139 13997
rect 36081 13988 36093 13991
rect 33888 13960 36093 13988
rect 36081 13957 36093 13960
rect 36127 13957 36139 13991
rect 36188 13988 36216 14028
rect 36449 14025 36461 14059
rect 36495 14056 36507 14059
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 36495 14028 37841 14056
rect 36495 14025 36507 14028
rect 36449 14019 36507 14025
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 37829 14019 37887 14025
rect 38197 14059 38255 14065
rect 38197 14025 38209 14059
rect 38243 14056 38255 14059
rect 41322 14056 41328 14068
rect 38243 14028 41328 14056
rect 38243 14025 38255 14028
rect 38197 14019 38255 14025
rect 41322 14016 41328 14028
rect 41380 14016 41386 14068
rect 45833 14059 45891 14065
rect 45833 14025 45845 14059
rect 45879 14056 45891 14059
rect 47854 14056 47860 14068
rect 45879 14028 47860 14056
rect 45879 14025 45891 14028
rect 45833 14019 45891 14025
rect 47854 14016 47860 14028
rect 47912 14016 47918 14068
rect 48406 14016 48412 14068
rect 48464 14016 48470 14068
rect 48866 14016 48872 14068
rect 48924 14056 48930 14068
rect 49145 14059 49203 14065
rect 49145 14056 49157 14059
rect 48924 14028 49157 14056
rect 48924 14016 48930 14028
rect 49145 14025 49157 14028
rect 49191 14025 49203 14059
rect 49145 14019 49203 14025
rect 36188 13960 36492 13988
rect 36081 13951 36139 13957
rect 26605 13923 26663 13929
rect 26605 13889 26617 13923
rect 26651 13889 26663 13923
rect 26605 13883 26663 13889
rect 28902 13880 28908 13932
rect 28960 13880 28966 13932
rect 31110 13880 31116 13932
rect 31168 13880 31174 13932
rect 34698 13880 34704 13932
rect 34756 13920 34762 13932
rect 34793 13923 34851 13929
rect 34793 13920 34805 13923
rect 34756 13892 34805 13920
rect 34756 13880 34762 13892
rect 34793 13889 34805 13892
rect 34839 13889 34851 13923
rect 36170 13920 36176 13932
rect 34793 13883 34851 13889
rect 35912 13892 36176 13920
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13821 14795 13855
rect 14737 13815 14795 13821
rect 15102 13812 15108 13864
rect 15160 13852 15166 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15160 13824 16129 13852
rect 15160 13812 15166 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 12124 13756 12434 13784
rect 12124 13744 12130 13756
rect 14458 13744 14464 13796
rect 14516 13784 14522 13796
rect 17788 13784 17816 13815
rect 18598 13812 18604 13864
rect 18656 13852 18662 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18656 13824 18889 13852
rect 18656 13812 18662 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19024 13824 19717 13852
rect 19024 13812 19030 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19981 13855 20039 13861
rect 19981 13821 19993 13855
rect 20027 13852 20039 13855
rect 20714 13852 20720 13864
rect 20027 13824 20720 13852
rect 20027 13821 20039 13824
rect 19981 13815 20039 13821
rect 20714 13812 20720 13824
rect 20772 13852 20778 13864
rect 21910 13852 21916 13864
rect 20772 13824 21916 13852
rect 20772 13812 20778 13824
rect 21910 13812 21916 13824
rect 21968 13852 21974 13864
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 21968 13824 22017 13852
rect 21968 13812 21974 13824
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 23753 13855 23811 13861
rect 23753 13821 23765 13855
rect 23799 13821 23811 13855
rect 23753 13815 23811 13821
rect 17954 13784 17960 13796
rect 14516 13756 16896 13784
rect 17788 13756 17960 13784
rect 14516 13744 14522 13756
rect 12342 13716 12348 13728
rect 9824 13688 12348 13716
rect 9824 13676 9830 13688
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12437 13719 12495 13725
rect 12437 13685 12449 13719
rect 12483 13716 12495 13719
rect 12710 13716 12716 13728
rect 12483 13688 12716 13716
rect 12483 13685 12495 13688
rect 12437 13679 12495 13685
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 15289 13719 15347 13725
rect 15289 13685 15301 13719
rect 15335 13716 15347 13719
rect 16298 13716 16304 13728
rect 15335 13688 16304 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 16868 13716 16896 13756
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 23768 13784 23796 13815
rect 23934 13812 23940 13864
rect 23992 13852 23998 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23992 13824 24225 13852
rect 23992 13812 23998 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 27062 13812 27068 13864
rect 27120 13852 27126 13864
rect 29365 13855 29423 13861
rect 29365 13852 29377 13855
rect 27120 13824 29377 13852
rect 27120 13812 27126 13824
rect 29365 13821 29377 13824
rect 29411 13821 29423 13855
rect 29365 13815 29423 13821
rect 30837 13855 30895 13861
rect 30837 13821 30849 13855
rect 30883 13852 30895 13855
rect 32306 13852 32312 13864
rect 30883 13824 31064 13852
rect 30883 13821 30895 13824
rect 30837 13815 30895 13821
rect 24578 13784 24584 13796
rect 23768 13756 24584 13784
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 31036 13784 31064 13824
rect 31726 13824 32312 13852
rect 31726 13784 31754 13824
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 34054 13812 34060 13864
rect 34112 13812 34118 13864
rect 35912 13861 35940 13892
rect 36170 13880 36176 13892
rect 36228 13920 36234 13932
rect 36354 13920 36360 13932
rect 36228 13892 36360 13920
rect 36228 13880 36234 13892
rect 36354 13880 36360 13892
rect 36412 13880 36418 13932
rect 36464 13920 36492 13960
rect 36722 13948 36728 14000
rect 36780 13988 36786 14000
rect 37737 13991 37795 13997
rect 37737 13988 37749 13991
rect 36780 13960 37749 13988
rect 36780 13948 36786 13960
rect 37737 13957 37749 13960
rect 37783 13957 37795 13991
rect 37737 13951 37795 13957
rect 38565 13991 38623 13997
rect 38565 13957 38577 13991
rect 38611 13988 38623 13991
rect 38654 13988 38660 14000
rect 38611 13960 38660 13988
rect 38611 13957 38623 13960
rect 38565 13951 38623 13957
rect 38654 13948 38660 13960
rect 38712 13988 38718 14000
rect 38838 13988 38844 14000
rect 38712 13960 38844 13988
rect 38712 13948 38718 13960
rect 38838 13948 38844 13960
rect 38896 13988 38902 14000
rect 38933 13991 38991 13997
rect 38933 13988 38945 13991
rect 38896 13960 38945 13988
rect 38896 13948 38902 13960
rect 38933 13957 38945 13960
rect 38979 13957 38991 13991
rect 38933 13951 38991 13957
rect 39482 13948 39488 14000
rect 39540 13988 39546 14000
rect 45005 13991 45063 13997
rect 45005 13988 45017 13991
rect 39540 13960 45017 13988
rect 39540 13948 39546 13960
rect 45005 13957 45017 13960
rect 45051 13957 45063 13991
rect 45005 13951 45063 13957
rect 48133 13991 48191 13997
rect 48133 13957 48145 13991
rect 48179 13988 48191 13991
rect 49234 13988 49240 14000
rect 48179 13960 49240 13988
rect 48179 13957 48191 13960
rect 48133 13951 48191 13957
rect 49234 13948 49240 13960
rect 49292 13948 49298 14000
rect 36909 13923 36967 13929
rect 36909 13920 36921 13923
rect 36464 13892 36921 13920
rect 36909 13889 36921 13892
rect 36955 13889 36967 13923
rect 36909 13883 36967 13889
rect 45646 13880 45652 13932
rect 45704 13880 45710 13932
rect 48222 13880 48228 13932
rect 48280 13920 48286 13932
rect 48593 13923 48651 13929
rect 48593 13920 48605 13923
rect 48280 13892 48605 13920
rect 48280 13880 48286 13892
rect 48593 13889 48605 13892
rect 48639 13889 48651 13923
rect 48593 13883 48651 13889
rect 34609 13855 34667 13861
rect 34609 13821 34621 13855
rect 34655 13821 34667 13855
rect 34609 13815 34667 13821
rect 35897 13855 35955 13861
rect 35897 13821 35909 13855
rect 35943 13821 35955 13855
rect 35897 13815 35955 13821
rect 31036 13756 31754 13784
rect 34624 13784 34652 13815
rect 35986 13812 35992 13864
rect 36044 13812 36050 13864
rect 36262 13812 36268 13864
rect 36320 13852 36326 13864
rect 36630 13852 36636 13864
rect 36320 13824 36636 13852
rect 36320 13812 36326 13824
rect 36630 13812 36636 13824
rect 36688 13852 36694 13864
rect 36725 13855 36783 13861
rect 36725 13852 36737 13855
rect 36688 13824 36737 13852
rect 36688 13812 36694 13824
rect 36725 13821 36737 13824
rect 36771 13821 36783 13855
rect 36725 13815 36783 13821
rect 37645 13855 37703 13861
rect 37645 13821 37657 13855
rect 37691 13821 37703 13855
rect 37645 13815 37703 13821
rect 45189 13855 45247 13861
rect 45189 13821 45201 13855
rect 45235 13852 45247 13855
rect 46566 13852 46572 13864
rect 45235 13824 46572 13852
rect 45235 13821 45247 13824
rect 45189 13815 45247 13821
rect 34698 13784 34704 13796
rect 34624 13756 34704 13784
rect 34698 13744 34704 13756
rect 34756 13744 34762 13796
rect 37660 13784 37688 13815
rect 46566 13812 46572 13824
rect 46624 13812 46630 13864
rect 38194 13784 38200 13796
rect 37660 13756 38200 13784
rect 38194 13744 38200 13756
rect 38252 13744 38258 13796
rect 23106 13716 23112 13728
rect 16868 13688 23112 13716
rect 23106 13676 23112 13688
rect 23164 13676 23170 13728
rect 24670 13676 24676 13728
rect 24728 13716 24734 13728
rect 25682 13716 25688 13728
rect 24728 13688 25688 13716
rect 24728 13676 24734 13688
rect 25682 13676 25688 13688
rect 25740 13676 25746 13728
rect 30834 13676 30840 13728
rect 30892 13716 30898 13728
rect 33799 13719 33857 13725
rect 33799 13716 33811 13719
rect 30892 13688 33811 13716
rect 30892 13676 30898 13688
rect 33799 13685 33811 13688
rect 33845 13716 33857 13719
rect 35894 13716 35900 13728
rect 33845 13688 35900 13716
rect 33845 13685 33857 13688
rect 33799 13679 33857 13685
rect 35894 13676 35900 13688
rect 35952 13676 35958 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 2976 13484 12664 13512
rect 1762 13336 1768 13388
rect 1820 13336 1826 13388
rect 2976 13317 3004 13484
rect 12636 13444 12664 13484
rect 13722 13472 13728 13524
rect 13780 13472 13786 13524
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 13998 13512 14004 13524
rect 13955 13484 14004 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 13998 13472 14004 13484
rect 14056 13512 14062 13524
rect 15010 13512 15016 13524
rect 14056 13484 15016 13512
rect 14056 13472 14062 13484
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 17954 13512 17960 13524
rect 15396 13484 17960 13512
rect 14277 13447 14335 13453
rect 14277 13444 14289 13447
rect 12636 13416 14289 13444
rect 14277 13413 14289 13416
rect 14323 13413 14335 13447
rect 14277 13407 14335 13413
rect 14734 13404 14740 13456
rect 14792 13444 14798 13456
rect 14829 13447 14887 13453
rect 14829 13444 14841 13447
rect 14792 13416 14841 13444
rect 14792 13404 14798 13416
rect 14829 13413 14841 13416
rect 14875 13413 14887 13447
rect 14829 13407 14887 13413
rect 10778 13336 10784 13388
rect 10836 13376 10842 13388
rect 12066 13376 12072 13388
rect 10836 13348 12072 13376
rect 10836 13336 10842 13348
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 12400 13348 12541 13376
rect 12400 13336 12406 13348
rect 12529 13345 12541 13348
rect 12575 13376 12587 13379
rect 12575 13348 12664 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 11057 13243 11115 13249
rect 11057 13240 11069 13243
rect 9088 13212 11069 13240
rect 9088 13200 9094 13212
rect 11057 13209 11069 13212
rect 11103 13209 11115 13243
rect 12342 13240 12348 13252
rect 12282 13212 12348 13240
rect 11057 13203 11115 13209
rect 10505 13175 10563 13181
rect 10505 13141 10517 13175
rect 10551 13172 10563 13175
rect 10870 13172 10876 13184
rect 10551 13144 10876 13172
rect 10551 13141 10563 13144
rect 10505 13135 10563 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11072 13172 11100 13203
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 12636 13240 12664 13348
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12860 13348 13093 13376
rect 12860 13336 12866 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 13998 13376 14004 13388
rect 13872 13348 14004 13376
rect 13872 13336 13878 13348
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 15102 13376 15108 13388
rect 14292 13348 15108 13376
rect 14292 13320 14320 13348
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15396 13385 15424 13484
rect 17954 13472 17960 13484
rect 18012 13512 18018 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 18012 13484 18153 13512
rect 18012 13472 18018 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 18414 13512 18420 13524
rect 18187 13484 18420 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19208 13484 19441 13512
rect 19208 13472 19214 13484
rect 19429 13481 19441 13484
rect 19475 13512 19487 13515
rect 20070 13512 20076 13524
rect 19475 13484 20076 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20254 13472 20260 13524
rect 20312 13512 20318 13524
rect 20441 13515 20499 13521
rect 20441 13512 20453 13515
rect 20312 13484 20453 13512
rect 20312 13472 20318 13484
rect 20441 13481 20453 13484
rect 20487 13481 20499 13515
rect 20441 13475 20499 13481
rect 20898 13472 20904 13524
rect 20956 13472 20962 13524
rect 22094 13472 22100 13524
rect 22152 13472 22158 13524
rect 22738 13512 22744 13524
rect 22572 13484 22744 13512
rect 16114 13404 16120 13456
rect 16172 13444 16178 13456
rect 16172 13416 16528 13444
rect 16172 13404 16178 13416
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 15470 13336 15476 13388
rect 15528 13336 15534 13388
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16298 13376 16304 13388
rect 15804 13348 16304 13376
rect 15804 13336 15810 13348
rect 16298 13336 16304 13348
rect 16356 13376 16362 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 16356 13348 16405 13376
rect 16356 13336 16362 13348
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16500 13376 16528 13416
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 22462 13444 22468 13456
rect 18564 13416 22468 13444
rect 18564 13404 18570 13416
rect 22462 13404 22468 13416
rect 22520 13404 22526 13456
rect 16669 13379 16727 13385
rect 16669 13376 16681 13379
rect 16500 13348 16681 13376
rect 16393 13339 16451 13345
rect 16669 13345 16681 13348
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13376 19947 13379
rect 20714 13376 20720 13388
rect 19935 13348 20720 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 21358 13336 21364 13388
rect 21416 13376 21422 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 21416 13348 21465 13376
rect 21416 13336 21422 13348
rect 21453 13345 21465 13348
rect 21499 13376 21511 13379
rect 22572 13376 22600 13484
rect 22738 13472 22744 13484
rect 22796 13472 22802 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 24029 13515 24087 13521
rect 24029 13512 24041 13515
rect 23716 13484 24041 13512
rect 23716 13472 23722 13484
rect 24029 13481 24041 13484
rect 24075 13481 24087 13515
rect 24029 13475 24087 13481
rect 25590 13472 25596 13524
rect 25648 13472 25654 13524
rect 25774 13472 25780 13524
rect 25832 13512 25838 13524
rect 26697 13515 26755 13521
rect 26697 13512 26709 13515
rect 25832 13484 26709 13512
rect 25832 13472 25838 13484
rect 26697 13481 26709 13484
rect 26743 13512 26755 13515
rect 27433 13515 27491 13521
rect 27433 13512 27445 13515
rect 26743 13484 27445 13512
rect 26743 13481 26755 13484
rect 26697 13475 26755 13481
rect 27433 13481 27445 13484
rect 27479 13512 27491 13515
rect 27522 13512 27528 13524
rect 27479 13484 27528 13512
rect 27479 13481 27491 13484
rect 27433 13475 27491 13481
rect 27522 13472 27528 13484
rect 27580 13472 27586 13524
rect 27706 13472 27712 13524
rect 27764 13472 27770 13524
rect 27798 13472 27804 13524
rect 27856 13472 27862 13524
rect 28169 13515 28227 13521
rect 28169 13481 28181 13515
rect 28215 13512 28227 13515
rect 28350 13512 28356 13524
rect 28215 13484 28356 13512
rect 28215 13481 28227 13484
rect 28169 13475 28227 13481
rect 28350 13472 28356 13484
rect 28408 13512 28414 13524
rect 28902 13512 28908 13524
rect 28408 13484 28908 13512
rect 28408 13472 28414 13484
rect 28902 13472 28908 13484
rect 28960 13472 28966 13524
rect 29181 13515 29239 13521
rect 29181 13481 29193 13515
rect 29227 13512 29239 13515
rect 33778 13512 33784 13524
rect 29227 13484 33784 13512
rect 29227 13481 29239 13484
rect 29181 13475 29239 13481
rect 33778 13472 33784 13484
rect 33836 13472 33842 13524
rect 35526 13472 35532 13524
rect 35584 13512 35590 13524
rect 35621 13515 35679 13521
rect 35621 13512 35633 13515
rect 35584 13484 35633 13512
rect 35584 13472 35590 13484
rect 35621 13481 35633 13484
rect 35667 13481 35679 13515
rect 35621 13475 35679 13481
rect 35989 13515 36047 13521
rect 35989 13481 36001 13515
rect 36035 13512 36047 13515
rect 36262 13512 36268 13524
rect 36035 13484 36268 13512
rect 36035 13481 36047 13484
rect 35989 13475 36047 13481
rect 36262 13472 36268 13484
rect 36320 13472 36326 13524
rect 36556 13484 38148 13512
rect 24854 13404 24860 13456
rect 24912 13444 24918 13456
rect 25792 13444 25820 13472
rect 29914 13444 29920 13456
rect 24912 13416 25820 13444
rect 28644 13416 29920 13444
rect 24912 13404 24918 13416
rect 21499 13348 22600 13376
rect 22741 13379 22799 13385
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 22741 13345 22753 13379
rect 22787 13376 22799 13379
rect 23014 13376 23020 13388
rect 22787 13348 23020 13376
rect 22787 13345 22799 13348
rect 22741 13339 22799 13345
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13345 23535 13379
rect 23477 13339 23535 13345
rect 23569 13379 23627 13385
rect 23569 13345 23581 13379
rect 23615 13376 23627 13379
rect 24026 13376 24032 13388
rect 23615 13348 24032 13376
rect 23615 13345 23627 13348
rect 23569 13339 23627 13345
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 14458 13268 14464 13320
rect 14516 13268 14522 13320
rect 15562 13268 15568 13320
rect 15620 13268 15626 13320
rect 23492 13308 23520 13339
rect 24026 13336 24032 13348
rect 24084 13376 24090 13388
rect 24394 13376 24400 13388
rect 24084 13348 24400 13376
rect 24084 13336 24090 13348
rect 24394 13336 24400 13348
rect 24452 13336 24458 13388
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13376 25099 13379
rect 27062 13376 27068 13388
rect 25087 13348 27068 13376
rect 25087 13345 25099 13348
rect 25041 13339 25099 13345
rect 27062 13336 27068 13348
rect 27120 13336 27126 13388
rect 28644 13385 28672 13416
rect 29914 13404 29920 13416
rect 29972 13404 29978 13456
rect 30374 13404 30380 13456
rect 30432 13444 30438 13456
rect 31113 13447 31171 13453
rect 31113 13444 31125 13447
rect 30432 13416 31125 13444
rect 30432 13404 30438 13416
rect 31113 13413 31125 13416
rect 31159 13413 31171 13447
rect 31113 13407 31171 13413
rect 33321 13447 33379 13453
rect 33321 13413 33333 13447
rect 33367 13413 33379 13447
rect 33321 13407 33379 13413
rect 28629 13379 28687 13385
rect 28629 13345 28641 13379
rect 28675 13345 28687 13379
rect 28629 13339 28687 13345
rect 29822 13336 29828 13388
rect 29880 13336 29886 13388
rect 30009 13379 30067 13385
rect 30009 13345 30021 13379
rect 30055 13376 30067 13379
rect 30466 13376 30472 13388
rect 30055 13348 30472 13376
rect 30055 13345 30067 13348
rect 30009 13339 30067 13345
rect 30466 13336 30472 13348
rect 30524 13336 30530 13388
rect 31570 13336 31576 13388
rect 31628 13376 31634 13388
rect 33336 13376 33364 13407
rect 33686 13404 33692 13456
rect 33744 13444 33750 13456
rect 36081 13447 36139 13453
rect 36081 13444 36093 13447
rect 33744 13416 36093 13444
rect 33744 13404 33750 13416
rect 36081 13413 36093 13416
rect 36127 13413 36139 13447
rect 36556 13444 36584 13484
rect 36081 13407 36139 13413
rect 36280 13416 36584 13444
rect 38120 13444 38148 13484
rect 38194 13472 38200 13524
rect 38252 13472 38258 13524
rect 38565 13515 38623 13521
rect 38565 13481 38577 13515
rect 38611 13512 38623 13515
rect 38838 13512 38844 13524
rect 38611 13484 38844 13512
rect 38611 13481 38623 13484
rect 38565 13475 38623 13481
rect 38838 13472 38844 13484
rect 38896 13512 38902 13524
rect 39577 13515 39635 13521
rect 39577 13512 39589 13515
rect 38896 13484 39589 13512
rect 38896 13472 38902 13484
rect 39577 13481 39589 13484
rect 39623 13481 39635 13515
rect 39577 13475 39635 13481
rect 39206 13444 39212 13456
rect 38120 13416 39212 13444
rect 31628 13348 33364 13376
rect 31628 13336 31634 13348
rect 33870 13336 33876 13388
rect 33928 13376 33934 13388
rect 34333 13379 34391 13385
rect 34333 13376 34345 13379
rect 33928 13348 34345 13376
rect 33928 13336 33934 13348
rect 34333 13345 34345 13348
rect 34379 13345 34391 13379
rect 34333 13339 34391 13345
rect 35069 13379 35127 13385
rect 35069 13345 35081 13379
rect 35115 13376 35127 13379
rect 36280 13376 36308 13416
rect 39206 13404 39212 13416
rect 39264 13404 39270 13456
rect 35115 13348 36308 13376
rect 35115 13345 35127 13348
rect 35069 13339 35127 13345
rect 36354 13336 36360 13388
rect 36412 13376 36418 13388
rect 36725 13379 36783 13385
rect 36725 13376 36737 13379
rect 36412 13348 36737 13376
rect 36412 13336 36418 13348
rect 36725 13345 36737 13348
rect 36771 13345 36783 13379
rect 36725 13339 36783 13345
rect 36814 13336 36820 13388
rect 36872 13376 36878 13388
rect 39482 13376 39488 13388
rect 36872 13348 39488 13376
rect 36872 13336 36878 13348
rect 39482 13336 39488 13348
rect 39540 13336 39546 13388
rect 24670 13308 24676 13320
rect 23492 13280 24676 13308
rect 24670 13268 24676 13280
rect 24728 13268 24734 13320
rect 25130 13268 25136 13320
rect 25188 13308 25194 13320
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 25188 13280 25237 13308
rect 25188 13268 25194 13280
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 27430 13308 27436 13320
rect 25225 13271 25283 13277
rect 25332 13280 27436 13308
rect 14918 13240 14924 13252
rect 12636 13212 14924 13240
rect 14918 13200 14924 13212
rect 14976 13200 14982 13252
rect 15856 13212 17080 13240
rect 13814 13172 13820 13184
rect 11020 13144 13820 13172
rect 11020 13132 11026 13144
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 15856 13172 15884 13212
rect 14148 13144 15884 13172
rect 14148 13132 14154 13144
rect 15930 13132 15936 13184
rect 15988 13132 15994 13184
rect 17052 13172 17080 13212
rect 17126 13200 17132 13252
rect 17184 13200 17190 13252
rect 18877 13243 18935 13249
rect 18877 13209 18889 13243
rect 18923 13240 18935 13243
rect 20073 13243 20131 13249
rect 20073 13240 20085 13243
rect 18923 13212 20085 13240
rect 18923 13209 18935 13212
rect 18877 13203 18935 13209
rect 20073 13209 20085 13212
rect 20119 13209 20131 13243
rect 20073 13203 20131 13209
rect 21174 13200 21180 13252
rect 21232 13240 21238 13252
rect 21361 13243 21419 13249
rect 21361 13240 21373 13243
rect 21232 13212 21373 13240
rect 21232 13200 21238 13212
rect 21361 13209 21373 13212
rect 21407 13240 21419 13243
rect 21634 13240 21640 13252
rect 21407 13212 21640 13240
rect 21407 13209 21419 13212
rect 21361 13203 21419 13209
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 22465 13243 22523 13249
rect 22465 13209 22477 13243
rect 22511 13240 22523 13243
rect 22830 13240 22836 13252
rect 22511 13212 22836 13240
rect 22511 13209 22523 13212
rect 22465 13203 22523 13209
rect 22830 13200 22836 13212
rect 22888 13200 22894 13252
rect 23658 13200 23664 13252
rect 23716 13200 23722 13252
rect 25332 13240 25360 13280
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 28813 13311 28871 13317
rect 28813 13277 28825 13311
rect 28859 13308 28871 13311
rect 28994 13308 29000 13320
rect 28859 13280 29000 13308
rect 28859 13277 28871 13280
rect 28813 13271 28871 13277
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30190 13308 30196 13320
rect 30147 13280 30196 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 32861 13311 32919 13317
rect 32861 13277 32873 13311
rect 32907 13308 32919 13311
rect 34054 13308 34060 13320
rect 32907 13280 34060 13308
rect 32907 13277 32919 13280
rect 32861 13271 32919 13277
rect 34054 13268 34060 13280
rect 34112 13268 34118 13320
rect 34882 13268 34888 13320
rect 34940 13308 34946 13320
rect 36449 13311 36507 13317
rect 36449 13308 36461 13311
rect 34940 13280 36461 13308
rect 34940 13268 34946 13280
rect 36449 13277 36461 13280
rect 36495 13277 36507 13311
rect 36449 13271 36507 13277
rect 23768 13212 25360 13240
rect 19886 13172 19892 13184
rect 17052 13144 19892 13172
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13172 20039 13175
rect 20254 13172 20260 13184
rect 20027 13144 20260 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 21266 13132 21272 13184
rect 21324 13172 21330 13184
rect 21726 13172 21732 13184
rect 21324 13144 21732 13172
rect 21324 13132 21330 13144
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 22557 13175 22615 13181
rect 22557 13141 22569 13175
rect 22603 13172 22615 13175
rect 23768 13172 23796 13212
rect 26050 13200 26056 13252
rect 26108 13200 26114 13252
rect 32585 13243 32643 13249
rect 30484 13212 31340 13240
rect 32154 13212 32536 13240
rect 22603 13144 23796 13172
rect 22603 13141 22615 13144
rect 22557 13135 22615 13141
rect 23842 13132 23848 13184
rect 23900 13172 23906 13184
rect 24489 13175 24547 13181
rect 24489 13172 24501 13175
rect 23900 13144 24501 13172
rect 23900 13132 23906 13144
rect 24489 13141 24501 13144
rect 24535 13172 24547 13175
rect 25133 13175 25191 13181
rect 25133 13172 25145 13175
rect 24535 13144 25145 13172
rect 24535 13141 24547 13144
rect 24489 13135 24547 13141
rect 25133 13141 25145 13144
rect 25179 13172 25191 13175
rect 26510 13172 26516 13184
rect 25179 13144 26516 13172
rect 25179 13141 25191 13144
rect 25133 13135 25191 13141
rect 26510 13132 26516 13144
rect 26568 13132 26574 13184
rect 28718 13132 28724 13184
rect 28776 13132 28782 13184
rect 30484 13181 30512 13212
rect 30469 13175 30527 13181
rect 30469 13141 30481 13175
rect 30515 13141 30527 13175
rect 31312 13172 31340 13212
rect 31662 13172 31668 13184
rect 31312 13144 31668 13172
rect 30469 13135 30527 13141
rect 31662 13132 31668 13144
rect 31720 13132 31726 13184
rect 31846 13132 31852 13184
rect 31904 13172 31910 13184
rect 32232 13172 32260 13212
rect 31904 13144 32260 13172
rect 32508 13172 32536 13212
rect 32585 13209 32597 13243
rect 32631 13240 32643 13243
rect 33962 13240 33968 13252
rect 32631 13212 33968 13240
rect 32631 13209 32643 13212
rect 32585 13203 32643 13209
rect 33962 13200 33968 13212
rect 34020 13200 34026 13252
rect 35158 13200 35164 13252
rect 35216 13200 35222 13252
rect 35253 13243 35311 13249
rect 35253 13209 35265 13243
rect 35299 13240 35311 13243
rect 36354 13240 36360 13252
rect 35299 13212 36360 13240
rect 35299 13209 35311 13212
rect 35253 13203 35311 13209
rect 36354 13200 36360 13212
rect 36412 13200 36418 13252
rect 36464 13240 36492 13271
rect 41322 13268 41328 13320
rect 41380 13268 41386 13320
rect 46566 13268 46572 13320
rect 46624 13308 46630 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 46624 13280 47961 13308
rect 46624 13268 46630 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 49142 13268 49148 13320
rect 49200 13268 49206 13320
rect 36464 13212 36584 13240
rect 33318 13172 33324 13184
rect 32508 13144 33324 13172
rect 31904 13132 31910 13144
rect 33318 13132 33324 13144
rect 33376 13132 33382 13184
rect 33686 13132 33692 13184
rect 33744 13132 33750 13184
rect 33781 13175 33839 13181
rect 33781 13141 33793 13175
rect 33827 13172 33839 13175
rect 34330 13172 34336 13184
rect 33827 13144 34336 13172
rect 33827 13141 33839 13144
rect 33781 13135 33839 13141
rect 34330 13132 34336 13144
rect 34388 13132 34394 13184
rect 36556 13172 36584 13212
rect 36630 13200 36636 13252
rect 36688 13240 36694 13252
rect 36688 13212 37214 13240
rect 36688 13200 36694 13212
rect 37458 13172 37464 13184
rect 36556 13144 37464 13172
rect 37458 13132 37464 13144
rect 37516 13132 37522 13184
rect 37642 13132 37648 13184
rect 37700 13172 37706 13184
rect 39298 13172 39304 13184
rect 37700 13144 39304 13172
rect 37700 13132 37706 13144
rect 39298 13132 39304 13144
rect 39356 13132 39362 13184
rect 41509 13175 41567 13181
rect 41509 13141 41521 13175
rect 41555 13172 41567 13175
rect 45922 13172 45928 13184
rect 41555 13144 45928 13172
rect 41555 13141 41567 13144
rect 41509 13135 41567 13141
rect 45922 13132 45928 13144
rect 45980 13132 45986 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12968 3111 12971
rect 5442 12968 5448 12980
rect 3099 12940 5448 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 10962 12928 10968 12980
rect 11020 12928 11026 12980
rect 11146 12928 11152 12980
rect 11204 12928 11210 12980
rect 11974 12928 11980 12980
rect 12032 12928 12038 12980
rect 12069 12971 12127 12977
rect 12069 12937 12081 12971
rect 12115 12968 12127 12971
rect 12158 12968 12164 12980
rect 12115 12940 12164 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12713 12971 12771 12977
rect 12713 12968 12725 12971
rect 12584 12940 12725 12968
rect 12584 12928 12590 12940
rect 12713 12937 12725 12940
rect 12759 12937 12771 12971
rect 12713 12931 12771 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13262 12968 13268 12980
rect 13127 12940 13268 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13630 12928 13636 12980
rect 13688 12968 13694 12980
rect 13688 12940 14964 12968
rect 13688 12928 13694 12940
rect 1302 12860 1308 12912
rect 1360 12900 1366 12912
rect 1673 12903 1731 12909
rect 1673 12900 1685 12903
rect 1360 12872 1685 12900
rect 1360 12860 1366 12872
rect 1673 12869 1685 12872
rect 1719 12900 1731 12903
rect 2133 12903 2191 12909
rect 2133 12900 2145 12903
rect 1719 12872 2145 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 2133 12869 2145 12872
rect 2179 12869 2191 12903
rect 14642 12900 14648 12912
rect 14122 12872 14648 12900
rect 2133 12863 2191 12869
rect 14642 12860 14648 12872
rect 14700 12860 14706 12912
rect 14936 12900 14964 12940
rect 15010 12928 15016 12980
rect 15068 12968 15074 12980
rect 15197 12971 15255 12977
rect 15197 12968 15209 12971
rect 15068 12940 15209 12968
rect 15068 12928 15074 12940
rect 15197 12937 15209 12940
rect 15243 12937 15255 12971
rect 15197 12931 15255 12937
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 15896 12940 19104 12968
rect 15896 12928 15902 12940
rect 15470 12900 15476 12912
rect 14936 12872 15476 12900
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 15933 12903 15991 12909
rect 15933 12869 15945 12903
rect 15979 12900 15991 12903
rect 16206 12900 16212 12912
rect 15979 12872 16212 12900
rect 15979 12869 15991 12872
rect 15933 12863 15991 12869
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 16298 12860 16304 12912
rect 16356 12900 16362 12912
rect 18693 12903 18751 12909
rect 18693 12900 18705 12903
rect 16356 12872 18705 12900
rect 16356 12860 16362 12872
rect 18693 12869 18705 12872
rect 18739 12900 18751 12903
rect 18966 12900 18972 12912
rect 18739 12872 18972 12900
rect 18739 12869 18751 12872
rect 18693 12863 18751 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 19076 12900 19104 12940
rect 20714 12928 20720 12980
rect 20772 12928 20778 12980
rect 21177 12971 21235 12977
rect 21177 12937 21189 12971
rect 21223 12968 21235 12971
rect 22646 12968 22652 12980
rect 21223 12940 22652 12968
rect 21223 12937 21235 12940
rect 21177 12931 21235 12937
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 22922 12928 22928 12980
rect 22980 12928 22986 12980
rect 23014 12928 23020 12980
rect 23072 12968 23078 12980
rect 23658 12968 23664 12980
rect 23072 12940 23664 12968
rect 23072 12928 23078 12940
rect 23658 12928 23664 12940
rect 23716 12928 23722 12980
rect 24578 12928 24584 12980
rect 24636 12968 24642 12980
rect 24636 12940 25636 12968
rect 24636 12928 24642 12940
rect 23842 12900 23848 12912
rect 19076 12872 23848 12900
rect 23842 12860 23848 12872
rect 23900 12860 23906 12912
rect 24854 12860 24860 12912
rect 24912 12860 24918 12912
rect 25314 12860 25320 12912
rect 25372 12860 25378 12912
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 1268 12804 2881 12832
rect 1268 12792 1274 12804
rect 2869 12801 2881 12804
rect 2915 12832 2927 12835
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 2915 12804 3341 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12832 17003 12835
rect 17034 12832 17040 12844
rect 16991 12804 17040 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18874 12832 18880 12844
rect 17911 12804 18880 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19610 12792 19616 12844
rect 19668 12792 19674 12844
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 21910 12832 21916 12844
rect 21131 12804 21916 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 22646 12832 22652 12844
rect 22244 12804 22652 12832
rect 22244 12792 22250 12804
rect 22646 12792 22652 12804
rect 22704 12832 22710 12844
rect 25608 12841 25636 12940
rect 25774 12928 25780 12980
rect 25832 12968 25838 12980
rect 26053 12971 26111 12977
rect 26053 12968 26065 12971
rect 25832 12940 26065 12968
rect 25832 12928 25838 12940
rect 26053 12937 26065 12940
rect 26099 12937 26111 12971
rect 26053 12931 26111 12937
rect 26329 12971 26387 12977
rect 26329 12937 26341 12971
rect 26375 12968 26387 12971
rect 26418 12968 26424 12980
rect 26375 12940 26424 12968
rect 26375 12937 26387 12940
rect 26329 12931 26387 12937
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 26510 12928 26516 12980
rect 26568 12968 26574 12980
rect 26697 12971 26755 12977
rect 26697 12968 26709 12971
rect 26568 12940 26709 12968
rect 26568 12928 26574 12940
rect 26697 12937 26709 12940
rect 26743 12968 26755 12971
rect 27062 12968 27068 12980
rect 26743 12940 27068 12968
rect 26743 12937 26755 12940
rect 26697 12931 26755 12937
rect 27062 12928 27068 12940
rect 27120 12928 27126 12980
rect 27890 12928 27896 12980
rect 27948 12968 27954 12980
rect 31757 12971 31815 12977
rect 27948 12940 31616 12968
rect 27948 12928 27954 12940
rect 27522 12860 27528 12912
rect 27580 12900 27586 12912
rect 27580 12872 27738 12900
rect 27580 12860 27586 12872
rect 29638 12860 29644 12912
rect 29696 12860 29702 12912
rect 30190 12860 30196 12912
rect 30248 12900 30254 12912
rect 30285 12903 30343 12909
rect 30285 12900 30297 12903
rect 30248 12872 30297 12900
rect 30248 12860 30254 12872
rect 30285 12869 30297 12872
rect 30331 12869 30343 12903
rect 31588 12900 31616 12940
rect 31757 12937 31769 12971
rect 31803 12968 31815 12971
rect 32398 12968 32404 12980
rect 31803 12940 32404 12968
rect 31803 12937 31815 12940
rect 31757 12931 31815 12937
rect 32398 12928 32404 12940
rect 32456 12968 32462 12980
rect 32582 12968 32588 12980
rect 32456 12940 32588 12968
rect 32456 12928 32462 12940
rect 32582 12928 32588 12940
rect 32640 12928 32646 12980
rect 33413 12971 33471 12977
rect 33413 12937 33425 12971
rect 33459 12968 33471 12971
rect 33686 12968 33692 12980
rect 33459 12940 33692 12968
rect 33459 12937 33471 12940
rect 33413 12931 33471 12937
rect 33686 12928 33692 12940
rect 33744 12928 33750 12980
rect 34054 12928 34060 12980
rect 34112 12968 34118 12980
rect 34112 12940 34836 12968
rect 34112 12928 34118 12940
rect 34808 12909 34836 12940
rect 35158 12928 35164 12980
rect 35216 12968 35222 12980
rect 36449 12971 36507 12977
rect 36449 12968 36461 12971
rect 35216 12940 36461 12968
rect 35216 12928 35222 12940
rect 36449 12937 36461 12940
rect 36495 12968 36507 12971
rect 40310 12968 40316 12980
rect 36495 12940 40316 12968
rect 36495 12937 36507 12940
rect 36449 12931 36507 12937
rect 40310 12928 40316 12940
rect 40368 12928 40374 12980
rect 32677 12903 32735 12909
rect 32677 12900 32689 12903
rect 31588 12872 32689 12900
rect 30285 12863 30343 12869
rect 32677 12869 32689 12872
rect 32723 12869 32735 12903
rect 32677 12863 32735 12869
rect 34793 12903 34851 12909
rect 34793 12869 34805 12903
rect 34839 12900 34851 12903
rect 34882 12900 34888 12912
rect 34839 12872 34888 12900
rect 34839 12869 34851 12872
rect 34793 12863 34851 12869
rect 34882 12860 34888 12872
rect 34940 12860 34946 12912
rect 35802 12860 35808 12912
rect 35860 12900 35866 12912
rect 35860 12872 35940 12900
rect 35860 12860 35866 12872
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22704 12804 23029 12832
rect 22704 12792 22710 12804
rect 23017 12801 23029 12804
rect 23063 12832 23075 12835
rect 25593 12835 25651 12841
rect 23063 12804 23980 12832
rect 23063 12801 23075 12804
rect 23017 12795 23075 12801
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 9490 12764 9496 12776
rect 1903 12736 9496 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 13538 12764 13544 12776
rect 12492 12736 13544 12764
rect 12492 12724 12498 12736
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14550 12724 14556 12776
rect 14608 12724 14614 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15470 12764 15476 12776
rect 14875 12736 15476 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 15749 12767 15807 12773
rect 15749 12733 15761 12767
rect 15795 12764 15807 12767
rect 16114 12764 16120 12776
rect 15795 12736 16120 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12764 17463 12767
rect 19518 12764 19524 12776
rect 17451 12736 19524 12764
rect 17451 12733 17463 12736
rect 17405 12727 17463 12733
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 19702 12724 19708 12776
rect 19760 12724 19766 12776
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20162 12764 20168 12776
rect 19935 12736 20168 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20162 12724 20168 12736
rect 20220 12724 20226 12776
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 20496 12736 21281 12764
rect 20496 12724 20502 12736
rect 21269 12733 21281 12736
rect 21315 12733 21327 12767
rect 21269 12727 21327 12733
rect 22002 12724 22008 12776
rect 22060 12724 22066 12776
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 22741 12767 22799 12773
rect 22741 12764 22753 12767
rect 22152 12736 22753 12764
rect 22152 12724 22158 12736
rect 22741 12733 22753 12736
rect 22787 12764 22799 12767
rect 22787 12736 23520 12764
rect 22787 12733 22799 12736
rect 22741 12727 22799 12733
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 12894 12696 12900 12708
rect 12768 12668 12900 12696
rect 12768 12656 12774 12668
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 15286 12656 15292 12708
rect 15344 12696 15350 12708
rect 15838 12696 15844 12708
rect 15344 12668 15844 12696
rect 15344 12656 15350 12668
rect 15838 12656 15844 12668
rect 15896 12656 15902 12708
rect 16669 12699 16727 12705
rect 16669 12696 16681 12699
rect 15948 12668 16681 12696
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11241 12631 11299 12637
rect 11241 12628 11253 12631
rect 11204 12600 11253 12628
rect 11204 12588 11210 12600
rect 11241 12597 11253 12600
rect 11287 12597 11299 12631
rect 11241 12591 11299 12597
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 12526 12628 12532 12640
rect 12483 12600 12532 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 15562 12628 15568 12640
rect 12676 12600 15568 12628
rect 12676 12588 12682 12600
rect 15562 12588 15568 12600
rect 15620 12628 15626 12640
rect 15948 12628 15976 12668
rect 16669 12665 16681 12668
rect 16715 12696 16727 12699
rect 17126 12696 17132 12708
rect 16715 12668 17132 12696
rect 16715 12665 16727 12668
rect 16669 12659 16727 12665
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 19245 12699 19303 12705
rect 19245 12696 19257 12699
rect 17828 12668 19257 12696
rect 17828 12656 17834 12668
rect 19245 12665 19257 12668
rect 19291 12665 19303 12699
rect 19245 12659 19303 12665
rect 20364 12668 21220 12696
rect 15620 12600 15976 12628
rect 15620 12588 15626 12600
rect 16298 12588 16304 12640
rect 16356 12588 16362 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20364 12637 20392 12668
rect 20349 12631 20407 12637
rect 20349 12628 20361 12631
rect 19392 12600 20361 12628
rect 19392 12588 19398 12600
rect 20349 12597 20361 12600
rect 20395 12597 20407 12631
rect 21192 12628 21220 12668
rect 21542 12656 21548 12708
rect 21600 12696 21606 12708
rect 22922 12696 22928 12708
rect 21600 12668 22928 12696
rect 21600 12656 21606 12668
rect 22922 12656 22928 12668
rect 22980 12656 22986 12708
rect 23382 12656 23388 12708
rect 23440 12656 23446 12708
rect 23492 12696 23520 12736
rect 23566 12724 23572 12776
rect 23624 12764 23630 12776
rect 23842 12764 23848 12776
rect 23624 12736 23848 12764
rect 23624 12724 23630 12736
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 23952 12764 23980 12804
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 29181 12835 29239 12841
rect 29181 12801 29193 12835
rect 29227 12832 29239 12835
rect 30006 12832 30012 12844
rect 29227 12804 30012 12832
rect 29227 12801 29239 12804
rect 29181 12795 29239 12801
rect 30006 12792 30012 12804
rect 30064 12792 30070 12844
rect 31846 12832 31852 12844
rect 31418 12804 31852 12832
rect 31846 12792 31852 12804
rect 31904 12792 31910 12844
rect 32122 12792 32128 12844
rect 32180 12832 32186 12844
rect 32585 12835 32643 12841
rect 32585 12832 32597 12835
rect 32180 12804 32597 12832
rect 32180 12792 32186 12804
rect 32585 12801 32597 12804
rect 32631 12801 32643 12835
rect 32585 12795 32643 12801
rect 34057 12835 34115 12841
rect 34057 12801 34069 12835
rect 34103 12832 34115 12835
rect 34422 12832 34428 12844
rect 34103 12804 34428 12832
rect 34103 12801 34115 12804
rect 34057 12795 34115 12801
rect 34422 12792 34428 12804
rect 34480 12792 34486 12844
rect 35912 12832 35940 12872
rect 36078 12860 36084 12912
rect 36136 12900 36142 12912
rect 36538 12900 36544 12912
rect 36136 12872 36544 12900
rect 36136 12860 36142 12872
rect 36538 12860 36544 12872
rect 36596 12860 36602 12912
rect 36906 12860 36912 12912
rect 36964 12900 36970 12912
rect 37642 12900 37648 12912
rect 36964 12872 37648 12900
rect 36964 12860 36970 12872
rect 37642 12860 37648 12872
rect 37700 12860 37706 12912
rect 36633 12835 36691 12841
rect 36633 12832 36645 12835
rect 35912 12804 36645 12832
rect 36633 12801 36645 12804
rect 36679 12832 36691 12835
rect 36814 12832 36820 12844
rect 36679 12804 36820 12832
rect 36679 12801 36691 12804
rect 36633 12795 36691 12801
rect 36814 12792 36820 12804
rect 36872 12792 36878 12844
rect 37458 12792 37464 12844
rect 37516 12792 37522 12844
rect 38838 12792 38844 12844
rect 38896 12792 38902 12844
rect 40034 12792 40040 12844
rect 40092 12832 40098 12844
rect 40497 12835 40555 12841
rect 40497 12832 40509 12835
rect 40092 12804 40509 12832
rect 40092 12792 40098 12804
rect 40497 12801 40509 12804
rect 40543 12801 40555 12835
rect 40497 12795 40555 12801
rect 45922 12792 45928 12844
rect 45980 12792 45986 12844
rect 47854 12792 47860 12844
rect 47912 12832 47918 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47912 12804 47961 12832
rect 47912 12792 47918 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 49142 12792 49148 12844
rect 49200 12792 49206 12844
rect 25869 12767 25927 12773
rect 25869 12764 25881 12767
rect 23952 12736 25881 12764
rect 25869 12733 25881 12736
rect 25915 12764 25927 12767
rect 26050 12764 26056 12776
rect 25915 12736 26056 12764
rect 25915 12733 25927 12736
rect 25869 12727 25927 12733
rect 26050 12724 26056 12736
rect 26108 12724 26114 12776
rect 26786 12764 26792 12776
rect 26436 12736 26792 12764
rect 23492 12668 24348 12696
rect 21266 12628 21272 12640
rect 21192 12600 21272 12628
rect 20349 12591 20407 12597
rect 21266 12588 21272 12600
rect 21324 12628 21330 12640
rect 24026 12628 24032 12640
rect 21324 12600 24032 12628
rect 21324 12588 21330 12600
rect 24026 12588 24032 12600
rect 24084 12588 24090 12640
rect 24320 12628 24348 12668
rect 26436 12637 26464 12736
rect 26786 12724 26792 12736
rect 26844 12764 26850 12776
rect 27157 12767 27215 12773
rect 27157 12764 27169 12767
rect 26844 12736 27169 12764
rect 26844 12724 26850 12736
rect 27157 12733 27169 12736
rect 27203 12733 27215 12767
rect 27157 12727 27215 12733
rect 28902 12724 28908 12776
rect 28960 12764 28966 12776
rect 32401 12767 32459 12773
rect 32401 12764 32413 12767
rect 28960 12736 32413 12764
rect 28960 12724 28966 12736
rect 32401 12733 32413 12736
rect 32447 12733 32459 12767
rect 33870 12764 33876 12776
rect 32401 12727 32459 12733
rect 32968 12736 33876 12764
rect 32968 12696 32996 12736
rect 33870 12724 33876 12736
rect 33928 12724 33934 12776
rect 34790 12724 34796 12776
rect 34848 12764 34854 12776
rect 35529 12767 35587 12773
rect 35529 12764 35541 12767
rect 34848 12736 35541 12764
rect 34848 12724 34854 12736
rect 35529 12733 35541 12736
rect 35575 12733 35587 12767
rect 35529 12727 35587 12733
rect 35713 12767 35771 12773
rect 35713 12733 35725 12767
rect 35759 12764 35771 12767
rect 36998 12764 37004 12776
rect 35759 12736 37004 12764
rect 35759 12733 35771 12736
rect 35713 12727 35771 12733
rect 31726 12668 32996 12696
rect 33045 12699 33103 12705
rect 26421 12631 26479 12637
rect 26421 12628 26433 12631
rect 24320 12600 26433 12628
rect 26421 12597 26433 12600
rect 26467 12597 26479 12631
rect 26421 12591 26479 12597
rect 27798 12588 27804 12640
rect 27856 12628 27862 12640
rect 31726 12628 31754 12668
rect 33045 12665 33057 12699
rect 33091 12696 33103 12699
rect 34514 12696 34520 12708
rect 33091 12668 34520 12696
rect 33091 12665 33103 12668
rect 33045 12659 33103 12665
rect 34514 12656 34520 12668
rect 34572 12656 34578 12708
rect 27856 12600 31754 12628
rect 27856 12588 27862 12600
rect 33318 12588 33324 12640
rect 33376 12628 33382 12640
rect 33597 12631 33655 12637
rect 33597 12628 33609 12631
rect 33376 12600 33609 12628
rect 33376 12588 33382 12600
rect 33597 12597 33609 12600
rect 33643 12628 33655 12631
rect 33781 12631 33839 12637
rect 33781 12628 33793 12631
rect 33643 12600 33793 12628
rect 33643 12597 33655 12600
rect 33597 12591 33655 12597
rect 33781 12597 33793 12600
rect 33827 12628 33839 12631
rect 34238 12628 34244 12640
rect 33827 12600 34244 12628
rect 33827 12597 33839 12600
rect 33781 12591 33839 12597
rect 34238 12588 34244 12600
rect 34296 12628 34302 12640
rect 35434 12628 35440 12640
rect 34296 12600 35440 12628
rect 34296 12588 34302 12600
rect 35434 12588 35440 12600
rect 35492 12588 35498 12640
rect 35544 12628 35572 12727
rect 36998 12724 37004 12736
rect 37056 12724 37062 12776
rect 37737 12767 37795 12773
rect 37737 12733 37749 12767
rect 37783 12764 37795 12767
rect 38286 12764 38292 12776
rect 37783 12736 38292 12764
rect 37783 12733 37795 12736
rect 37737 12727 37795 12733
rect 38286 12724 38292 12736
rect 38344 12724 38350 12776
rect 39298 12724 39304 12776
rect 39356 12764 39362 12776
rect 39485 12767 39543 12773
rect 39485 12764 39497 12767
rect 39356 12736 39497 12764
rect 39356 12724 39362 12736
rect 39485 12733 39497 12736
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 36173 12699 36231 12705
rect 36173 12665 36185 12699
rect 36219 12696 36231 12699
rect 40221 12699 40279 12705
rect 36219 12668 37596 12696
rect 36219 12665 36231 12668
rect 36173 12659 36231 12665
rect 36817 12631 36875 12637
rect 36817 12628 36829 12631
rect 35544 12600 36829 12628
rect 36817 12597 36829 12600
rect 36863 12628 36875 12631
rect 36906 12628 36912 12640
rect 36863 12600 36912 12628
rect 36863 12597 36875 12600
rect 36817 12591 36875 12597
rect 36906 12588 36912 12600
rect 36964 12588 36970 12640
rect 36998 12588 37004 12640
rect 37056 12588 37062 12640
rect 37568 12628 37596 12668
rect 40221 12665 40233 12699
rect 40267 12696 40279 12699
rect 46750 12696 46756 12708
rect 40267 12668 46756 12696
rect 40267 12665 40279 12668
rect 40221 12659 40279 12665
rect 46750 12656 46756 12668
rect 46808 12656 46814 12708
rect 39114 12628 39120 12640
rect 37568 12600 39120 12628
rect 39114 12588 39120 12600
rect 39172 12588 39178 12640
rect 46109 12631 46167 12637
rect 46109 12597 46121 12631
rect 46155 12628 46167 12631
rect 47946 12628 47952 12640
rect 46155 12600 47952 12628
rect 46155 12597 46167 12600
rect 46109 12591 46167 12597
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11790 12424 11796 12436
rect 11287 12396 11796 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 12032 12396 16405 12424
rect 12032 12384 12038 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 16393 12387 16451 12393
rect 1302 12248 1308 12300
rect 1360 12288 1366 12300
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 1360 12260 2421 12288
rect 1360 12248 1366 12260
rect 2409 12257 2421 12260
rect 2455 12288 2467 12291
rect 2685 12291 2743 12297
rect 2685 12288 2697 12291
rect 2455 12260 2697 12288
rect 2455 12257 2467 12260
rect 2409 12251 2467 12257
rect 2685 12257 2697 12260
rect 2731 12257 2743 12291
rect 2685 12251 2743 12257
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 10778 12288 10784 12300
rect 9539 12260 10784 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 10778 12248 10784 12260
rect 10836 12288 10842 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 10836 12260 11713 12288
rect 10836 12248 10842 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 13725 12291 13783 12297
rect 12400 12260 13124 12288
rect 12400 12248 12406 12260
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 5810 12220 5816 12232
rect 2179 12192 5816 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 10870 12180 10876 12232
rect 10928 12180 10934 12232
rect 13096 12220 13124 12260
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 14826 12288 14832 12300
rect 13771 12260 14832 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15746 12288 15752 12300
rect 15528 12260 15752 12288
rect 15528 12248 15534 12260
rect 15746 12248 15752 12260
rect 15804 12288 15810 12300
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 15804 12260 16129 12288
rect 15804 12248 15810 12260
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 14734 12220 14740 12232
rect 13096 12206 14740 12220
rect 13110 12192 14740 12206
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 16408 12220 16436 12387
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 16724 12396 19441 12424
rect 16724 12384 16730 12396
rect 19429 12393 19441 12396
rect 19475 12393 19487 12427
rect 21542 12424 21548 12436
rect 19429 12387 19487 12393
rect 19536 12396 21548 12424
rect 19536 12356 19564 12396
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 21637 12427 21695 12433
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 21683 12396 22416 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 17144 12328 19564 12356
rect 22388 12356 22416 12396
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 23293 12427 23351 12433
rect 23293 12424 23305 12427
rect 22520 12396 23305 12424
rect 22520 12384 22526 12396
rect 23293 12393 23305 12396
rect 23339 12393 23351 12427
rect 26694 12424 26700 12436
rect 23293 12387 23351 12393
rect 23860 12396 26700 12424
rect 23474 12356 23480 12368
rect 22388 12328 23480 12356
rect 17144 12229 17172 12328
rect 23474 12316 23480 12328
rect 23532 12316 23538 12368
rect 17402 12248 17408 12300
rect 17460 12248 17466 12300
rect 17512 12260 19472 12288
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16408 12192 17141 12220
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17512 12220 17540 12260
rect 17276 12192 17540 12220
rect 17276 12180 17282 12192
rect 9766 12112 9772 12164
rect 9824 12112 9830 12164
rect 11054 12112 11060 12164
rect 11112 12152 11118 12164
rect 11977 12155 12035 12161
rect 11977 12152 11989 12155
rect 11112 12124 11989 12152
rect 11112 12112 11118 12124
rect 11977 12121 11989 12124
rect 12023 12121 12035 12155
rect 11977 12115 12035 12121
rect 13446 12112 13452 12164
rect 13504 12152 13510 12164
rect 13504 12124 14504 12152
rect 13504 12112 13510 12124
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 14240 12056 14381 12084
rect 14240 12044 14246 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14476 12084 14504 12124
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 15841 12155 15899 12161
rect 15841 12152 15853 12155
rect 15620 12124 15853 12152
rect 15620 12112 15626 12124
rect 15841 12121 15853 12124
rect 15887 12121 15899 12155
rect 15841 12115 15899 12121
rect 18141 12155 18199 12161
rect 18141 12121 18153 12155
rect 18187 12152 18199 12155
rect 18598 12152 18604 12164
rect 18187 12124 18604 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 18874 12112 18880 12164
rect 18932 12152 18938 12164
rect 19242 12152 19248 12164
rect 18932 12124 19248 12152
rect 18932 12112 18938 12124
rect 19242 12112 19248 12124
rect 19300 12112 19306 12164
rect 19444 12152 19472 12260
rect 19886 12248 19892 12300
rect 19944 12288 19950 12300
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19944 12260 19993 12288
rect 19944 12248 19950 12260
rect 19981 12257 19993 12260
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20625 12291 20683 12297
rect 20625 12257 20637 12291
rect 20671 12288 20683 12291
rect 21085 12291 21143 12297
rect 21085 12288 21097 12291
rect 20671 12260 21097 12288
rect 20671 12257 20683 12260
rect 20625 12251 20683 12257
rect 21085 12257 21097 12260
rect 21131 12288 21143 12291
rect 22094 12288 22100 12300
rect 21131 12260 22100 12288
rect 21131 12257 21143 12260
rect 21085 12251 21143 12257
rect 22094 12248 22100 12260
rect 22152 12248 22158 12300
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12288 22339 12291
rect 23753 12291 23811 12297
rect 22327 12260 23704 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 19576 12192 19809 12220
rect 19576 12180 19582 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 20990 12180 20996 12232
rect 21048 12220 21054 12232
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 21048 12192 21189 12220
rect 21048 12180 21054 12192
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 21726 12220 21732 12232
rect 21315 12192 21732 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21726 12180 21732 12192
rect 21784 12180 21790 12232
rect 23676 12220 23704 12260
rect 23753 12257 23765 12291
rect 23799 12288 23811 12291
rect 23860 12288 23888 12396
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 27709 12427 27767 12433
rect 27709 12393 27721 12427
rect 27755 12424 27767 12427
rect 27890 12424 27896 12436
rect 27755 12396 27896 12424
rect 27755 12393 27767 12396
rect 27709 12387 27767 12393
rect 27890 12384 27896 12396
rect 27948 12384 27954 12436
rect 31846 12384 31852 12436
rect 31904 12384 31910 12436
rect 33870 12384 33876 12436
rect 33928 12424 33934 12436
rect 33928 12396 37228 12424
rect 33928 12384 33934 12396
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 27338 12356 27344 12368
rect 26384 12328 27344 12356
rect 26384 12316 26390 12328
rect 27338 12316 27344 12328
rect 27396 12316 27402 12368
rect 34238 12316 34244 12368
rect 34296 12316 34302 12368
rect 23799 12260 23888 12288
rect 23937 12291 23995 12297
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 23937 12257 23949 12291
rect 23983 12288 23995 12291
rect 24854 12288 24860 12300
rect 23983 12260 24860 12288
rect 23983 12257 23995 12260
rect 23937 12251 23995 12257
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 26878 12248 26884 12300
rect 26936 12288 26942 12300
rect 27062 12288 27068 12300
rect 26936 12260 27068 12288
rect 26936 12248 26942 12260
rect 27062 12248 27068 12260
rect 27120 12248 27126 12300
rect 28445 12291 28503 12297
rect 28445 12257 28457 12291
rect 28491 12288 28503 12291
rect 29733 12291 29791 12297
rect 29733 12288 29745 12291
rect 28491 12260 29745 12288
rect 28491 12257 28503 12260
rect 28445 12251 28503 12257
rect 29733 12257 29745 12260
rect 29779 12288 29791 12291
rect 30006 12288 30012 12300
rect 29779 12260 30012 12288
rect 29779 12257 29791 12260
rect 29733 12251 29791 12257
rect 30006 12248 30012 12260
rect 30064 12248 30070 12300
rect 32398 12248 32404 12300
rect 32456 12248 32462 12300
rect 23676 12192 23796 12220
rect 19444 12124 20760 12152
rect 16666 12084 16672 12096
rect 14476 12056 16672 12084
rect 14369 12047 14427 12053
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 16758 12044 16764 12096
rect 16816 12044 16822 12096
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 20622 12084 20628 12096
rect 19935 12056 20628 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 20732 12084 20760 12124
rect 22370 12112 22376 12164
rect 22428 12112 22434 12164
rect 22462 12112 22468 12164
rect 22520 12112 22526 12164
rect 23661 12155 23719 12161
rect 23661 12152 23673 12155
rect 22848 12124 23673 12152
rect 22388 12084 22416 12112
rect 22848 12093 22876 12124
rect 23661 12121 23673 12124
rect 23707 12121 23719 12155
rect 23661 12115 23719 12121
rect 20732 12056 22416 12084
rect 22833 12087 22891 12093
rect 22833 12053 22845 12087
rect 22879 12053 22891 12087
rect 23768 12084 23796 12192
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 25866 12180 25872 12232
rect 25924 12220 25930 12232
rect 26697 12223 26755 12229
rect 26697 12220 26709 12223
rect 25924 12192 26709 12220
rect 25924 12180 25930 12192
rect 26697 12189 26709 12192
rect 26743 12220 26755 12223
rect 27522 12220 27528 12232
rect 26743 12192 27528 12220
rect 26743 12189 26755 12192
rect 26697 12183 26755 12189
rect 27522 12180 27528 12192
rect 27580 12180 27586 12232
rect 32122 12180 32128 12232
rect 32180 12180 32186 12232
rect 33502 12180 33508 12232
rect 33560 12220 33566 12232
rect 34256 12220 34284 12316
rect 34790 12248 34796 12300
rect 34848 12288 34854 12300
rect 37200 12297 37228 12396
rect 38838 12384 38844 12436
rect 38896 12424 38902 12436
rect 38896 12396 39160 12424
rect 38896 12384 38902 12396
rect 39025 12359 39083 12365
rect 39025 12325 39037 12359
rect 39071 12325 39083 12359
rect 39132 12356 39160 12396
rect 39298 12384 39304 12436
rect 39356 12384 39362 12436
rect 39485 12359 39543 12365
rect 39485 12356 39497 12359
rect 39132 12328 39497 12356
rect 39025 12319 39083 12325
rect 39485 12325 39497 12328
rect 39531 12325 39543 12359
rect 39485 12319 39543 12325
rect 40313 12359 40371 12365
rect 40313 12325 40325 12359
rect 40359 12356 40371 12359
rect 47210 12356 47216 12368
rect 40359 12328 47216 12356
rect 40359 12325 40371 12328
rect 40313 12319 40371 12325
rect 35161 12291 35219 12297
rect 35161 12288 35173 12291
rect 34848 12260 35173 12288
rect 34848 12248 34854 12260
rect 35161 12257 35173 12260
rect 35207 12257 35219 12291
rect 35161 12251 35219 12257
rect 37185 12291 37243 12297
rect 37185 12257 37197 12291
rect 37231 12257 37243 12291
rect 37185 12251 37243 12257
rect 37366 12248 37372 12300
rect 37424 12248 37430 12300
rect 38378 12248 38384 12300
rect 38436 12248 38442 12300
rect 38565 12291 38623 12297
rect 38565 12257 38577 12291
rect 38611 12288 38623 12291
rect 38746 12288 38752 12300
rect 38611 12260 38752 12288
rect 38611 12257 38623 12260
rect 38565 12251 38623 12257
rect 38746 12248 38752 12260
rect 38804 12248 38810 12300
rect 39040 12288 39068 12319
rect 47210 12316 47216 12328
rect 47268 12316 47274 12368
rect 39040 12260 41460 12288
rect 33560 12192 34284 12220
rect 33560 12180 33566 12192
rect 34882 12180 34888 12232
rect 34940 12180 34946 12232
rect 41432 12229 41460 12260
rect 49142 12248 49148 12300
rect 49200 12248 49206 12300
rect 40773 12223 40831 12229
rect 40773 12220 40785 12223
rect 37844 12192 40785 12220
rect 23842 12112 23848 12164
rect 23900 12152 23906 12164
rect 24857 12155 24915 12161
rect 24857 12152 24869 12155
rect 23900 12124 24869 12152
rect 23900 12112 23906 12124
rect 24857 12121 24869 12124
rect 24903 12121 24915 12155
rect 24857 12115 24915 12121
rect 28810 12112 28816 12164
rect 28868 12152 28874 12164
rect 29181 12155 29239 12161
rect 29181 12152 29193 12155
rect 28868 12124 29193 12152
rect 28868 12112 28874 12124
rect 29181 12121 29193 12124
rect 29227 12121 29239 12155
rect 29181 12115 29239 12121
rect 29914 12112 29920 12164
rect 29972 12152 29978 12164
rect 30009 12155 30067 12161
rect 30009 12152 30021 12155
rect 29972 12124 30021 12152
rect 29972 12112 29978 12124
rect 30009 12121 30021 12124
rect 30055 12121 30067 12155
rect 31846 12152 31852 12164
rect 31234 12124 31852 12152
rect 30009 12115 30067 12121
rect 31846 12112 31852 12124
rect 31904 12112 31910 12164
rect 35434 12112 35440 12164
rect 35492 12152 35498 12164
rect 35492 12124 35650 12152
rect 35492 12112 35498 12124
rect 24210 12084 24216 12096
rect 23768 12056 24216 12084
rect 22833 12047 22891 12053
rect 24210 12044 24216 12056
rect 24268 12084 24274 12096
rect 26326 12084 26332 12096
rect 24268 12056 26332 12084
rect 24268 12044 24274 12056
rect 26326 12044 26332 12056
rect 26384 12044 26390 12096
rect 26970 12044 26976 12096
rect 27028 12084 27034 12096
rect 27246 12084 27252 12096
rect 27028 12056 27252 12084
rect 27028 12044 27034 12056
rect 27246 12044 27252 12056
rect 27304 12044 27310 12096
rect 27338 12044 27344 12096
rect 27396 12044 27402 12096
rect 31386 12044 31392 12096
rect 31444 12084 31450 12096
rect 31481 12087 31539 12093
rect 31481 12084 31493 12087
rect 31444 12056 31493 12084
rect 31444 12044 31450 12056
rect 31481 12053 31493 12056
rect 31527 12053 31539 12087
rect 31481 12047 31539 12053
rect 34330 12044 34336 12096
rect 34388 12044 34394 12096
rect 36633 12087 36691 12093
rect 36633 12053 36645 12087
rect 36679 12084 36691 12087
rect 36722 12084 36728 12096
rect 36679 12056 36728 12084
rect 36679 12053 36691 12056
rect 36633 12047 36691 12053
rect 36722 12044 36728 12056
rect 36780 12044 36786 12096
rect 37461 12087 37519 12093
rect 37461 12053 37473 12087
rect 37507 12084 37519 12087
rect 37550 12084 37556 12096
rect 37507 12056 37556 12084
rect 37507 12053 37519 12056
rect 37461 12047 37519 12053
rect 37550 12044 37556 12056
rect 37608 12044 37614 12096
rect 37844 12093 37872 12192
rect 40773 12189 40785 12192
rect 40819 12189 40831 12223
rect 40773 12183 40831 12189
rect 41417 12223 41475 12229
rect 41417 12189 41429 12223
rect 41463 12189 41475 12223
rect 45925 12223 45983 12229
rect 45925 12220 45937 12223
rect 41417 12183 41475 12189
rect 45526 12192 45937 12220
rect 40129 12155 40187 12161
rect 40129 12121 40141 12155
rect 40175 12152 40187 12155
rect 40402 12152 40408 12164
rect 40175 12124 40408 12152
rect 40175 12121 40187 12124
rect 40129 12115 40187 12121
rect 40402 12112 40408 12124
rect 40460 12112 40466 12164
rect 37829 12087 37887 12093
rect 37829 12053 37841 12087
rect 37875 12053 37887 12087
rect 37829 12047 37887 12053
rect 38654 12044 38660 12096
rect 38712 12044 38718 12096
rect 40954 12044 40960 12096
rect 41012 12044 41018 12096
rect 41601 12087 41659 12093
rect 41601 12053 41613 12087
rect 41647 12084 41659 12087
rect 45526 12084 45554 12192
rect 45925 12189 45937 12192
rect 45971 12189 45983 12223
rect 45925 12183 45983 12189
rect 47946 12180 47952 12232
rect 48004 12180 48010 12232
rect 41647 12056 45554 12084
rect 41647 12053 41659 12056
rect 41601 12047 41659 12053
rect 46106 12044 46112 12096
rect 46164 12044 46170 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 4246 11880 4252 11892
rect 2547 11852 4252 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11609 11883 11667 11889
rect 11609 11880 11621 11883
rect 10928 11852 11621 11880
rect 10928 11840 10934 11852
rect 11609 11849 11621 11852
rect 11655 11880 11667 11883
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 11655 11852 12081 11880
rect 11655 11849 11667 11852
rect 11609 11843 11667 11849
rect 12069 11849 12081 11852
rect 12115 11880 12127 11883
rect 12342 11880 12348 11892
rect 12115 11852 12348 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12710 11840 12716 11892
rect 12768 11840 12774 11892
rect 13354 11840 13360 11892
rect 13412 11840 13418 11892
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 14185 11883 14243 11889
rect 14185 11880 14197 11883
rect 13688 11852 14197 11880
rect 13688 11840 13694 11852
rect 14185 11849 14197 11852
rect 14231 11849 14243 11883
rect 14185 11843 14243 11849
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 15194 11880 15200 11892
rect 14323 11852 15200 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15473 11883 15531 11889
rect 15473 11849 15485 11883
rect 15519 11880 15531 11883
rect 15838 11880 15844 11892
rect 15519 11852 15844 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 15838 11840 15844 11852
rect 15896 11880 15902 11892
rect 16390 11880 16396 11892
rect 15896 11852 16396 11880
rect 15896 11840 15902 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16485 11883 16543 11889
rect 16485 11849 16497 11883
rect 16531 11880 16543 11883
rect 17034 11880 17040 11892
rect 16531 11852 17040 11880
rect 16531 11849 16543 11852
rect 16485 11843 16543 11849
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 19242 11840 19248 11892
rect 19300 11880 19306 11892
rect 26605 11883 26663 11889
rect 19300 11852 22324 11880
rect 19300 11840 19306 11852
rect 2130 11772 2136 11824
rect 2188 11812 2194 11824
rect 13998 11812 14004 11824
rect 2188 11784 14004 11812
rect 2188 11772 2194 11784
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 17052 11812 17080 11840
rect 20346 11812 20352 11824
rect 14884 11784 15792 11812
rect 17052 11784 17158 11812
rect 19720 11784 20352 11812
rect 14884 11772 14890 11784
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1268 11716 1593 11744
rect 1268 11704 1274 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 2332 11676 2360 11707
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 13541 11747 13599 11753
rect 11848 11716 12940 11744
rect 11848 11704 11854 11716
rect 12912 11685 12940 11716
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 14734 11744 14740 11756
rect 13587 11716 14740 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 2777 11679 2835 11685
rect 2777 11676 2789 11679
rect 1360 11648 2789 11676
rect 1360 11636 1366 11648
rect 2777 11645 2789 11648
rect 2823 11645 2835 11679
rect 2777 11639 2835 11645
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 11422 11608 11428 11620
rect 1811 11580 11428 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 12250 11568 12256 11620
rect 12308 11608 12314 11620
rect 12710 11608 12716 11620
rect 12308 11580 12716 11608
rect 12308 11568 12314 11580
rect 12710 11568 12716 11580
rect 12768 11568 12774 11620
rect 12820 11608 12848 11639
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13630 11676 13636 11688
rect 13320 11648 13636 11676
rect 13320 11636 13326 11648
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13998 11636 14004 11688
rect 14056 11636 14062 11688
rect 15562 11636 15568 11688
rect 15620 11636 15626 11688
rect 15764 11685 15792 11784
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11744 19303 11747
rect 19334 11744 19340 11756
rect 19291 11716 19340 11744
rect 19291 11713 19303 11716
rect 19245 11707 19303 11713
rect 19334 11704 19340 11716
rect 19392 11704 19398 11756
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11645 15807 11679
rect 15749 11639 15807 11645
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 16172 11648 16865 11676
rect 16172 11636 16178 11648
rect 16853 11645 16865 11648
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11676 18383 11679
rect 18371 11648 18552 11676
rect 18371 11645 18383 11648
rect 18325 11639 18383 11645
rect 14366 11608 14372 11620
rect 12820 11580 14372 11608
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 14645 11611 14703 11617
rect 14645 11577 14657 11611
rect 14691 11608 14703 11611
rect 15470 11608 15476 11620
rect 14691 11580 15476 11608
rect 14691 11577 14703 11580
rect 14645 11571 14703 11577
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 16942 11608 16948 11620
rect 15580 11580 16948 11608
rect 12342 11500 12348 11552
rect 12400 11500 12406 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14884 11512 15117 11540
rect 14884 11500 14890 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15580 11540 15608 11580
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 15436 11512 15608 11540
rect 15436 11500 15442 11512
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16264 11512 16313 11540
rect 16264 11500 16270 11512
rect 16301 11509 16313 11512
rect 16347 11540 16359 11543
rect 17954 11540 17960 11552
rect 16347 11512 17960 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 17954 11500 17960 11512
rect 18012 11500 18018 11552
rect 18524 11540 18552 11648
rect 18598 11636 18604 11688
rect 18656 11676 18662 11688
rect 18874 11676 18880 11688
rect 18656 11648 18880 11676
rect 18656 11636 18662 11648
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 19720 11685 19748 11784
rect 20346 11772 20352 11784
rect 20404 11772 20410 11824
rect 20990 11772 20996 11824
rect 21048 11812 21054 11824
rect 21177 11815 21235 11821
rect 21177 11812 21189 11815
rect 21048 11784 21189 11812
rect 21048 11772 21054 11784
rect 21177 11781 21189 11784
rect 21223 11812 21235 11815
rect 21266 11812 21272 11824
rect 21223 11784 21272 11812
rect 21223 11781 21235 11784
rect 21177 11775 21235 11781
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11744 19947 11747
rect 20070 11744 20076 11756
rect 19935 11716 20076 11744
rect 19935 11713 19947 11716
rect 19889 11707 19947 11713
rect 20070 11704 20076 11716
rect 20128 11744 20134 11756
rect 20530 11744 20536 11756
rect 20128 11716 20536 11744
rect 20128 11704 20134 11716
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11744 21143 11747
rect 22002 11744 22008 11756
rect 21131 11716 22008 11744
rect 21131 11713 21143 11716
rect 21085 11707 21143 11713
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22296 11753 22324 11852
rect 26605 11849 26617 11883
rect 26651 11880 26663 11883
rect 27338 11880 27344 11892
rect 26651 11852 27344 11880
rect 26651 11849 26663 11852
rect 26605 11843 26663 11849
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 27893 11883 27951 11889
rect 27893 11849 27905 11883
rect 27939 11880 27951 11883
rect 28718 11880 28724 11892
rect 27939 11852 28724 11880
rect 27939 11849 27951 11852
rect 27893 11843 27951 11849
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 31481 11883 31539 11889
rect 31481 11849 31493 11883
rect 31527 11880 31539 11883
rect 31754 11880 31760 11892
rect 31527 11852 31760 11880
rect 31527 11849 31539 11852
rect 31481 11843 31539 11849
rect 31754 11840 31760 11852
rect 31812 11840 31818 11892
rect 31846 11840 31852 11892
rect 31904 11840 31910 11892
rect 31938 11840 31944 11892
rect 31996 11880 32002 11892
rect 32585 11883 32643 11889
rect 32585 11880 32597 11883
rect 31996 11852 32597 11880
rect 31996 11840 32002 11852
rect 32585 11849 32597 11852
rect 32631 11849 32643 11883
rect 32585 11843 32643 11849
rect 32677 11883 32735 11889
rect 32677 11849 32689 11883
rect 32723 11880 32735 11883
rect 32766 11880 32772 11892
rect 32723 11852 32772 11880
rect 32723 11849 32735 11852
rect 32677 11843 32735 11849
rect 32766 11840 32772 11852
rect 32824 11840 32830 11892
rect 34793 11883 34851 11889
rect 34793 11849 34805 11883
rect 34839 11880 34851 11883
rect 35434 11880 35440 11892
rect 34839 11852 35440 11880
rect 34839 11849 34851 11852
rect 34793 11843 34851 11849
rect 35434 11840 35440 11852
rect 35492 11880 35498 11892
rect 35492 11852 35664 11880
rect 35492 11840 35498 11852
rect 24210 11772 24216 11824
rect 24268 11772 24274 11824
rect 25866 11812 25872 11824
rect 25438 11784 25872 11812
rect 25866 11772 25872 11784
rect 25924 11772 25930 11824
rect 26142 11772 26148 11824
rect 26200 11812 26206 11824
rect 26970 11812 26976 11824
rect 26200 11784 26976 11812
rect 26200 11772 26206 11784
rect 26970 11772 26976 11784
rect 27028 11812 27034 11824
rect 27525 11815 27583 11821
rect 27525 11812 27537 11815
rect 27028 11784 27537 11812
rect 27028 11772 27034 11784
rect 27525 11781 27537 11784
rect 27571 11781 27583 11815
rect 27525 11775 27583 11781
rect 27614 11772 27620 11824
rect 27672 11812 27678 11824
rect 30009 11815 30067 11821
rect 27672 11784 28842 11812
rect 27672 11772 27678 11784
rect 30009 11781 30021 11815
rect 30055 11812 30067 11815
rect 31386 11812 31392 11824
rect 30055 11784 31392 11812
rect 30055 11781 30067 11784
rect 30009 11775 30067 11781
rect 31386 11772 31392 11784
rect 31444 11772 31450 11824
rect 31570 11772 31576 11824
rect 31628 11812 31634 11824
rect 35526 11812 35532 11824
rect 31628 11784 33732 11812
rect 31628 11772 31634 11784
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22554 11744 22560 11756
rect 22327 11716 22560 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 31110 11704 31116 11756
rect 31168 11704 31174 11756
rect 31404 11744 31432 11772
rect 33704 11744 33732 11784
rect 33980 11784 35532 11812
rect 33781 11747 33839 11753
rect 33781 11744 33793 11747
rect 31404 11716 33640 11744
rect 33704 11716 33793 11744
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11645 19763 11679
rect 19705 11639 19763 11645
rect 19797 11679 19855 11685
rect 19797 11645 19809 11679
rect 19843 11676 19855 11679
rect 19843 11648 20944 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 19061 11611 19119 11617
rect 19061 11577 19073 11611
rect 19107 11608 19119 11611
rect 19812 11608 19840 11639
rect 19107 11580 19840 11608
rect 19107 11577 19119 11580
rect 19061 11571 19119 11577
rect 20254 11568 20260 11620
rect 20312 11568 20318 11620
rect 20717 11611 20775 11617
rect 20717 11577 20729 11611
rect 20763 11608 20775 11611
rect 20806 11608 20812 11620
rect 20763 11580 20812 11608
rect 20763 11577 20775 11580
rect 20717 11571 20775 11577
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 20916 11608 20944 11648
rect 21358 11636 21364 11688
rect 21416 11636 21422 11688
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11676 22155 11679
rect 22370 11676 22376 11688
rect 22143 11648 22376 11676
rect 22143 11645 22155 11648
rect 22097 11639 22155 11645
rect 22370 11636 22376 11648
rect 22428 11636 22434 11688
rect 23385 11679 23443 11685
rect 23385 11645 23397 11679
rect 23431 11676 23443 11679
rect 23937 11679 23995 11685
rect 23937 11676 23949 11679
rect 23431 11648 23949 11676
rect 23431 11645 23443 11648
rect 23385 11639 23443 11645
rect 23937 11645 23949 11648
rect 23983 11645 23995 11679
rect 23937 11639 23995 11645
rect 22646 11608 22652 11620
rect 20916 11580 22652 11608
rect 22646 11568 22652 11580
rect 22704 11568 22710 11620
rect 20438 11540 20444 11552
rect 18524 11512 20444 11540
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 21634 11500 21640 11552
rect 21692 11540 21698 11552
rect 21913 11543 21971 11549
rect 21913 11540 21925 11543
rect 21692 11512 21925 11540
rect 21692 11500 21698 11512
rect 21913 11509 21925 11512
rect 21959 11540 21971 11543
rect 22002 11540 22008 11552
rect 21959 11512 22008 11540
rect 21959 11509 21971 11512
rect 21913 11503 21971 11509
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 23952 11540 23980 11639
rect 24854 11636 24860 11688
rect 24912 11676 24918 11688
rect 25685 11679 25743 11685
rect 25685 11676 25697 11679
rect 24912 11648 25697 11676
rect 24912 11636 24918 11648
rect 25685 11645 25697 11648
rect 25731 11645 25743 11679
rect 25685 11639 25743 11645
rect 27154 11636 27160 11688
rect 27212 11676 27218 11688
rect 27249 11679 27307 11685
rect 27249 11676 27261 11679
rect 27212 11648 27261 11676
rect 27212 11636 27218 11648
rect 27249 11645 27261 11648
rect 27295 11645 27307 11679
rect 27249 11639 27307 11645
rect 27430 11636 27436 11688
rect 27488 11636 27494 11688
rect 28537 11679 28595 11685
rect 28537 11645 28549 11679
rect 28583 11676 28595 11679
rect 29546 11676 29552 11688
rect 28583 11648 29552 11676
rect 28583 11645 28595 11648
rect 28537 11639 28595 11645
rect 27338 11568 27344 11620
rect 27396 11608 27402 11620
rect 28552 11608 28580 11639
rect 29546 11636 29552 11648
rect 29604 11636 29610 11688
rect 29638 11636 29644 11688
rect 29696 11676 29702 11688
rect 30285 11679 30343 11685
rect 30285 11676 30297 11679
rect 29696 11648 30297 11676
rect 29696 11636 29702 11648
rect 30285 11645 30297 11648
rect 30331 11645 30343 11679
rect 30285 11639 30343 11645
rect 30834 11636 30840 11688
rect 30892 11636 30898 11688
rect 31021 11679 31079 11685
rect 31021 11645 31033 11679
rect 31067 11676 31079 11679
rect 31938 11676 31944 11688
rect 31067 11648 31944 11676
rect 31067 11645 31079 11648
rect 31021 11639 31079 11645
rect 31938 11636 31944 11648
rect 31996 11636 32002 11688
rect 32493 11679 32551 11685
rect 32493 11645 32505 11679
rect 32539 11676 32551 11679
rect 32674 11676 32680 11688
rect 32539 11648 32680 11676
rect 32539 11645 32551 11648
rect 32493 11639 32551 11645
rect 32674 11636 32680 11648
rect 32732 11636 32738 11688
rect 33612 11685 33640 11716
rect 33781 11713 33793 11716
rect 33827 11713 33839 11747
rect 33781 11707 33839 11713
rect 33870 11704 33876 11756
rect 33928 11704 33934 11756
rect 33597 11679 33655 11685
rect 33597 11645 33609 11679
rect 33643 11645 33655 11679
rect 33597 11639 33655 11645
rect 27396 11580 28580 11608
rect 30392 11580 31524 11608
rect 27396 11568 27402 11580
rect 24578 11540 24584 11552
rect 23952 11512 24584 11540
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 29270 11500 29276 11552
rect 29328 11540 29334 11552
rect 30392 11540 30420 11580
rect 29328 11512 30420 11540
rect 29328 11500 29334 11512
rect 30466 11500 30472 11552
rect 30524 11540 30530 11552
rect 31386 11540 31392 11552
rect 30524 11512 31392 11540
rect 30524 11500 30530 11512
rect 31386 11500 31392 11512
rect 31444 11500 31450 11552
rect 31496 11540 31524 11580
rect 31570 11568 31576 11620
rect 31628 11608 31634 11620
rect 33980 11608 34008 11784
rect 35526 11772 35532 11784
rect 35584 11772 35590 11824
rect 35636 11812 35664 11852
rect 35802 11840 35808 11892
rect 35860 11880 35866 11892
rect 37737 11883 37795 11889
rect 37737 11880 37749 11883
rect 35860 11852 37749 11880
rect 35860 11840 35866 11852
rect 37737 11849 37749 11852
rect 37783 11849 37795 11883
rect 37737 11843 37795 11849
rect 38654 11840 38660 11892
rect 38712 11840 38718 11892
rect 39114 11840 39120 11892
rect 39172 11840 39178 11892
rect 35894 11812 35900 11824
rect 35636 11784 35900 11812
rect 35894 11772 35900 11784
rect 35952 11772 35958 11824
rect 37366 11772 37372 11824
rect 37424 11812 37430 11824
rect 39945 11815 40003 11821
rect 39945 11812 39957 11815
rect 37424 11784 39957 11812
rect 37424 11772 37430 11784
rect 39945 11781 39957 11784
rect 39991 11812 40003 11815
rect 40589 11815 40647 11821
rect 40589 11812 40601 11815
rect 39991 11784 40601 11812
rect 39991 11781 40003 11784
rect 39945 11775 40003 11781
rect 40589 11781 40601 11784
rect 40635 11781 40647 11815
rect 40589 11775 40647 11781
rect 40954 11772 40960 11824
rect 41012 11812 41018 11824
rect 45097 11815 45155 11821
rect 45097 11812 45109 11815
rect 41012 11784 45109 11812
rect 41012 11772 41018 11784
rect 45097 11781 45109 11784
rect 45143 11781 45155 11815
rect 45097 11775 45155 11781
rect 49142 11772 49148 11824
rect 49200 11772 49206 11824
rect 36814 11704 36820 11756
rect 36872 11744 36878 11756
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 36872 11716 37841 11744
rect 36872 11704 36878 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 39022 11704 39028 11756
rect 39080 11704 39086 11756
rect 40402 11704 40408 11756
rect 40460 11704 40466 11756
rect 46106 11704 46112 11756
rect 46164 11744 46170 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 46164 11716 47961 11744
rect 46164 11704 46170 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 34422 11636 34428 11688
rect 34480 11676 34486 11688
rect 34517 11679 34575 11685
rect 34517 11676 34529 11679
rect 34480 11648 34529 11676
rect 34480 11636 34486 11648
rect 34517 11645 34529 11648
rect 34563 11645 34575 11679
rect 34517 11639 34575 11645
rect 34882 11636 34888 11688
rect 34940 11676 34946 11688
rect 35161 11679 35219 11685
rect 35161 11676 35173 11679
rect 34940 11648 35173 11676
rect 34940 11636 34946 11648
rect 35161 11645 35173 11648
rect 35207 11645 35219 11679
rect 35161 11639 35219 11645
rect 35437 11679 35495 11685
rect 35437 11645 35449 11679
rect 35483 11676 35495 11679
rect 36170 11676 36176 11688
rect 35483 11648 36176 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 31628 11580 34008 11608
rect 34241 11611 34299 11617
rect 31628 11568 31634 11580
rect 34241 11577 34253 11611
rect 34287 11608 34299 11611
rect 35066 11608 35072 11620
rect 34287 11580 35072 11608
rect 34287 11577 34299 11580
rect 34241 11571 34299 11577
rect 35066 11568 35072 11580
rect 35124 11568 35130 11620
rect 32858 11540 32864 11552
rect 31496 11512 32864 11540
rect 32858 11500 32864 11512
rect 32916 11500 32922 11552
rect 33045 11543 33103 11549
rect 33045 11509 33057 11543
rect 33091 11540 33103 11543
rect 34606 11540 34612 11552
rect 33091 11512 34612 11540
rect 33091 11509 33103 11512
rect 33045 11503 33103 11509
rect 34606 11500 34612 11512
rect 34664 11500 34670 11552
rect 35176 11540 35204 11639
rect 36170 11636 36176 11648
rect 36228 11676 36234 11688
rect 36228 11648 36584 11676
rect 36228 11636 36234 11648
rect 36556 11608 36584 11648
rect 36630 11636 36636 11688
rect 36688 11676 36694 11688
rect 37553 11679 37611 11685
rect 37553 11676 37565 11679
rect 36688 11648 37565 11676
rect 36688 11636 36694 11648
rect 37553 11645 37565 11648
rect 37599 11645 37611 11679
rect 39209 11679 39267 11685
rect 39209 11676 39221 11679
rect 37553 11639 37611 11645
rect 37660 11648 39221 11676
rect 36909 11611 36967 11617
rect 36556 11580 36768 11608
rect 36740 11552 36768 11580
rect 36909 11577 36921 11611
rect 36955 11608 36967 11611
rect 37182 11608 37188 11620
rect 36955 11580 37188 11608
rect 36955 11577 36967 11580
rect 36909 11571 36967 11577
rect 37182 11568 37188 11580
rect 37240 11568 37246 11620
rect 35618 11540 35624 11552
rect 35176 11512 35624 11540
rect 35618 11500 35624 11512
rect 35676 11500 35682 11552
rect 35802 11500 35808 11552
rect 35860 11540 35866 11552
rect 35986 11540 35992 11552
rect 35860 11512 35992 11540
rect 35860 11500 35866 11512
rect 35986 11500 35992 11512
rect 36044 11500 36050 11552
rect 36722 11500 36728 11552
rect 36780 11540 36786 11552
rect 37660 11540 37688 11648
rect 39209 11645 39221 11648
rect 39255 11645 39267 11679
rect 39209 11639 39267 11645
rect 40129 11611 40187 11617
rect 40129 11577 40141 11611
rect 40175 11608 40187 11611
rect 45281 11611 45339 11617
rect 40175 11580 42840 11608
rect 40175 11577 40187 11580
rect 40129 11571 40187 11577
rect 36780 11512 37688 11540
rect 38197 11543 38255 11549
rect 36780 11500 36786 11512
rect 38197 11509 38209 11543
rect 38243 11540 38255 11543
rect 40218 11540 40224 11552
rect 38243 11512 40224 11540
rect 38243 11509 38255 11512
rect 38197 11503 38255 11509
rect 40218 11500 40224 11512
rect 40276 11500 40282 11552
rect 42812 11540 42840 11580
rect 45281 11577 45293 11611
rect 45327 11608 45339 11611
rect 46566 11608 46572 11620
rect 45327 11580 46572 11608
rect 45327 11577 45339 11580
rect 45281 11571 45339 11577
rect 46566 11568 46572 11580
rect 46624 11568 46630 11620
rect 47026 11540 47032 11552
rect 42812 11512 47032 11540
rect 47026 11500 47032 11512
rect 47084 11500 47090 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 1210 11296 1216 11348
rect 1268 11336 1274 11348
rect 2133 11339 2191 11345
rect 2133 11336 2145 11339
rect 1268 11308 2145 11336
rect 1268 11296 1274 11308
rect 2133 11305 2145 11308
rect 2179 11305 2191 11339
rect 2133 11299 2191 11305
rect 2746 11308 12664 11336
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11268 1823 11271
rect 2746 11268 2774 11308
rect 1811 11240 2774 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11054 11200 11060 11212
rect 11011 11172 11060 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11790 11160 11796 11212
rect 11848 11200 11854 11212
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 11848 11172 12449 11200
rect 11848 11160 11854 11172
rect 12437 11169 12449 11172
rect 12483 11169 12495 11203
rect 12636 11200 12664 11308
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 13964 11308 14381 11336
rect 13964 11296 13970 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 16114 11336 16120 11348
rect 14608 11308 16120 11336
rect 14608 11296 14614 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16301 11339 16359 11345
rect 16301 11305 16313 11339
rect 16347 11336 16359 11339
rect 16390 11336 16396 11348
rect 16347 11308 16396 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 17126 11336 17132 11348
rect 16908 11308 17132 11336
rect 16908 11296 16914 11308
rect 17126 11296 17132 11308
rect 17184 11336 17190 11348
rect 19061 11339 19119 11345
rect 17184 11308 18460 11336
rect 17184 11296 17190 11308
rect 12710 11228 12716 11280
rect 12768 11268 12774 11280
rect 16761 11271 16819 11277
rect 16761 11268 16773 11271
rect 12768 11240 16773 11268
rect 12768 11228 12774 11240
rect 16761 11237 16773 11240
rect 16807 11237 16819 11271
rect 17957 11271 18015 11277
rect 17957 11268 17969 11271
rect 16761 11231 16819 11237
rect 16868 11240 17969 11268
rect 14458 11200 14464 11212
rect 12636 11172 14464 11200
rect 12437 11163 12495 11169
rect 14458 11160 14464 11172
rect 14516 11160 14522 11212
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11200 15071 11203
rect 15286 11200 15292 11212
rect 15059 11172 15292 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15746 11160 15752 11212
rect 15804 11160 15810 11212
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 15930 11200 15936 11212
rect 15887 11172 15936 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 16868 11200 16896 11240
rect 17957 11237 17969 11240
rect 18003 11237 18015 11271
rect 18432 11268 18460 11308
rect 19061 11305 19073 11339
rect 19107 11336 19119 11339
rect 19242 11336 19248 11348
rect 19107 11308 19248 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19521 11339 19579 11345
rect 19521 11336 19533 11339
rect 19484 11308 19533 11336
rect 19484 11296 19490 11308
rect 19521 11305 19533 11308
rect 19567 11336 19579 11339
rect 20070 11336 20076 11348
rect 19567 11308 20076 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 20438 11296 20444 11348
rect 20496 11296 20502 11348
rect 21931 11339 21989 11345
rect 21931 11305 21943 11339
rect 21977 11336 21989 11339
rect 21977 11308 23244 11336
rect 21977 11305 21989 11308
rect 21931 11299 21989 11305
rect 19150 11268 19156 11280
rect 18432 11240 19156 11268
rect 17957 11231 18015 11237
rect 18524 11209 18552 11240
rect 19150 11228 19156 11240
rect 19208 11228 19214 11280
rect 23216 11268 23244 11308
rect 23290 11296 23296 11348
rect 23348 11296 23354 11348
rect 25222 11336 25228 11348
rect 24596 11308 25228 11336
rect 23750 11268 23756 11280
rect 23216 11240 23756 11268
rect 23750 11228 23756 11240
rect 23808 11228 23814 11280
rect 16172 11172 16896 11200
rect 17405 11203 17463 11209
rect 16172 11160 16178 11172
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 18509 11203 18567 11209
rect 17451 11172 18460 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 1636 11104 2329 11132
rect 1636 11092 1642 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 12710 11092 12716 11144
rect 12768 11092 12774 11144
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 17034 11132 17040 11144
rect 13771 11104 17040 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 17034 11092 17040 11104
rect 17092 11092 17098 11144
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11132 17279 11135
rect 18322 11132 18328 11144
rect 17267 11104 18328 11132
rect 17267 11101 17279 11104
rect 17221 11095 17279 11101
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 18432 11132 18460 11172
rect 18509 11169 18521 11203
rect 18555 11169 18567 11203
rect 18509 11163 18567 11169
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 23842 11200 23848 11212
rect 20364 11172 23848 11200
rect 19518 11132 19524 11144
rect 18432 11104 19524 11132
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 12006 11036 12572 11064
rect 12544 11008 12572 11036
rect 12894 11024 12900 11076
rect 12952 11064 12958 11076
rect 12989 11067 13047 11073
rect 12989 11064 13001 11067
rect 12952 11036 13001 11064
rect 12952 11024 12958 11036
rect 12989 11033 13001 11036
rect 13035 11064 13047 11067
rect 15562 11064 15568 11076
rect 13035 11036 15568 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 16574 11064 16580 11076
rect 15979 11036 16580 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 17129 11067 17187 11073
rect 17129 11033 17141 11067
rect 17175 11064 17187 11067
rect 17770 11064 17776 11076
rect 17175 11036 17776 11064
rect 17175 11033 17187 11036
rect 17129 11027 17187 11033
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 17954 11024 17960 11076
rect 18012 11064 18018 11076
rect 18506 11064 18512 11076
rect 18012 11036 18512 11064
rect 18012 11024 18018 11036
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 13265 10999 13323 11005
rect 13265 10996 13277 10999
rect 12584 10968 13277 10996
rect 12584 10956 12590 10968
rect 13265 10965 13277 10968
rect 13311 10996 13323 10999
rect 14642 10996 14648 11008
rect 13311 10968 14648 10996
rect 13311 10965 13323 10968
rect 13265 10959 13323 10965
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 14734 10956 14740 11008
rect 14792 10956 14798 11008
rect 18340 11005 18368 11036
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 18598 11024 18604 11076
rect 18656 11064 18662 11076
rect 20364 11064 20392 11172
rect 23842 11160 23848 11172
rect 23900 11160 23906 11212
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11200 23995 11203
rect 24596 11200 24624 11308
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 26602 11336 26608 11348
rect 26375 11308 26608 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 28810 11296 28816 11348
rect 28868 11336 28874 11348
rect 28997 11339 29055 11345
rect 28997 11336 29009 11339
rect 28868 11308 29009 11336
rect 28868 11296 28874 11308
rect 28997 11305 29009 11308
rect 29043 11336 29055 11339
rect 33318 11336 33324 11348
rect 29043 11308 33324 11336
rect 29043 11305 29055 11308
rect 28997 11299 29055 11305
rect 33318 11296 33324 11308
rect 33376 11336 33382 11348
rect 34422 11336 34428 11348
rect 33376 11308 34428 11336
rect 33376 11296 33382 11308
rect 34422 11296 34428 11308
rect 34480 11336 34486 11348
rect 34701 11339 34759 11345
rect 34701 11336 34713 11339
rect 34480 11308 34713 11336
rect 34480 11296 34486 11308
rect 34701 11305 34713 11308
rect 34747 11305 34759 11339
rect 34701 11299 34759 11305
rect 35066 11296 35072 11348
rect 35124 11336 35130 11348
rect 38381 11339 38439 11345
rect 35124 11308 38240 11336
rect 35124 11296 35130 11308
rect 28629 11271 28687 11277
rect 28629 11237 28641 11271
rect 28675 11268 28687 11271
rect 28902 11268 28908 11280
rect 28675 11240 28908 11268
rect 28675 11237 28687 11240
rect 28629 11231 28687 11237
rect 28902 11228 28908 11240
rect 28960 11228 28966 11280
rect 30466 11228 30472 11280
rect 30524 11228 30530 11280
rect 32674 11228 32680 11280
rect 32732 11268 32738 11280
rect 32861 11271 32919 11277
rect 32861 11268 32873 11271
rect 32732 11240 32873 11268
rect 32732 11228 32738 11240
rect 32861 11237 32873 11240
rect 32907 11237 32919 11271
rect 32861 11231 32919 11237
rect 32950 11228 32956 11280
rect 33008 11268 33014 11280
rect 33008 11240 35894 11268
rect 33008 11228 33014 11240
rect 23983 11172 24624 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24854 11160 24860 11212
rect 24912 11160 24918 11212
rect 29181 11203 29239 11209
rect 29181 11169 29193 11203
rect 29227 11200 29239 11203
rect 29273 11203 29331 11209
rect 29273 11200 29285 11203
rect 29227 11172 29285 11200
rect 29227 11169 29239 11172
rect 29181 11163 29239 11169
rect 29273 11169 29285 11172
rect 29319 11169 29331 11203
rect 29273 11163 29331 11169
rect 29917 11203 29975 11209
rect 29917 11169 29929 11203
rect 29963 11200 29975 11203
rect 31478 11200 31484 11212
rect 29963 11172 31484 11200
rect 29963 11169 29975 11172
rect 29917 11163 29975 11169
rect 20806 11092 20812 11144
rect 20864 11092 20870 11144
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11132 22247 11135
rect 24578 11132 24584 11144
rect 22235 11104 24584 11132
rect 22235 11101 22247 11104
rect 22189 11095 22247 11101
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 28902 11092 28908 11144
rect 28960 11132 28966 11144
rect 29196 11132 29224 11163
rect 31478 11160 31484 11172
rect 31536 11160 31542 11212
rect 32122 11160 32128 11212
rect 32180 11200 32186 11212
rect 34057 11203 34115 11209
rect 34057 11200 34069 11203
rect 32180 11172 34069 11200
rect 32180 11160 32186 11172
rect 34057 11169 34069 11172
rect 34103 11200 34115 11203
rect 34882 11200 34888 11212
rect 34103 11172 34888 11200
rect 34103 11169 34115 11172
rect 34057 11163 34115 11169
rect 34882 11160 34888 11172
rect 34940 11160 34946 11212
rect 35866 11200 35894 11240
rect 37366 11200 37372 11212
rect 35866 11172 37372 11200
rect 37366 11160 37372 11172
rect 37424 11160 37430 11212
rect 37458 11160 37464 11212
rect 37516 11200 37522 11212
rect 37737 11203 37795 11209
rect 37737 11200 37749 11203
rect 37516 11172 37749 11200
rect 37516 11160 37522 11172
rect 37737 11169 37749 11172
rect 37783 11169 37795 11203
rect 37737 11163 37795 11169
rect 28960 11104 29224 11132
rect 28960 11092 28966 11104
rect 29638 11092 29644 11144
rect 29696 11132 29702 11144
rect 31113 11135 31171 11141
rect 31113 11132 31125 11135
rect 29696 11104 31125 11132
rect 29696 11092 29702 11104
rect 31113 11101 31125 11104
rect 31159 11101 31171 11135
rect 33226 11132 33232 11144
rect 32522 11104 33232 11132
rect 31113 11095 31171 11101
rect 33226 11092 33232 11104
rect 33284 11092 33290 11144
rect 33318 11092 33324 11144
rect 33376 11092 33382 11144
rect 35894 11092 35900 11144
rect 35952 11132 35958 11144
rect 36446 11132 36452 11144
rect 35952 11104 36452 11132
rect 35952 11092 35958 11104
rect 36446 11092 36452 11104
rect 36504 11092 36510 11144
rect 38212 11141 38240 11308
rect 38381 11305 38393 11339
rect 38427 11336 38439 11339
rect 44358 11336 44364 11348
rect 38427 11308 44364 11336
rect 38427 11305 38439 11308
rect 38381 11299 38439 11305
rect 44358 11296 44364 11308
rect 44416 11296 44422 11348
rect 38749 11271 38807 11277
rect 38749 11237 38761 11271
rect 38795 11268 38807 11271
rect 38838 11268 38844 11280
rect 38795 11240 38844 11268
rect 38795 11237 38807 11240
rect 38749 11231 38807 11237
rect 38838 11228 38844 11240
rect 38896 11228 38902 11280
rect 39482 11228 39488 11280
rect 39540 11268 39546 11280
rect 39577 11271 39635 11277
rect 39577 11268 39589 11271
rect 39540 11240 39589 11268
rect 39540 11228 39546 11240
rect 39577 11237 39589 11240
rect 39623 11237 39635 11271
rect 39577 11231 39635 11237
rect 40957 11271 41015 11277
rect 40957 11237 40969 11271
rect 41003 11268 41015 11271
rect 41003 11240 45554 11268
rect 41003 11237 41015 11240
rect 40957 11231 41015 11237
rect 38197 11135 38255 11141
rect 38197 11101 38209 11135
rect 38243 11101 38255 11135
rect 39592 11132 39620 11231
rect 40129 11135 40187 11141
rect 40129 11132 40141 11135
rect 39592 11104 40141 11132
rect 38197 11095 38255 11101
rect 40129 11101 40141 11104
rect 40175 11101 40187 11135
rect 40129 11095 40187 11101
rect 40218 11092 40224 11144
rect 40276 11132 40282 11144
rect 40773 11135 40831 11141
rect 40773 11132 40785 11135
rect 40276 11104 40785 11132
rect 40276 11092 40282 11104
rect 40773 11101 40785 11104
rect 40819 11101 40831 11135
rect 45526 11132 45554 11240
rect 49142 11160 49148 11212
rect 49200 11160 49206 11212
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 45526 11104 45661 11132
rect 40773 11095 40831 11101
rect 45649 11101 45661 11104
rect 45695 11101 45707 11135
rect 45649 11095 45707 11101
rect 46750 11092 46756 11144
rect 46808 11132 46814 11144
rect 47949 11135 48007 11141
rect 47949 11132 47961 11135
rect 46808 11104 47961 11132
rect 46808 11092 46814 11104
rect 47949 11101 47961 11104
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 18656 11036 20392 11064
rect 18656 11024 18662 11036
rect 21634 11024 21640 11076
rect 21692 11064 21698 11076
rect 23661 11067 23719 11073
rect 21692 11036 22784 11064
rect 21692 11024 21698 11036
rect 18325 10999 18383 11005
rect 18325 10965 18337 10999
rect 18371 10965 18383 10999
rect 18325 10959 18383 10965
rect 18417 10999 18475 11005
rect 18417 10965 18429 10999
rect 18463 10996 18475 10999
rect 18616 10996 18644 11024
rect 18463 10968 18644 10996
rect 18463 10965 18475 10968
rect 18417 10959 18475 10965
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 22002 10996 22008 11008
rect 19484 10968 22008 10996
rect 19484 10956 19490 10968
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 22646 10956 22652 11008
rect 22704 10956 22710 11008
rect 22756 10996 22784 11036
rect 23661 11033 23673 11067
rect 23707 11064 23719 11067
rect 23934 11064 23940 11076
rect 23707 11036 23940 11064
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 25866 11024 25872 11076
rect 25924 11024 25930 11076
rect 27154 11024 27160 11076
rect 27212 11024 27218 11076
rect 27614 11024 27620 11076
rect 27672 11024 27678 11076
rect 29012 11036 29224 11064
rect 23566 10996 23572 11008
rect 22756 10968 23572 10996
rect 23566 10956 23572 10968
rect 23624 10956 23630 11008
rect 23753 10999 23811 11005
rect 23753 10965 23765 10999
rect 23799 10996 23811 10999
rect 23842 10996 23848 11008
rect 23799 10968 23848 10996
rect 23799 10965 23811 10968
rect 23753 10959 23811 10965
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 24486 10956 24492 11008
rect 24544 10996 24550 11008
rect 29012 10996 29040 11036
rect 24544 10968 29040 10996
rect 29196 10996 29224 11036
rect 29270 11024 29276 11076
rect 29328 11064 29334 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 29328 11036 30021 11064
rect 29328 11024 29334 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 31386 11024 31392 11076
rect 31444 11024 31450 11076
rect 31478 11024 31484 11076
rect 31536 11064 31542 11076
rect 35158 11064 35164 11076
rect 31536 11036 31754 11064
rect 31536 11024 31542 11036
rect 30101 10999 30159 11005
rect 30101 10996 30113 10999
rect 29196 10968 30113 10996
rect 24544 10956 24550 10968
rect 30101 10965 30113 10968
rect 30147 10996 30159 10999
rect 30742 10996 30748 11008
rect 30147 10968 30748 10996
rect 30147 10965 30159 10968
rect 30101 10959 30159 10965
rect 30742 10956 30748 10968
rect 30800 10956 30806 11008
rect 31726 10996 31754 11036
rect 32692 11036 35164 11064
rect 32692 10996 32720 11036
rect 35158 11024 35164 11036
rect 35216 11024 35222 11076
rect 35713 11067 35771 11073
rect 35713 11033 35725 11067
rect 35759 11064 35771 11067
rect 36078 11064 36084 11076
rect 35759 11036 36084 11064
rect 35759 11033 35771 11036
rect 35713 11027 35771 11033
rect 36078 11024 36084 11036
rect 36136 11024 36142 11076
rect 37182 11024 37188 11076
rect 37240 11064 37246 11076
rect 37461 11067 37519 11073
rect 37461 11064 37473 11067
rect 37240 11036 37473 11064
rect 37240 11024 37246 11036
rect 37461 11033 37473 11036
rect 37507 11064 37519 11067
rect 38378 11064 38384 11076
rect 37507 11036 38384 11064
rect 37507 11033 37519 11036
rect 37461 11027 37519 11033
rect 38378 11024 38384 11036
rect 38436 11024 38442 11076
rect 40313 11067 40371 11073
rect 40313 11033 40325 11067
rect 40359 11064 40371 11067
rect 45833 11067 45891 11073
rect 40359 11036 45554 11064
rect 40359 11033 40371 11036
rect 40313 11027 40371 11033
rect 31726 10968 32720 10996
rect 33686 10956 33692 11008
rect 33744 10996 33750 11008
rect 33962 10996 33968 11008
rect 33744 10968 33968 10996
rect 33744 10956 33750 10968
rect 33962 10956 33968 10968
rect 34020 10996 34026 11008
rect 38562 10996 38568 11008
rect 34020 10968 38568 10996
rect 34020 10956 34026 10968
rect 38562 10956 38568 10968
rect 38620 10956 38626 11008
rect 45526 10996 45554 11036
rect 45833 11033 45845 11067
rect 45879 11064 45891 11067
rect 46934 11064 46940 11076
rect 45879 11036 46940 11064
rect 45879 11033 45891 11036
rect 45833 11027 45891 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 46106 10996 46112 11008
rect 45526 10968 46112 10996
rect 46106 10956 46112 10968
rect 46164 10956 46170 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 1811 10764 2774 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 1210 10684 1216 10736
rect 1268 10724 1274 10736
rect 2746 10724 2774 10764
rect 12526 10752 12532 10804
rect 12584 10752 12590 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12860 10764 13185 10792
rect 12860 10752 12866 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 14366 10752 14372 10804
rect 14424 10752 14430 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 15979 10764 17141 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 19426 10792 19432 10804
rect 17644 10764 19432 10792
rect 17644 10752 17650 10764
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19702 10792 19708 10804
rect 19567 10764 19708 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 22646 10792 22652 10804
rect 21131 10764 22652 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 22922 10752 22928 10804
rect 22980 10792 22986 10804
rect 24213 10795 24271 10801
rect 24213 10792 24225 10795
rect 22980 10764 24225 10792
rect 22980 10752 22986 10764
rect 24213 10761 24225 10764
rect 24259 10761 24271 10795
rect 24213 10755 24271 10761
rect 25866 10752 25872 10804
rect 25924 10792 25930 10804
rect 26421 10795 26479 10801
rect 26421 10792 26433 10795
rect 25924 10764 26433 10792
rect 25924 10752 25930 10764
rect 26421 10761 26433 10764
rect 26467 10792 26479 10795
rect 26694 10792 26700 10804
rect 26467 10764 26700 10792
rect 26467 10761 26479 10764
rect 26421 10755 26479 10761
rect 26694 10752 26700 10764
rect 26752 10752 26758 10804
rect 27062 10752 27068 10804
rect 27120 10792 27126 10804
rect 30190 10792 30196 10804
rect 27120 10764 30196 10792
rect 27120 10752 27126 10764
rect 30190 10752 30196 10764
rect 30248 10792 30254 10804
rect 30834 10792 30840 10804
rect 30248 10764 30840 10792
rect 30248 10752 30254 10764
rect 30834 10752 30840 10764
rect 30892 10752 30898 10804
rect 31110 10752 31116 10804
rect 31168 10792 31174 10804
rect 31389 10795 31447 10801
rect 31389 10792 31401 10795
rect 31168 10764 31401 10792
rect 31168 10752 31174 10764
rect 31389 10761 31401 10764
rect 31435 10761 31447 10795
rect 31389 10755 31447 10761
rect 32306 10752 32312 10804
rect 32364 10792 32370 10804
rect 32490 10792 32496 10804
rect 32364 10764 32496 10792
rect 32364 10752 32370 10764
rect 32490 10752 32496 10764
rect 32548 10792 32554 10804
rect 33873 10795 33931 10801
rect 33873 10792 33885 10795
rect 32548 10764 33885 10792
rect 32548 10752 32554 10764
rect 33873 10761 33885 10764
rect 33919 10761 33931 10795
rect 33873 10755 33931 10761
rect 35866 10764 36768 10792
rect 14090 10724 14096 10736
rect 1268 10696 2360 10724
rect 2746 10696 14096 10724
rect 1268 10684 1274 10696
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 2332 10665 2360 10696
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 16758 10724 16764 10736
rect 14875 10696 16764 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 16758 10684 16764 10696
rect 16816 10684 16822 10736
rect 17034 10684 17040 10736
rect 17092 10724 17098 10736
rect 17497 10727 17555 10733
rect 17497 10724 17509 10727
rect 17092 10696 17509 10724
rect 17092 10684 17098 10696
rect 17497 10693 17509 10696
rect 17543 10693 17555 10727
rect 19981 10727 20039 10733
rect 19981 10724 19993 10727
rect 17497 10687 17555 10693
rect 18064 10696 19993 10724
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1360 10628 1593 10656
rect 1360 10616 1366 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2363 10628 2881 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 1596 10588 1624 10619
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 12308 10628 13553 10656
rect 12308 10616 12314 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 13541 10619 13599 10625
rect 13740 10628 14749 10656
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 1596 10560 3065 10588
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 13262 10588 13268 10600
rect 12759 10560 13268 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 13262 10548 13268 10560
rect 13320 10588 13326 10600
rect 13633 10591 13691 10597
rect 13633 10588 13645 10591
rect 13320 10560 13645 10588
rect 13320 10548 13326 10560
rect 13633 10557 13645 10560
rect 13679 10557 13691 10591
rect 13633 10551 13691 10557
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 13446 10520 13452 10532
rect 2547 10492 13452 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 12250 10412 12256 10464
rect 12308 10412 12314 10464
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12584 10424 12909 10452
rect 12584 10412 12590 10424
rect 12897 10421 12909 10424
rect 12943 10452 12955 10455
rect 13740 10452 13768 10628
rect 14737 10625 14749 10628
rect 14783 10656 14795 10659
rect 16206 10656 16212 10668
rect 14783 10628 16212 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 17310 10656 17316 10668
rect 16899 10628 17316 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 17310 10616 17316 10628
rect 17368 10656 17374 10668
rect 18064 10656 18092 10696
rect 19981 10693 19993 10696
rect 20027 10693 20039 10727
rect 20990 10724 20996 10736
rect 19981 10687 20039 10693
rect 20180 10696 20996 10724
rect 17368 10628 18092 10656
rect 17368 10616 17374 10628
rect 18414 10616 18420 10668
rect 18472 10656 18478 10668
rect 18472 10628 18552 10656
rect 18472 10616 18478 10628
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 14550 10588 14556 10600
rect 13863 10560 14556 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15068 10560 16037 10588
rect 15068 10548 15074 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 13998 10480 14004 10532
rect 14056 10520 14062 10532
rect 16132 10520 16160 10551
rect 16666 10548 16672 10600
rect 16724 10588 16730 10600
rect 17586 10588 17592 10600
rect 16724 10560 17592 10588
rect 16724 10548 16730 10560
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 17678 10548 17684 10600
rect 17736 10548 17742 10600
rect 18524 10520 18552 10628
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 18966 10656 18972 10668
rect 18831 10628 18972 10656
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 18966 10616 18972 10628
rect 19024 10656 19030 10668
rect 19889 10659 19947 10665
rect 19024 10628 19334 10656
rect 19024 10616 19030 10628
rect 18877 10591 18935 10597
rect 18877 10557 18889 10591
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 18892 10520 18920 10551
rect 14056 10492 16160 10520
rect 16960 10492 18460 10520
rect 18524 10492 18920 10520
rect 19306 10520 19334 10628
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 20180 10656 20208 10696
rect 20990 10684 20996 10696
rect 21048 10684 21054 10736
rect 21177 10727 21235 10733
rect 21177 10693 21189 10727
rect 21223 10724 21235 10727
rect 22278 10724 22284 10736
rect 21223 10696 22284 10724
rect 21223 10693 21235 10696
rect 21177 10687 21235 10693
rect 22278 10684 22284 10696
rect 22336 10684 22342 10736
rect 23566 10684 23572 10736
rect 23624 10724 23630 10736
rect 26142 10724 26148 10736
rect 23624 10696 26148 10724
rect 23624 10684 23630 10696
rect 26142 10684 26148 10696
rect 26200 10684 26206 10736
rect 27430 10684 27436 10736
rect 27488 10724 27494 10736
rect 28537 10727 28595 10733
rect 27488 10696 27660 10724
rect 27488 10684 27494 10696
rect 19935 10628 20208 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 19904 10588 19932 10619
rect 20254 10616 20260 10668
rect 20312 10656 20318 10668
rect 20312 10628 21496 10656
rect 20312 10616 20318 10628
rect 19978 10588 19984 10600
rect 19904 10560 19984 10588
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 21082 10588 21088 10600
rect 20211 10560 21088 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 21082 10548 21088 10560
rect 21140 10548 21146 10600
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 21266 10520 21272 10532
rect 19306 10492 21272 10520
rect 14056 10480 14062 10492
rect 12943 10424 13768 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 15562 10412 15568 10464
rect 15620 10412 15626 10464
rect 15654 10412 15660 10464
rect 15712 10452 15718 10464
rect 16960 10452 16988 10492
rect 15712 10424 16988 10452
rect 15712 10412 15718 10424
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 17092 10424 18337 10452
rect 17092 10412 17098 10424
rect 18325 10421 18337 10424
rect 18371 10421 18383 10455
rect 18432 10452 18460 10492
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 18432 10424 20729 10452
rect 18325 10415 18383 10421
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 21376 10452 21404 10551
rect 21468 10520 21496 10628
rect 23382 10616 23388 10668
rect 23440 10616 23446 10668
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25409 10659 25467 10665
rect 25409 10656 25421 10659
rect 24627 10628 25421 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 25409 10625 25421 10628
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 26326 10616 26332 10668
rect 26384 10616 26390 10668
rect 26789 10659 26847 10665
rect 26789 10625 26801 10659
rect 26835 10656 26847 10659
rect 27448 10656 27476 10684
rect 26835 10628 27476 10656
rect 26835 10625 26847 10628
rect 26789 10619 26847 10625
rect 27522 10616 27528 10668
rect 27580 10616 27586 10668
rect 27632 10656 27660 10696
rect 28537 10693 28549 10727
rect 28583 10724 28595 10727
rect 28810 10724 28816 10736
rect 28583 10696 28816 10724
rect 28583 10693 28595 10696
rect 28537 10687 28595 10693
rect 28810 10684 28816 10696
rect 28868 10684 28874 10736
rect 28966 10696 32812 10724
rect 28966 10656 28994 10696
rect 27632 10628 28994 10656
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 30561 10659 30619 10665
rect 30561 10656 30573 10659
rect 29972 10628 30573 10656
rect 29972 10616 29978 10628
rect 30561 10625 30573 10628
rect 30607 10625 30619 10659
rect 30561 10619 30619 10625
rect 30650 10616 30656 10668
rect 30708 10656 30714 10668
rect 32677 10659 32735 10665
rect 32677 10656 32689 10659
rect 30708 10628 32689 10656
rect 30708 10616 30714 10628
rect 32677 10625 32689 10628
rect 32723 10625 32735 10659
rect 32677 10619 32735 10625
rect 22002 10548 22008 10600
rect 22060 10548 22066 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22112 10560 22293 10588
rect 22112 10520 22140 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 23934 10548 23940 10600
rect 23992 10588 23998 10600
rect 24486 10588 24492 10600
rect 23992 10560 24492 10588
rect 23992 10548 23998 10560
rect 24486 10548 24492 10560
rect 24544 10588 24550 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 24544 10560 24685 10588
rect 24544 10548 24550 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 24857 10591 24915 10597
rect 24857 10557 24869 10591
rect 24903 10588 24915 10591
rect 26602 10588 26608 10600
rect 24903 10560 26608 10588
rect 24903 10557 24915 10560
rect 24857 10551 24915 10557
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 27062 10548 27068 10600
rect 27120 10588 27126 10600
rect 27249 10591 27307 10597
rect 27249 10588 27261 10591
rect 27120 10560 27261 10588
rect 27120 10548 27126 10560
rect 27249 10557 27261 10560
rect 27295 10557 27307 10591
rect 27249 10551 27307 10557
rect 27433 10591 27491 10597
rect 27433 10557 27445 10591
rect 27479 10557 27491 10591
rect 27433 10551 27491 10557
rect 21468 10492 22140 10520
rect 23566 10480 23572 10532
rect 23624 10520 23630 10532
rect 26053 10523 26111 10529
rect 26053 10520 26065 10523
rect 23624 10492 26065 10520
rect 23624 10480 23630 10492
rect 26053 10489 26065 10492
rect 26099 10520 26111 10523
rect 27448 10520 27476 10551
rect 29546 10548 29552 10600
rect 29604 10548 29610 10600
rect 29822 10548 29828 10600
rect 29880 10588 29886 10600
rect 30377 10591 30435 10597
rect 30377 10588 30389 10591
rect 29880 10560 30389 10588
rect 29880 10548 29886 10560
rect 30377 10557 30389 10560
rect 30423 10557 30435 10591
rect 30377 10551 30435 10557
rect 30466 10548 30472 10600
rect 30524 10548 30530 10600
rect 30834 10548 30840 10600
rect 30892 10588 30898 10600
rect 32306 10588 32312 10600
rect 30892 10560 32312 10588
rect 30892 10548 30898 10560
rect 32306 10548 32312 10560
rect 32364 10548 32370 10600
rect 32398 10548 32404 10600
rect 32456 10548 32462 10600
rect 32585 10591 32643 10597
rect 32585 10557 32597 10591
rect 32631 10557 32643 10591
rect 32784 10588 32812 10696
rect 33226 10684 33232 10736
rect 33284 10724 33290 10736
rect 33413 10727 33471 10733
rect 33413 10724 33425 10727
rect 33284 10696 33425 10724
rect 33284 10684 33290 10696
rect 33413 10693 33425 10696
rect 33459 10724 33471 10727
rect 33502 10724 33508 10736
rect 33459 10696 33508 10724
rect 33459 10693 33471 10696
rect 33413 10687 33471 10693
rect 33502 10684 33508 10696
rect 33560 10724 33566 10736
rect 33560 10696 34178 10724
rect 33560 10684 33566 10696
rect 35250 10684 35256 10736
rect 35308 10724 35314 10736
rect 35866 10724 35894 10764
rect 35308 10696 35894 10724
rect 35308 10684 35314 10696
rect 35618 10616 35624 10668
rect 35676 10616 35682 10668
rect 35710 10616 35716 10668
rect 35768 10656 35774 10668
rect 35768 10628 36216 10656
rect 35768 10616 35774 10628
rect 35250 10588 35256 10600
rect 32784 10560 35256 10588
rect 32585 10551 32643 10557
rect 26099 10492 27476 10520
rect 26099 10489 26111 10492
rect 26053 10483 26111 10489
rect 22094 10452 22100 10464
rect 21376 10424 22100 10452
rect 20717 10415 20775 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 23750 10412 23756 10464
rect 23808 10452 23814 10464
rect 24762 10452 24768 10464
rect 23808 10424 24768 10452
rect 23808 10412 23814 10424
rect 24762 10412 24768 10424
rect 24820 10412 24826 10464
rect 27448 10452 27476 10492
rect 27893 10523 27951 10529
rect 27893 10489 27905 10523
rect 27939 10520 27951 10523
rect 32600 10520 32628 10551
rect 35250 10548 35256 10560
rect 35308 10548 35314 10600
rect 36188 10597 36216 10628
rect 36446 10616 36452 10668
rect 36504 10616 36510 10668
rect 36740 10656 36768 10764
rect 36814 10752 36820 10804
rect 36872 10752 36878 10804
rect 38562 10684 38568 10736
rect 38620 10724 38626 10736
rect 39761 10727 39819 10733
rect 39761 10724 39773 10727
rect 38620 10696 39773 10724
rect 38620 10684 38626 10696
rect 39761 10693 39773 10696
rect 39807 10724 39819 10727
rect 40221 10727 40279 10733
rect 40221 10724 40233 10727
rect 39807 10696 40233 10724
rect 39807 10693 39819 10696
rect 39761 10687 39819 10693
rect 40221 10693 40233 10696
rect 40267 10693 40279 10727
rect 40221 10687 40279 10693
rect 49145 10727 49203 10733
rect 49145 10693 49157 10727
rect 49191 10724 49203 10727
rect 49234 10724 49240 10736
rect 49191 10696 49240 10724
rect 49191 10693 49203 10696
rect 49145 10687 49203 10693
rect 49234 10684 49240 10696
rect 49292 10684 49298 10736
rect 38930 10656 38936 10668
rect 36740 10628 38936 10656
rect 38930 10616 38936 10628
rect 38988 10616 38994 10668
rect 46934 10616 46940 10668
rect 46992 10656 46998 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 46992 10628 47961 10656
rect 46992 10616 46998 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 35345 10591 35403 10597
rect 35345 10557 35357 10591
rect 35391 10588 35403 10591
rect 36173 10591 36231 10597
rect 35391 10560 35894 10588
rect 35391 10557 35403 10560
rect 35345 10551 35403 10557
rect 27939 10492 32628 10520
rect 33045 10523 33103 10529
rect 27939 10489 27951 10492
rect 27893 10483 27951 10489
rect 33045 10489 33057 10523
rect 33091 10520 33103 10523
rect 35866 10520 35894 10560
rect 36173 10557 36185 10591
rect 36219 10557 36231 10591
rect 36173 10551 36231 10557
rect 36354 10548 36360 10600
rect 36412 10548 36418 10600
rect 36538 10548 36544 10600
rect 36596 10588 36602 10600
rect 36906 10588 36912 10600
rect 36596 10560 36912 10588
rect 36596 10548 36602 10560
rect 36906 10548 36912 10560
rect 36964 10588 36970 10600
rect 37277 10591 37335 10597
rect 37277 10588 37289 10591
rect 36964 10560 37289 10588
rect 36964 10548 36970 10560
rect 37277 10557 37289 10560
rect 37323 10588 37335 10591
rect 37461 10591 37519 10597
rect 37461 10588 37473 10591
rect 37323 10560 37473 10588
rect 37323 10557 37335 10560
rect 37277 10551 37335 10557
rect 37461 10557 37473 10560
rect 37507 10557 37519 10591
rect 37461 10551 37519 10557
rect 36630 10520 36636 10532
rect 33091 10492 34376 10520
rect 35866 10492 36636 10520
rect 33091 10489 33103 10492
rect 33045 10483 33103 10489
rect 30834 10452 30840 10464
rect 27448 10424 30840 10452
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 30929 10455 30987 10461
rect 30929 10421 30941 10455
rect 30975 10452 30987 10455
rect 31754 10452 31760 10464
rect 30975 10424 31760 10452
rect 30975 10421 30987 10424
rect 30929 10415 30987 10421
rect 31754 10412 31760 10424
rect 31812 10412 31818 10464
rect 31938 10412 31944 10464
rect 31996 10452 32002 10464
rect 32858 10452 32864 10464
rect 31996 10424 32864 10452
rect 31996 10412 32002 10424
rect 32858 10412 32864 10424
rect 32916 10412 32922 10464
rect 34348 10452 34376 10492
rect 36630 10480 36636 10492
rect 36688 10480 36694 10532
rect 37550 10520 37556 10532
rect 36740 10492 37556 10520
rect 36740 10452 36768 10492
rect 37550 10480 37556 10492
rect 37608 10480 37614 10532
rect 39945 10523 40003 10529
rect 39945 10489 39957 10523
rect 39991 10520 40003 10523
rect 47118 10520 47124 10532
rect 39991 10492 47124 10520
rect 39991 10489 40003 10492
rect 39945 10483 40003 10489
rect 47118 10480 47124 10492
rect 47176 10480 47182 10532
rect 34348 10424 36768 10452
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 13449 10251 13507 10257
rect 13449 10217 13461 10251
rect 13495 10248 13507 10251
rect 15010 10248 15016 10260
rect 13495 10220 15016 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 16114 10248 16120 10260
rect 16040 10220 16120 10248
rect 4798 10140 4804 10192
rect 4856 10180 4862 10192
rect 12526 10180 12532 10192
rect 4856 10152 12532 10180
rect 4856 10140 4862 10152
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 13909 10183 13967 10189
rect 13909 10149 13921 10183
rect 13955 10180 13967 10183
rect 14734 10180 14740 10192
rect 13955 10152 14740 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 2130 10072 2136 10124
rect 2188 10072 2194 10124
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 16040 10112 16068 10220
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 16482 10208 16488 10260
rect 16540 10208 16546 10260
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 18322 10248 18328 10260
rect 18187 10220 18328 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 20220 10220 20269 10248
rect 20220 10208 20226 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 20364 10220 22094 10248
rect 17678 10180 17684 10192
rect 13035 10084 16068 10112
rect 16132 10152 17684 10180
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 2406 10004 2412 10056
rect 2464 10004 2470 10056
rect 12912 9976 12940 10075
rect 13078 10004 13084 10056
rect 13136 10044 13142 10056
rect 14274 10044 14280 10056
rect 13136 10016 14280 10044
rect 13136 10004 13142 10016
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 14182 9976 14188 9988
rect 12912 9948 14188 9976
rect 14182 9936 14188 9948
rect 14240 9976 14246 9988
rect 15749 9979 15807 9985
rect 14240 9948 14412 9976
rect 14240 9936 14246 9948
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13078 9908 13084 9920
rect 12492 9880 13084 9908
rect 12492 9868 12498 9880
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14277 9911 14335 9917
rect 14277 9908 14289 9911
rect 13964 9880 14289 9908
rect 13964 9868 13970 9880
rect 14277 9877 14289 9880
rect 14323 9877 14335 9911
rect 14384 9908 14412 9948
rect 15749 9945 15761 9979
rect 15795 9976 15807 9979
rect 16132 9976 16160 10152
rect 17678 10140 17684 10152
rect 17736 10140 17742 10192
rect 16298 10072 16304 10124
rect 16356 10112 16362 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 16356 10084 17417 10112
rect 16356 10072 16362 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10112 17647 10115
rect 17862 10112 17868 10124
rect 17635 10084 17868 10112
rect 17635 10081 17647 10084
rect 17589 10075 17647 10081
rect 17862 10072 17868 10084
rect 17920 10112 17926 10124
rect 18414 10112 18420 10124
rect 17920 10084 18420 10112
rect 17920 10072 17926 10084
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 18598 10072 18604 10124
rect 18656 10072 18662 10124
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 19426 10112 19432 10124
rect 18831 10084 19432 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19668 10084 19717 10112
rect 19668 10072 19674 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 16206 10004 16212 10056
rect 16264 10044 16270 10056
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 16264 10016 18521 10044
rect 16264 10004 16270 10016
rect 18509 10013 18521 10016
rect 18555 10044 18567 10047
rect 20364 10044 20392 10220
rect 22066 10180 22094 10220
rect 23658 10208 23664 10260
rect 23716 10248 23722 10260
rect 24486 10248 24492 10260
rect 23716 10220 24492 10248
rect 23716 10208 23722 10220
rect 24486 10208 24492 10220
rect 24544 10248 24550 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 24544 10220 24593 10248
rect 24544 10208 24550 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 26326 10248 26332 10260
rect 24581 10211 24639 10217
rect 24688 10220 26332 10248
rect 24688 10180 24716 10220
rect 26326 10208 26332 10220
rect 26384 10248 26390 10260
rect 27430 10248 27436 10260
rect 26384 10220 27436 10248
rect 26384 10208 26390 10220
rect 27430 10208 27436 10220
rect 27488 10208 27494 10260
rect 28721 10251 28779 10257
rect 28721 10217 28733 10251
rect 28767 10248 28779 10251
rect 29086 10248 29092 10260
rect 28767 10220 29092 10248
rect 28767 10217 28779 10220
rect 28721 10211 28779 10217
rect 29086 10208 29092 10220
rect 29144 10248 29150 10260
rect 29822 10248 29828 10260
rect 29144 10220 29828 10248
rect 29144 10208 29150 10220
rect 29822 10208 29828 10220
rect 29880 10208 29886 10260
rect 30377 10251 30435 10257
rect 30377 10217 30389 10251
rect 30423 10248 30435 10251
rect 31386 10248 31392 10260
rect 30423 10220 31392 10248
rect 30423 10217 30435 10220
rect 30377 10211 30435 10217
rect 31386 10208 31392 10220
rect 31444 10208 31450 10260
rect 32582 10248 32588 10260
rect 32048 10220 32588 10248
rect 26602 10180 26608 10192
rect 22066 10152 24716 10180
rect 26252 10152 26608 10180
rect 20438 10072 20444 10124
rect 20496 10112 20502 10124
rect 20714 10112 20720 10124
rect 20496 10084 20720 10112
rect 20496 10072 20502 10084
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21729 10115 21787 10121
rect 21729 10112 21741 10115
rect 21140 10084 21741 10112
rect 21140 10072 21146 10084
rect 21729 10081 21741 10084
rect 21775 10081 21787 10115
rect 21729 10075 21787 10081
rect 23753 10115 23811 10121
rect 23753 10081 23765 10115
rect 23799 10112 23811 10115
rect 23842 10112 23848 10124
rect 23799 10084 23848 10112
rect 23799 10081 23811 10084
rect 23753 10075 23811 10081
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10112 26111 10115
rect 26252 10112 26280 10152
rect 26602 10140 26608 10152
rect 26660 10140 26666 10192
rect 26694 10140 26700 10192
rect 26752 10140 26758 10192
rect 29270 10140 29276 10192
rect 29328 10140 29334 10192
rect 26099 10084 26280 10112
rect 26329 10115 26387 10121
rect 26099 10081 26111 10084
rect 26053 10075 26111 10081
rect 26329 10081 26341 10115
rect 26375 10112 26387 10115
rect 26878 10112 26884 10124
rect 26375 10084 26884 10112
rect 26375 10081 26387 10084
rect 26329 10075 26387 10081
rect 26878 10072 26884 10084
rect 26936 10112 26942 10124
rect 26973 10115 27031 10121
rect 26973 10112 26985 10115
rect 26936 10084 26985 10112
rect 26936 10072 26942 10084
rect 26973 10081 26985 10084
rect 27019 10112 27031 10115
rect 29546 10112 29552 10124
rect 27019 10084 29552 10112
rect 27019 10081 27031 10084
rect 26973 10075 27031 10081
rect 29546 10072 29552 10084
rect 29604 10072 29610 10124
rect 29917 10115 29975 10121
rect 29917 10081 29929 10115
rect 29963 10112 29975 10115
rect 30650 10112 30656 10124
rect 29963 10084 30656 10112
rect 29963 10081 29975 10084
rect 29917 10075 29975 10081
rect 30650 10072 30656 10084
rect 30708 10072 30714 10124
rect 30834 10072 30840 10124
rect 30892 10112 30898 10124
rect 32048 10112 32076 10220
rect 32582 10208 32588 10220
rect 32640 10248 32646 10260
rect 35710 10248 35716 10260
rect 32640 10220 35716 10248
rect 32640 10208 32646 10220
rect 35710 10208 35716 10220
rect 35768 10208 35774 10260
rect 36630 10208 36636 10260
rect 36688 10208 36694 10260
rect 36906 10208 36912 10260
rect 36964 10208 36970 10260
rect 32214 10140 32220 10192
rect 32272 10180 32278 10192
rect 32272 10152 32904 10180
rect 32272 10140 32278 10152
rect 30892 10084 32076 10112
rect 30892 10072 30898 10084
rect 32122 10072 32128 10124
rect 32180 10072 32186 10124
rect 32582 10072 32588 10124
rect 32640 10112 32646 10124
rect 32876 10121 32904 10152
rect 32677 10115 32735 10121
rect 32677 10112 32689 10115
rect 32640 10084 32689 10112
rect 32640 10072 32646 10084
rect 32677 10081 32689 10084
rect 32723 10081 32735 10115
rect 32677 10075 32735 10081
rect 32861 10115 32919 10121
rect 32861 10081 32873 10115
rect 32907 10081 32919 10115
rect 32861 10075 32919 10081
rect 34698 10072 34704 10124
rect 34756 10112 34762 10124
rect 35161 10115 35219 10121
rect 35161 10112 35173 10115
rect 34756 10084 35173 10112
rect 34756 10072 34762 10084
rect 35161 10081 35173 10084
rect 35207 10112 35219 10115
rect 35618 10112 35624 10124
rect 35207 10084 35624 10112
rect 35207 10081 35219 10084
rect 35161 10075 35219 10081
rect 35618 10072 35624 10084
rect 35676 10072 35682 10124
rect 35710 10072 35716 10124
rect 35768 10112 35774 10124
rect 40589 10115 40647 10121
rect 40589 10112 40601 10115
rect 35768 10084 38332 10112
rect 35768 10072 35774 10084
rect 18555 10016 20392 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 15795 9948 16160 9976
rect 15795 9945 15807 9948
rect 15749 9939 15807 9945
rect 15764 9908 15792 9939
rect 16758 9936 16764 9988
rect 16816 9976 16822 9988
rect 16816 9948 20392 9976
rect 20732 9962 20760 10072
rect 22002 10004 22008 10056
rect 22060 10044 22066 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 22060 10016 23213 10044
rect 22060 10004 22066 10016
rect 23201 10013 23213 10016
rect 23247 10044 23259 10047
rect 24026 10044 24032 10056
rect 23247 10016 24032 10044
rect 23247 10013 23259 10016
rect 23201 10007 23259 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 32766 10004 32772 10056
rect 32824 10044 32830 10056
rect 33781 10047 33839 10053
rect 33781 10044 33793 10047
rect 32824 10016 33793 10044
rect 32824 10004 32830 10016
rect 33781 10013 33793 10016
rect 33827 10013 33839 10047
rect 33781 10007 33839 10013
rect 34882 10004 34888 10056
rect 34940 10004 34946 10056
rect 36538 10044 36544 10056
rect 36294 10016 36544 10044
rect 36538 10004 36544 10016
rect 36596 10004 36602 10056
rect 38304 10053 38332 10084
rect 40144 10084 40601 10112
rect 38289 10047 38347 10053
rect 38289 10013 38301 10047
rect 38335 10044 38347 10047
rect 38749 10047 38807 10053
rect 38749 10044 38761 10047
rect 38335 10016 38761 10044
rect 38335 10013 38347 10016
rect 38289 10007 38347 10013
rect 38749 10013 38761 10016
rect 38795 10013 38807 10047
rect 38749 10007 38807 10013
rect 38930 10004 38936 10056
rect 38988 10044 38994 10056
rect 40144 10053 40172 10084
rect 40589 10081 40601 10084
rect 40635 10081 40647 10115
rect 40589 10075 40647 10081
rect 49142 10072 49148 10124
rect 49200 10072 49206 10124
rect 40129 10047 40187 10053
rect 40129 10044 40141 10047
rect 38988 10016 40141 10044
rect 38988 10004 38994 10016
rect 40129 10013 40141 10016
rect 40175 10013 40187 10047
rect 40129 10007 40187 10013
rect 40313 10047 40371 10053
rect 40313 10013 40325 10047
rect 40359 10044 40371 10047
rect 45830 10044 45836 10056
rect 40359 10016 45836 10044
rect 40359 10013 40371 10016
rect 40313 10007 40371 10013
rect 45830 10004 45836 10016
rect 45888 10004 45894 10056
rect 46106 10004 46112 10056
rect 46164 10004 46170 10056
rect 46566 10004 46572 10056
rect 46624 10044 46630 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46624 10016 47961 10044
rect 46624 10004 46630 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 22465 9979 22523 9985
rect 16816 9936 16822 9948
rect 14384 9880 15792 9908
rect 14277 9871 14335 9877
rect 16574 9868 16580 9920
rect 16632 9868 16638 9920
rect 16942 9868 16948 9920
rect 17000 9868 17006 9920
rect 17310 9868 17316 9920
rect 17368 9868 17374 9920
rect 20364 9908 20392 9948
rect 22465 9945 22477 9979
rect 22511 9976 22523 9979
rect 22554 9976 22560 9988
rect 22511 9948 22560 9976
rect 22511 9945 22523 9948
rect 22465 9939 22523 9945
rect 22554 9936 22560 9948
rect 22612 9936 22618 9988
rect 23382 9936 23388 9988
rect 23440 9976 23446 9988
rect 23845 9979 23903 9985
rect 23845 9976 23857 9979
rect 23440 9948 23857 9976
rect 23440 9936 23446 9948
rect 23845 9945 23857 9948
rect 23891 9976 23903 9979
rect 24394 9976 24400 9988
rect 23891 9948 24400 9976
rect 23891 9945 23903 9948
rect 23845 9939 23903 9945
rect 24394 9936 24400 9948
rect 24452 9936 24458 9988
rect 25590 9936 25596 9988
rect 25648 9976 25654 9988
rect 25774 9976 25780 9988
rect 25648 9948 25780 9976
rect 25648 9936 25654 9948
rect 25774 9936 25780 9948
rect 25832 9936 25838 9988
rect 27249 9979 27307 9985
rect 27249 9945 27261 9979
rect 27295 9976 27307 9979
rect 27338 9976 27344 9988
rect 27295 9948 27344 9976
rect 27295 9945 27307 9948
rect 27249 9939 27307 9945
rect 27338 9936 27344 9948
rect 27396 9936 27402 9988
rect 27448 9948 27738 9976
rect 23566 9908 23572 9920
rect 20364 9880 23572 9908
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 23934 9868 23940 9920
rect 23992 9908 23998 9920
rect 24029 9911 24087 9917
rect 24029 9908 24041 9911
rect 23992 9880 24041 9908
rect 23992 9868 23998 9880
rect 24029 9877 24041 9880
rect 24075 9877 24087 9911
rect 24029 9871 24087 9877
rect 26694 9868 26700 9920
rect 26752 9908 26758 9920
rect 27448 9908 27476 9948
rect 30834 9936 30840 9988
rect 30892 9936 30898 9988
rect 31846 9936 31852 9988
rect 31904 9936 31910 9988
rect 31938 9936 31944 9988
rect 31996 9976 32002 9988
rect 32953 9979 33011 9985
rect 32953 9976 32965 9979
rect 31996 9948 32965 9976
rect 31996 9936 32002 9948
rect 32953 9945 32965 9948
rect 32999 9945 33011 9979
rect 37458 9976 37464 9988
rect 32953 9939 33011 9945
rect 33336 9948 34652 9976
rect 28902 9908 28908 9920
rect 26752 9880 28908 9908
rect 26752 9868 26758 9880
rect 28902 9868 28908 9880
rect 28960 9908 28966 9920
rect 28997 9911 29055 9917
rect 28997 9908 29009 9911
rect 28960 9880 29009 9908
rect 28960 9868 28966 9880
rect 28997 9877 29009 9880
rect 29043 9877 29055 9911
rect 28997 9871 29055 9877
rect 30098 9868 30104 9920
rect 30156 9908 30162 9920
rect 33226 9908 33232 9920
rect 30156 9880 33232 9908
rect 30156 9868 30162 9880
rect 33226 9868 33232 9880
rect 33284 9868 33290 9920
rect 33336 9917 33364 9948
rect 33321 9911 33379 9917
rect 33321 9877 33333 9911
rect 33367 9877 33379 9911
rect 34624 9908 34652 9948
rect 36556 9948 37464 9976
rect 36556 9908 36584 9948
rect 37458 9936 37464 9948
rect 37516 9936 37522 9988
rect 44358 9936 44364 9988
rect 44416 9936 44422 9988
rect 44545 9979 44603 9985
rect 44545 9945 44557 9979
rect 44591 9976 44603 9979
rect 46750 9976 46756 9988
rect 44591 9948 46756 9976
rect 44591 9945 44603 9948
rect 44545 9939 44603 9945
rect 46750 9936 46756 9948
rect 46808 9936 46814 9988
rect 47302 9936 47308 9988
rect 47360 9936 47366 9988
rect 34624 9880 36584 9908
rect 33321 9871 33379 9877
rect 38378 9868 38384 9920
rect 38436 9868 38442 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 2133 9707 2191 9713
rect 2133 9704 2145 9707
rect 1360 9676 2145 9704
rect 1360 9664 1366 9676
rect 2133 9673 2145 9676
rect 2179 9704 2191 9707
rect 2406 9704 2412 9716
rect 2179 9676 2412 9704
rect 2179 9673 2191 9676
rect 2133 9667 2191 9673
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 16574 9704 16580 9716
rect 14792 9676 16580 9704
rect 14792 9664 14798 9676
rect 16574 9664 16580 9676
rect 16632 9704 16638 9716
rect 19978 9704 19984 9716
rect 16632 9676 19984 9704
rect 16632 9664 16638 9676
rect 19978 9664 19984 9676
rect 20036 9664 20042 9716
rect 21082 9664 21088 9716
rect 21140 9664 21146 9716
rect 22278 9664 22284 9716
rect 22336 9664 22342 9716
rect 22554 9664 22560 9716
rect 22612 9704 22618 9716
rect 24578 9704 24584 9716
rect 22612 9676 24584 9704
rect 22612 9664 22618 9676
rect 24578 9664 24584 9676
rect 24636 9704 24642 9716
rect 28810 9704 28816 9716
rect 24636 9676 28816 9704
rect 24636 9664 24642 9676
rect 28810 9664 28816 9676
rect 28868 9664 28874 9716
rect 28902 9664 28908 9716
rect 28960 9704 28966 9716
rect 30650 9704 30656 9716
rect 28960 9676 30656 9704
rect 28960 9664 28966 9676
rect 30650 9664 30656 9676
rect 30708 9704 30714 9716
rect 30834 9704 30840 9716
rect 30708 9676 30840 9704
rect 30708 9664 30714 9676
rect 30834 9664 30840 9676
rect 30892 9664 30898 9716
rect 31478 9664 31484 9716
rect 31536 9704 31542 9716
rect 31757 9707 31815 9713
rect 31757 9704 31769 9707
rect 31536 9676 31769 9704
rect 31536 9664 31542 9676
rect 31757 9673 31769 9676
rect 31803 9673 31815 9707
rect 32861 9707 32919 9713
rect 32861 9704 32873 9707
rect 31757 9667 31815 9673
rect 32048 9676 32873 9704
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12618 9636 12624 9648
rect 12483 9608 12624 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 13357 9639 13415 9645
rect 13357 9605 13369 9639
rect 13403 9636 13415 9639
rect 13722 9636 13728 9648
rect 13403 9608 13728 9636
rect 13403 9605 13415 9608
rect 13357 9599 13415 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 15102 9636 15108 9648
rect 14674 9608 15108 9636
rect 15102 9596 15108 9608
rect 15160 9596 15166 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 16022 9636 16028 9648
rect 15252 9608 16028 9636
rect 15252 9596 15258 9608
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1360 9540 1593 9568
rect 1360 9528 1366 9540
rect 1581 9537 1593 9540
rect 1627 9568 1639 9571
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1627 9540 2329 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 15396 9577 15424 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 16117 9639 16175 9645
rect 16117 9605 16129 9639
rect 16163 9636 16175 9639
rect 16206 9636 16212 9648
rect 16163 9608 16212 9636
rect 16163 9605 16175 9608
rect 16117 9599 16175 9605
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 16301 9639 16359 9645
rect 16301 9605 16313 9639
rect 16347 9636 16359 9639
rect 16666 9636 16672 9648
rect 16347 9608 16672 9636
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 16850 9596 16856 9648
rect 16908 9596 16914 9648
rect 18322 9636 18328 9648
rect 18170 9608 18328 9636
rect 18322 9596 18328 9608
rect 18380 9596 18386 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 19613 9639 19671 9645
rect 19613 9636 19625 9639
rect 19576 9608 19625 9636
rect 19576 9596 19582 9608
rect 19613 9605 19625 9608
rect 19659 9605 19671 9639
rect 19613 9599 19671 9605
rect 20346 9596 20352 9648
rect 20404 9596 20410 9648
rect 21266 9596 21272 9648
rect 21324 9636 21330 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 21324 9608 21373 9636
rect 21324 9596 21330 9608
rect 21361 9605 21373 9608
rect 21407 9605 21419 9639
rect 21361 9599 21419 9605
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12400 9540 12541 9568
rect 12400 9528 12406 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 15838 9528 15844 9580
rect 15896 9528 15902 9580
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11112 9472 12265 9500
rect 11112 9460 11118 9472
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 15102 9460 15108 9512
rect 15160 9460 15166 9512
rect 18598 9460 18604 9512
rect 18656 9460 18662 9512
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 19337 9503 19395 9509
rect 19337 9500 19349 9503
rect 18932 9472 19349 9500
rect 18932 9460 18938 9472
rect 19337 9469 19349 9472
rect 19383 9469 19395 9503
rect 21376 9500 21404 9599
rect 24394 9596 24400 9648
rect 24452 9596 24458 9648
rect 24670 9596 24676 9648
rect 24728 9636 24734 9648
rect 27338 9636 27344 9648
rect 24728 9608 25268 9636
rect 24728 9596 24734 9608
rect 22646 9528 22652 9580
rect 22704 9528 22710 9580
rect 25240 9577 25268 9608
rect 25976 9608 27344 9636
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 25225 9571 25283 9577
rect 22787 9540 23612 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 22756 9500 22784 9531
rect 21376 9472 22784 9500
rect 22925 9503 22983 9509
rect 19337 9463 19395 9469
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23584 9500 23612 9540
rect 25225 9537 25237 9571
rect 25271 9537 25283 9571
rect 25976 9568 26004 9608
rect 27338 9596 27344 9608
rect 27396 9596 27402 9648
rect 28920 9636 28948 9664
rect 28566 9608 28948 9636
rect 28997 9639 29055 9645
rect 28997 9605 29009 9639
rect 29043 9636 29055 9639
rect 30098 9636 30104 9648
rect 29043 9608 30104 9636
rect 29043 9605 29055 9608
rect 28997 9599 29055 9605
rect 30098 9596 30104 9608
rect 30156 9596 30162 9648
rect 31662 9596 31668 9648
rect 31720 9636 31726 9648
rect 32048 9636 32076 9676
rect 32861 9673 32873 9676
rect 32907 9673 32919 9707
rect 32861 9667 32919 9673
rect 33502 9664 33508 9716
rect 33560 9704 33566 9716
rect 34422 9704 34428 9716
rect 33560 9676 34428 9704
rect 33560 9664 33566 9676
rect 34422 9664 34428 9676
rect 34480 9664 34486 9716
rect 35618 9664 35624 9716
rect 35676 9664 35682 9716
rect 36173 9707 36231 9713
rect 36173 9673 36185 9707
rect 36219 9704 36231 9707
rect 36538 9704 36544 9716
rect 36219 9676 36544 9704
rect 36219 9673 36231 9676
rect 36173 9667 36231 9673
rect 36538 9664 36544 9676
rect 36596 9664 36602 9716
rect 38378 9664 38384 9716
rect 38436 9704 38442 9716
rect 46934 9704 46940 9716
rect 38436 9676 46940 9704
rect 38436 9664 38442 9676
rect 46934 9664 46940 9676
rect 46992 9664 46998 9716
rect 31720 9608 32076 9636
rect 31720 9596 31726 9608
rect 32122 9596 32128 9648
rect 32180 9636 32186 9648
rect 32180 9608 33916 9636
rect 32180 9596 32186 9608
rect 25225 9531 25283 9537
rect 25884 9540 26004 9568
rect 26053 9571 26111 9577
rect 22971 9472 23520 9500
rect 23584 9472 23888 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 17310 9432 17316 9444
rect 15672 9404 17316 9432
rect 15672 9376 15700 9404
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 14918 9364 14924 9376
rect 12943 9336 14924 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 15654 9324 15660 9376
rect 15712 9324 15718 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16356 9336 16405 9364
rect 16356 9324 16362 9336
rect 16393 9333 16405 9336
rect 16439 9364 16451 9367
rect 18414 9364 18420 9376
rect 16439 9336 18420 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 21542 9324 21548 9376
rect 21600 9324 21606 9376
rect 21818 9324 21824 9376
rect 21876 9324 21882 9376
rect 23492 9373 23520 9472
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23750 9364 23756 9376
rect 23523 9336 23756 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 23860 9364 23888 9472
rect 24486 9460 24492 9512
rect 24544 9500 24550 9512
rect 25884 9509 25912 9540
rect 26053 9537 26065 9571
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 24949 9503 25007 9509
rect 24949 9500 24961 9503
rect 24544 9472 24961 9500
rect 24544 9460 24550 9472
rect 24949 9469 24961 9472
rect 24995 9469 25007 9503
rect 24949 9463 25007 9469
rect 25869 9503 25927 9509
rect 25869 9469 25881 9503
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 25958 9460 25964 9512
rect 26016 9460 26022 9512
rect 25682 9392 25688 9444
rect 25740 9432 25746 9444
rect 26068 9432 26096 9531
rect 31110 9528 31116 9580
rect 31168 9528 31174 9580
rect 31754 9528 31760 9580
rect 31812 9568 31818 9580
rect 33888 9577 33916 9608
rect 34698 9596 34704 9648
rect 34756 9596 34762 9648
rect 49145 9639 49203 9645
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 49234 9636 49240 9648
rect 49191 9608 49240 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 49234 9596 49240 9608
rect 49292 9596 49298 9648
rect 32953 9571 33011 9577
rect 32953 9568 32965 9571
rect 31812 9540 32965 9568
rect 31812 9528 31818 9540
rect 32953 9537 32965 9540
rect 32999 9537 33011 9571
rect 32953 9531 33011 9537
rect 33873 9571 33931 9577
rect 33873 9537 33885 9571
rect 33919 9537 33931 9571
rect 33873 9531 33931 9537
rect 47210 9528 47216 9580
rect 47268 9568 47274 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 47268 9540 47961 9568
rect 47268 9528 47274 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 27154 9460 27160 9512
rect 27212 9500 27218 9512
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27212 9472 27537 9500
rect 27212 9460 27218 9472
rect 27525 9469 27537 9472
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 28000 9472 29224 9500
rect 25740 9404 26096 9432
rect 26421 9435 26479 9441
rect 25740 9392 25746 9404
rect 26421 9401 26433 9435
rect 26467 9432 26479 9435
rect 28000 9432 28028 9472
rect 26467 9404 28028 9432
rect 29196 9432 29224 9472
rect 29270 9460 29276 9512
rect 29328 9500 29334 9512
rect 29546 9500 29552 9512
rect 29328 9472 29552 9500
rect 29328 9460 29334 9472
rect 29546 9460 29552 9472
rect 29604 9500 29610 9512
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29604 9472 29745 9500
rect 29604 9460 29610 9472
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 30006 9500 30012 9512
rect 29733 9463 29791 9469
rect 29840 9472 30012 9500
rect 29196 9404 29408 9432
rect 26467 9401 26479 9404
rect 26421 9395 26479 9401
rect 25866 9364 25872 9376
rect 23860 9336 25872 9364
rect 25866 9324 25872 9336
rect 25924 9324 25930 9376
rect 29380 9364 29408 9404
rect 29454 9392 29460 9444
rect 29512 9432 29518 9444
rect 29840 9432 29868 9472
rect 30006 9460 30012 9472
rect 30064 9460 30070 9512
rect 30098 9460 30104 9512
rect 30156 9500 30162 9512
rect 31481 9503 31539 9509
rect 31481 9500 31493 9503
rect 30156 9472 31493 9500
rect 30156 9460 30162 9472
rect 31481 9469 31493 9472
rect 31527 9500 31539 9503
rect 31527 9472 31754 9500
rect 31527 9469 31539 9472
rect 31481 9463 31539 9469
rect 29512 9404 29868 9432
rect 31726 9432 31754 9472
rect 31846 9460 31852 9512
rect 31904 9500 31910 9512
rect 32677 9503 32735 9509
rect 32677 9500 32689 9503
rect 31904 9472 32689 9500
rect 31904 9460 31910 9472
rect 32677 9469 32689 9472
rect 32723 9469 32735 9503
rect 32677 9463 32735 9469
rect 34149 9503 34207 9509
rect 34149 9469 34161 9503
rect 34195 9500 34207 9503
rect 34238 9500 34244 9512
rect 34195 9472 34244 9500
rect 34195 9469 34207 9472
rect 34149 9463 34207 9469
rect 34238 9460 34244 9472
rect 34296 9500 34302 9512
rect 35897 9503 35955 9509
rect 35897 9500 35909 9503
rect 34296 9472 35909 9500
rect 34296 9460 34302 9472
rect 35897 9469 35909 9472
rect 35943 9500 35955 9503
rect 36078 9500 36084 9512
rect 35943 9472 36084 9500
rect 35943 9469 35955 9472
rect 35897 9463 35955 9469
rect 36078 9460 36084 9472
rect 36136 9460 36142 9512
rect 32582 9432 32588 9444
rect 31726 9404 32588 9432
rect 29512 9392 29518 9404
rect 32582 9392 32588 9404
rect 32640 9392 32646 9444
rect 30466 9364 30472 9376
rect 29380 9336 30472 9364
rect 30466 9324 30472 9336
rect 30524 9324 30530 9376
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 32125 9367 32183 9373
rect 32125 9364 32137 9367
rect 31168 9336 32137 9364
rect 31168 9324 31174 9336
rect 32125 9333 32137 9336
rect 32171 9333 32183 9367
rect 32125 9327 32183 9333
rect 33321 9367 33379 9373
rect 33321 9333 33333 9367
rect 33367 9364 33379 9367
rect 35158 9364 35164 9376
rect 33367 9336 35164 9364
rect 33367 9333 33379 9336
rect 33321 9327 33379 9333
rect 35158 9324 35164 9336
rect 35216 9324 35222 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 1765 9163 1823 9169
rect 1765 9129 1777 9163
rect 1811 9160 1823 9163
rect 1811 9132 15700 9160
rect 1811 9129 1823 9132
rect 1765 9123 1823 9129
rect 2130 9052 2136 9104
rect 2188 9092 2194 9104
rect 15378 9092 15384 9104
rect 2188 9064 15384 9092
rect 2188 9052 2194 9064
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 15672 9092 15700 9132
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 16393 9163 16451 9169
rect 16393 9160 16405 9163
rect 15804 9132 16405 9160
rect 15804 9120 15810 9132
rect 16393 9129 16405 9132
rect 16439 9160 16451 9163
rect 17126 9160 17132 9172
rect 16439 9132 17132 9160
rect 16439 9129 16451 9132
rect 16393 9123 16451 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17862 9120 17868 9172
rect 17920 9169 17926 9172
rect 17920 9163 17935 9169
rect 17923 9129 17935 9163
rect 17920 9123 17935 9129
rect 19429 9163 19487 9169
rect 19429 9129 19441 9163
rect 19475 9160 19487 9163
rect 19518 9160 19524 9172
rect 19475 9132 19524 9160
rect 19475 9129 19487 9132
rect 19429 9123 19487 9129
rect 17920 9120 17926 9123
rect 19518 9120 19524 9132
rect 19576 9120 19582 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22152 9132 22293 9160
rect 22152 9120 22158 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 24489 9163 24547 9169
rect 22281 9123 22339 9129
rect 22480 9132 23980 9160
rect 16758 9092 16764 9104
rect 15672 9064 16764 9092
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2332 8996 2881 9024
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 2332 8965 2360 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 13354 9024 13360 9036
rect 3200 8996 13360 9024
rect 3200 8984 3206 8996
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15160 8996 15301 9024
rect 15160 8984 15166 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15470 8984 15476 9036
rect 15528 8984 15534 9036
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 18141 9027 18199 9033
rect 18141 9024 18153 9027
rect 16540 8996 18153 9024
rect 16540 8984 16546 8996
rect 18141 8993 18153 8996
rect 18187 9024 18199 9027
rect 18874 9024 18880 9036
rect 18187 8996 18880 9024
rect 18187 8993 18199 8996
rect 18141 8987 18199 8993
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 19484 8996 20913 9024
rect 19484 8984 19490 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 1268 8928 2329 8956
rect 1268 8916 1274 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2317 8919 2375 8925
rect 2424 8928 3065 8956
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 1673 8891 1731 8897
rect 1673 8888 1685 8891
rect 1360 8860 1685 8888
rect 1360 8848 1366 8860
rect 1673 8857 1685 8860
rect 1719 8888 1731 8891
rect 2424 8888 2452 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13596 8928 14289 8956
rect 13596 8916 13602 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 15562 8916 15568 8968
rect 15620 8916 15626 8968
rect 18690 8916 18696 8968
rect 18748 8916 18754 8968
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8956 21235 8959
rect 21450 8956 21456 8968
rect 21223 8928 21456 8956
rect 21223 8925 21235 8928
rect 21177 8919 21235 8925
rect 21450 8916 21456 8928
rect 21508 8956 21514 8968
rect 22002 8956 22008 8968
rect 21508 8928 22008 8956
rect 21508 8916 21514 8928
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 1719 8860 2452 8888
rect 2516 8860 3280 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 2516 8829 2544 8860
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 3142 8820 3148 8832
rect 2648 8792 3148 8820
rect 2648 8780 2654 8792
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3252 8820 3280 8860
rect 13722 8848 13728 8900
rect 13780 8888 13786 8900
rect 13780 8860 16068 8888
rect 13780 8848 13786 8860
rect 13814 8820 13820 8832
rect 3252 8792 13820 8820
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14458 8780 14464 8832
rect 14516 8780 14522 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15286 8820 15292 8832
rect 14967 8792 15292 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15930 8780 15936 8832
rect 15988 8780 15994 8832
rect 16040 8820 16068 8860
rect 17402 8848 17408 8900
rect 17460 8888 17466 8900
rect 18414 8888 18420 8900
rect 17460 8860 18420 8888
rect 17460 8848 17466 8860
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 20438 8848 20444 8900
rect 20496 8848 20502 8900
rect 22480 8888 22508 9132
rect 23952 9092 23980 9132
rect 24489 9129 24501 9163
rect 24535 9160 24547 9163
rect 24578 9160 24584 9172
rect 24535 9132 24584 9160
rect 24535 9129 24547 9132
rect 24489 9123 24547 9129
rect 24578 9120 24584 9132
rect 24636 9120 24642 9172
rect 25593 9163 25651 9169
rect 25593 9129 25605 9163
rect 25639 9160 25651 9163
rect 25958 9160 25964 9172
rect 25639 9132 25964 9160
rect 25639 9129 25651 9132
rect 25593 9123 25651 9129
rect 25608 9092 25636 9123
rect 25958 9120 25964 9132
rect 26016 9160 26022 9172
rect 32861 9163 32919 9169
rect 26016 9132 32444 9160
rect 26016 9120 26022 9132
rect 30006 9092 30012 9104
rect 23952 9064 25636 9092
rect 28368 9064 30012 9092
rect 23750 8984 23756 9036
rect 23808 8984 23814 9036
rect 24026 8984 24032 9036
rect 24084 8984 24090 9036
rect 24394 8984 24400 9036
rect 24452 9024 24458 9036
rect 24673 9027 24731 9033
rect 24673 9024 24685 9027
rect 24452 8996 24685 9024
rect 24452 8984 24458 8996
rect 24673 8993 24685 8996
rect 24719 9024 24731 9027
rect 24857 9027 24915 9033
rect 24857 9024 24869 9027
rect 24719 8996 24869 9024
rect 24719 8993 24731 8996
rect 24673 8987 24731 8993
rect 24857 8993 24869 8996
rect 24903 9024 24915 9027
rect 25409 9027 25467 9033
rect 25409 9024 25421 9027
rect 24903 8996 25421 9024
rect 24903 8993 24915 8996
rect 24857 8987 24915 8993
rect 25409 8993 25421 8996
rect 25455 9024 25467 9027
rect 25590 9024 25596 9036
rect 25455 8996 25596 9024
rect 25455 8993 25467 8996
rect 25409 8987 25467 8993
rect 25590 8984 25596 8996
rect 25648 8984 25654 9036
rect 28368 9033 28396 9064
rect 30006 9052 30012 9064
rect 30064 9092 30070 9104
rect 30745 9095 30803 9101
rect 30745 9092 30757 9095
rect 30064 9064 30757 9092
rect 30064 9052 30070 9064
rect 30745 9061 30757 9064
rect 30791 9061 30803 9095
rect 32416 9092 32444 9132
rect 32861 9129 32873 9163
rect 32907 9160 32919 9163
rect 33045 9163 33103 9169
rect 33045 9160 33057 9163
rect 32907 9132 33057 9160
rect 32907 9129 32919 9132
rect 32861 9123 32919 9129
rect 33045 9129 33057 9132
rect 33091 9160 33103 9163
rect 33502 9160 33508 9172
rect 33091 9132 33508 9160
rect 33091 9129 33103 9132
rect 33045 9123 33103 9129
rect 33502 9120 33508 9132
rect 33560 9120 33566 9172
rect 34057 9163 34115 9169
rect 34057 9129 34069 9163
rect 34103 9160 34115 9163
rect 36354 9160 36360 9172
rect 34103 9132 36360 9160
rect 34103 9129 34115 9132
rect 34057 9123 34115 9129
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 37090 9160 37096 9172
rect 36648 9132 37096 9160
rect 36648 9092 36676 9132
rect 37090 9120 37096 9132
rect 37148 9120 37154 9172
rect 32416 9064 36676 9092
rect 36725 9095 36783 9101
rect 30745 9055 30803 9061
rect 36725 9061 36737 9095
rect 36771 9092 36783 9095
rect 39942 9092 39948 9104
rect 36771 9064 39948 9092
rect 36771 9061 36783 9064
rect 36725 9055 36783 9061
rect 39942 9052 39948 9064
rect 40000 9052 40006 9104
rect 28353 9027 28411 9033
rect 28353 8993 28365 9027
rect 28399 8993 28411 9027
rect 31754 9024 31760 9036
rect 28353 8987 28411 8993
rect 28460 8996 31760 9024
rect 24394 8888 24400 8900
rect 20548 8860 22508 8888
rect 23322 8860 24400 8888
rect 20548 8820 20576 8860
rect 24394 8848 24400 8860
rect 24452 8848 24458 8900
rect 16040 8792 20576 8820
rect 21821 8823 21879 8829
rect 21821 8789 21833 8823
rect 21867 8820 21879 8823
rect 22186 8820 22192 8832
rect 21867 8792 22192 8820
rect 21867 8789 21879 8792
rect 21821 8783 21879 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 27798 8780 27804 8832
rect 27856 8820 27862 8832
rect 28460 8829 28488 8996
rect 31754 8984 31760 8996
rect 31812 8984 31818 9036
rect 32122 8984 32128 9036
rect 32180 9024 32186 9036
rect 32493 9027 32551 9033
rect 32493 9024 32505 9027
rect 32180 8996 32505 9024
rect 32180 8984 32186 8996
rect 32493 8993 32505 8996
rect 32539 8993 32551 9027
rect 32493 8987 32551 8993
rect 33505 9027 33563 9033
rect 33505 8993 33517 9027
rect 33551 8993 33563 9027
rect 33505 8987 33563 8993
rect 30650 8916 30656 8968
rect 30708 8956 30714 8968
rect 31110 8956 31116 8968
rect 30708 8928 31116 8956
rect 30708 8916 30714 8928
rect 31110 8916 31116 8928
rect 31168 8916 31174 8968
rect 32582 8916 32588 8968
rect 32640 8956 32646 8968
rect 33520 8956 33548 8987
rect 33594 8984 33600 9036
rect 33652 8984 33658 9036
rect 34054 8984 34060 9036
rect 34112 9024 34118 9036
rect 34977 9027 35035 9033
rect 34977 9024 34989 9027
rect 34112 8996 34989 9024
rect 34112 8984 34118 8996
rect 34977 8993 34989 8996
rect 35023 8993 35035 9027
rect 34977 8987 35035 8993
rect 35158 8984 35164 9036
rect 35216 9024 35222 9036
rect 49145 9027 49203 9033
rect 35216 8996 37688 9024
rect 35216 8984 35222 8996
rect 34238 8956 34244 8968
rect 32640 8928 34244 8956
rect 32640 8916 32646 8928
rect 34238 8916 34244 8928
rect 34296 8916 34302 8968
rect 34514 8916 34520 8968
rect 34572 8956 34578 8968
rect 37660 8965 37688 8996
rect 49145 8993 49157 9027
rect 49191 9024 49203 9027
rect 49326 9024 49332 9036
rect 49191 8996 49332 9024
rect 49191 8993 49203 8996
rect 49145 8987 49203 8993
rect 49326 8984 49332 8996
rect 49384 8984 49390 9036
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 34572 8928 36553 8956
rect 34572 8916 34578 8928
rect 36541 8925 36553 8928
rect 36587 8925 36599 8959
rect 36541 8919 36599 8925
rect 37645 8959 37703 8965
rect 37645 8925 37657 8959
rect 37691 8925 37703 8959
rect 39853 8959 39911 8965
rect 39853 8956 39865 8959
rect 37645 8919 37703 8925
rect 39316 8928 39865 8956
rect 28537 8891 28595 8897
rect 28537 8857 28549 8891
rect 28583 8888 28595 8891
rect 29733 8891 29791 8897
rect 29733 8888 29745 8891
rect 28583 8860 29745 8888
rect 28583 8857 28595 8860
rect 28537 8851 28595 8857
rect 29733 8857 29745 8860
rect 29779 8857 29791 8891
rect 32217 8891 32275 8897
rect 29733 8851 29791 8857
rect 30116 8860 30880 8888
rect 28445 8823 28503 8829
rect 28445 8820 28457 8823
rect 27856 8792 28457 8820
rect 27856 8780 27862 8792
rect 28445 8789 28457 8792
rect 28491 8789 28503 8823
rect 28445 8783 28503 8789
rect 28905 8823 28963 8829
rect 28905 8789 28917 8823
rect 28951 8820 28963 8823
rect 30116 8820 30144 8860
rect 28951 8792 30144 8820
rect 30285 8823 30343 8829
rect 28951 8789 28963 8792
rect 28905 8783 28963 8789
rect 30285 8789 30297 8823
rect 30331 8820 30343 8823
rect 30650 8820 30656 8832
rect 30331 8792 30656 8820
rect 30331 8789 30343 8792
rect 30285 8783 30343 8789
rect 30650 8780 30656 8792
rect 30708 8780 30714 8832
rect 30852 8820 30880 8860
rect 32217 8857 32229 8891
rect 32263 8888 32275 8891
rect 34054 8888 34060 8900
rect 32263 8860 34060 8888
rect 32263 8857 32275 8860
rect 32217 8851 32275 8857
rect 34054 8848 34060 8860
rect 34112 8848 34118 8900
rect 34146 8848 34152 8900
rect 34204 8888 34210 8900
rect 35253 8891 35311 8897
rect 35253 8888 35265 8891
rect 34204 8860 35265 8888
rect 34204 8848 34210 8860
rect 35253 8857 35265 8860
rect 35299 8857 35311 8891
rect 35253 8851 35311 8857
rect 37090 8848 37096 8900
rect 37148 8888 37154 8900
rect 39316 8897 39344 8928
rect 39853 8925 39865 8928
rect 39899 8925 39911 8959
rect 39853 8919 39911 8925
rect 47026 8916 47032 8968
rect 47084 8956 47090 8968
rect 47949 8959 48007 8965
rect 47949 8956 47961 8959
rect 47084 8928 47961 8956
rect 47084 8916 47090 8928
rect 47949 8925 47961 8928
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 39301 8891 39359 8897
rect 39301 8888 39313 8891
rect 37148 8860 39313 8888
rect 37148 8848 37154 8860
rect 39301 8857 39313 8860
rect 39347 8857 39359 8891
rect 39301 8851 39359 8857
rect 39485 8891 39543 8897
rect 39485 8857 39497 8891
rect 39531 8888 39543 8891
rect 47578 8888 47584 8900
rect 39531 8860 47584 8888
rect 39531 8857 39543 8860
rect 39485 8851 39543 8857
rect 47578 8848 47584 8860
rect 47636 8848 47642 8900
rect 31938 8820 31944 8832
rect 30852 8792 31944 8820
rect 31938 8780 31944 8792
rect 31996 8780 32002 8832
rect 33686 8780 33692 8832
rect 33744 8820 33750 8832
rect 34333 8823 34391 8829
rect 34333 8820 34345 8823
rect 33744 8792 34345 8820
rect 33744 8780 33750 8792
rect 34333 8789 34345 8792
rect 34379 8789 34391 8823
rect 34333 8783 34391 8789
rect 34606 8780 34612 8832
rect 34664 8820 34670 8832
rect 35161 8823 35219 8829
rect 35161 8820 35173 8823
rect 34664 8792 35173 8820
rect 34664 8780 34670 8792
rect 35161 8789 35173 8792
rect 35207 8789 35219 8823
rect 35161 8783 35219 8789
rect 35618 8780 35624 8832
rect 35676 8780 35682 8832
rect 37829 8823 37887 8829
rect 37829 8789 37841 8823
rect 37875 8820 37887 8823
rect 39758 8820 39764 8832
rect 37875 8792 39764 8820
rect 37875 8789 37887 8792
rect 37829 8783 37887 8789
rect 39758 8780 39764 8792
rect 39816 8780 39822 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 15194 8616 15200 8628
rect 12768 8588 15200 8616
rect 12768 8576 12774 8588
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 13648 8489 13676 8588
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 15795 8588 16221 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 16209 8585 16221 8588
rect 16255 8616 16267 8619
rect 17402 8616 17408 8628
rect 16255 8588 17408 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 13906 8508 13912 8560
rect 13964 8508 13970 8560
rect 15286 8548 15292 8560
rect 15134 8520 15292 8548
rect 15286 8508 15292 8520
rect 15344 8548 15350 8560
rect 15764 8548 15792 8579
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 19886 8616 19892 8628
rect 19751 8588 19892 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21192 8588 22017 8616
rect 15344 8520 15792 8548
rect 15344 8508 15350 8520
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17126 8548 17132 8560
rect 16816 8520 17132 8548
rect 16816 8508 16822 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 18414 8548 18420 8560
rect 18354 8520 18420 8548
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 20438 8508 20444 8560
rect 20496 8508 20502 8560
rect 21192 8557 21220 8588
rect 21177 8551 21235 8557
rect 21177 8517 21189 8551
rect 21223 8517 21235 8551
rect 21177 8511 21235 8517
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 16482 8480 16488 8492
rect 15252 8452 16488 8480
rect 15252 8440 15258 8452
rect 16482 8440 16488 8452
rect 16540 8480 16546 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16540 8452 16865 8480
rect 16540 8440 16546 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 2406 8372 2412 8424
rect 2464 8372 2470 8424
rect 15102 8372 15108 8424
rect 15160 8412 15166 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15160 8384 15393 8412
rect 15160 8372 15166 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 17828 8384 19073 8412
rect 17828 8372 17834 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 21450 8372 21456 8424
rect 21508 8372 21514 8424
rect 21928 8344 21956 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 24121 8619 24179 8625
rect 22005 8579 22063 8585
rect 22388 8588 23152 8616
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 22388 8480 22416 8588
rect 23124 8548 23152 8588
rect 24121 8585 24133 8619
rect 24167 8616 24179 8619
rect 24394 8616 24400 8628
rect 24167 8588 24400 8616
rect 24167 8585 24179 8588
rect 24121 8579 24179 8585
rect 24136 8548 24164 8579
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 31110 8576 31116 8628
rect 31168 8616 31174 8628
rect 31389 8619 31447 8625
rect 31389 8616 31401 8619
rect 31168 8588 31401 8616
rect 31168 8576 31174 8588
rect 31389 8585 31401 8588
rect 31435 8585 31447 8619
rect 31389 8579 31447 8585
rect 31757 8619 31815 8625
rect 31757 8585 31769 8619
rect 31803 8616 31815 8619
rect 33870 8616 33876 8628
rect 31803 8588 33876 8616
rect 31803 8585 31815 8588
rect 31757 8579 31815 8585
rect 33870 8576 33876 8588
rect 33928 8576 33934 8628
rect 34054 8576 34060 8628
rect 34112 8576 34118 8628
rect 34238 8576 34244 8628
rect 34296 8616 34302 8628
rect 34333 8619 34391 8625
rect 34333 8616 34345 8619
rect 34296 8588 34345 8616
rect 34296 8576 34302 8588
rect 34333 8585 34345 8588
rect 34379 8585 34391 8619
rect 34333 8579 34391 8585
rect 37645 8619 37703 8625
rect 37645 8585 37657 8619
rect 37691 8616 37703 8619
rect 41414 8616 41420 8628
rect 37691 8588 41420 8616
rect 37691 8585 37703 8588
rect 37645 8579 37703 8585
rect 41414 8576 41420 8588
rect 41472 8576 41478 8628
rect 23046 8520 24164 8548
rect 29086 8508 29092 8560
rect 29144 8508 29150 8560
rect 30650 8548 30656 8560
rect 30314 8520 30656 8548
rect 30650 8508 30656 8520
rect 30708 8508 30714 8560
rect 31938 8548 31944 8560
rect 31312 8520 31944 8548
rect 22060 8466 22416 8480
rect 23753 8483 23811 8489
rect 22060 8452 22402 8466
rect 22060 8440 22066 8452
rect 23753 8449 23765 8483
rect 23799 8480 23811 8483
rect 24026 8480 24032 8492
rect 23799 8452 24032 8480
rect 23799 8449 23811 8452
rect 23753 8443 23811 8449
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 31312 8480 31340 8520
rect 31938 8508 31944 8520
rect 31996 8548 32002 8560
rect 32582 8548 32588 8560
rect 31996 8520 32588 8548
rect 31996 8508 32002 8520
rect 32582 8508 32588 8520
rect 32640 8508 32646 8560
rect 34698 8548 34704 8560
rect 33810 8520 34704 8548
rect 34698 8508 34704 8520
rect 34756 8508 34762 8560
rect 35618 8508 35624 8560
rect 35676 8548 35682 8560
rect 35676 8520 38976 8548
rect 35676 8508 35682 8520
rect 31220 8452 31340 8480
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 23477 8415 23535 8421
rect 23477 8412 23489 8415
rect 22152 8384 23489 8412
rect 22152 8372 22158 8384
rect 23477 8381 23489 8384
rect 23523 8381 23535 8415
rect 23477 8375 23535 8381
rect 28810 8372 28816 8424
rect 28868 8412 28874 8424
rect 29178 8412 29184 8424
rect 28868 8384 29184 8412
rect 28868 8372 28874 8384
rect 29178 8372 29184 8384
rect 29236 8372 29242 8424
rect 31220 8421 31248 8452
rect 31754 8440 31760 8492
rect 31812 8480 31818 8492
rect 32030 8480 32036 8492
rect 31812 8452 32036 8480
rect 31812 8440 31818 8452
rect 32030 8440 32036 8452
rect 32088 8440 32094 8492
rect 32122 8440 32128 8492
rect 32180 8480 32186 8492
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 32180 8452 32321 8480
rect 32180 8440 32186 8452
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 33796 8452 37412 8480
rect 31205 8415 31263 8421
rect 31205 8381 31217 8415
rect 31251 8381 31263 8415
rect 31205 8375 31263 8381
rect 31294 8372 31300 8424
rect 31352 8372 31358 8424
rect 32214 8372 32220 8424
rect 32272 8412 32278 8424
rect 32585 8415 32643 8421
rect 32585 8412 32597 8415
rect 32272 8384 32597 8412
rect 32272 8372 32278 8384
rect 32585 8381 32597 8384
rect 32631 8412 32643 8415
rect 32674 8412 32680 8424
rect 32631 8384 32680 8412
rect 32631 8381 32643 8384
rect 32585 8375 32643 8381
rect 32674 8372 32680 8384
rect 32732 8372 32738 8424
rect 32950 8372 32956 8424
rect 33008 8412 33014 8424
rect 33796 8412 33824 8452
rect 33008 8384 33824 8412
rect 33008 8372 33014 8384
rect 33870 8372 33876 8424
rect 33928 8412 33934 8424
rect 36446 8412 36452 8424
rect 33928 8384 36452 8412
rect 33928 8372 33934 8384
rect 36446 8372 36452 8384
rect 36504 8372 36510 8424
rect 37384 8412 37412 8452
rect 37458 8440 37464 8492
rect 37516 8440 37522 8492
rect 38948 8489 38976 8520
rect 39758 8508 39764 8560
rect 39816 8548 39822 8560
rect 44177 8551 44235 8557
rect 44177 8548 44189 8551
rect 39816 8520 44189 8548
rect 39816 8508 39822 8520
rect 44177 8517 44189 8520
rect 44223 8517 44235 8551
rect 44177 8511 44235 8517
rect 44361 8551 44419 8557
rect 44361 8517 44373 8551
rect 44407 8548 44419 8551
rect 47854 8548 47860 8560
rect 44407 8520 47860 8548
rect 44407 8517 44419 8520
rect 44361 8511 44419 8517
rect 47854 8508 47860 8520
rect 47912 8508 47918 8560
rect 49142 8508 49148 8560
rect 49200 8508 49206 8560
rect 38933 8483 38991 8489
rect 38933 8449 38945 8483
rect 38979 8449 38991 8483
rect 38933 8443 38991 8449
rect 40310 8440 40316 8492
rect 40368 8480 40374 8492
rect 40773 8483 40831 8489
rect 40773 8480 40785 8483
rect 40368 8452 40785 8480
rect 40368 8440 40374 8452
rect 40773 8449 40785 8452
rect 40819 8449 40831 8483
rect 40773 8443 40831 8449
rect 45830 8440 45836 8492
rect 45888 8440 45894 8492
rect 46750 8440 46756 8492
rect 46808 8480 46814 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46808 8452 47961 8480
rect 46808 8440 46814 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 38746 8412 38752 8424
rect 37384 8384 38752 8412
rect 38746 8372 38752 8384
rect 38804 8372 38810 8424
rect 40497 8415 40555 8421
rect 40497 8381 40509 8415
rect 40543 8412 40555 8415
rect 40543 8384 45554 8412
rect 40543 8381 40555 8384
rect 40497 8375 40555 8381
rect 22462 8344 22468 8356
rect 21928 8316 22468 8344
rect 22462 8304 22468 8316
rect 22520 8304 22526 8356
rect 30561 8347 30619 8353
rect 30561 8313 30573 8347
rect 30607 8344 30619 8347
rect 31846 8344 31852 8356
rect 30607 8316 31852 8344
rect 30607 8313 30619 8316
rect 30561 8307 30619 8313
rect 31846 8304 31852 8316
rect 31904 8304 31910 8356
rect 33594 8304 33600 8356
rect 33652 8344 33658 8356
rect 34517 8347 34575 8353
rect 34517 8344 34529 8347
rect 33652 8316 34529 8344
rect 33652 8304 33658 8316
rect 34517 8313 34529 8316
rect 34563 8344 34575 8347
rect 38930 8344 38936 8356
rect 34563 8316 38936 8344
rect 34563 8313 34575 8316
rect 34517 8307 34575 8313
rect 38930 8304 38936 8316
rect 38988 8304 38994 8356
rect 39117 8347 39175 8353
rect 39117 8313 39129 8347
rect 39163 8344 39175 8347
rect 44910 8344 44916 8356
rect 39163 8316 44916 8344
rect 39163 8313 39175 8316
rect 39117 8307 39175 8313
rect 44910 8304 44916 8316
rect 44968 8304 44974 8356
rect 45526 8344 45554 8384
rect 46842 8372 46848 8424
rect 46900 8372 46906 8424
rect 47670 8344 47676 8356
rect 45526 8316 47676 8344
rect 47670 8304 47676 8316
rect 47728 8304 47734 8356
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 1360 8044 2145 8072
rect 1360 8032 1366 8044
rect 2133 8041 2145 8044
rect 2179 8072 2191 8075
rect 2406 8072 2412 8084
rect 2179 8044 2412 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 18564 8044 18981 8072
rect 18564 8032 18570 8044
rect 18969 8041 18981 8044
rect 19015 8041 19027 8075
rect 18969 8035 19027 8041
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22005 8075 22063 8081
rect 22005 8072 22017 8075
rect 21968 8044 22017 8072
rect 21968 8032 21974 8044
rect 22005 8041 22017 8044
rect 22051 8041 22063 8075
rect 22005 8035 22063 8041
rect 30377 8075 30435 8081
rect 30377 8041 30389 8075
rect 30423 8072 30435 8075
rect 30558 8072 30564 8084
rect 30423 8044 30564 8072
rect 30423 8041 30435 8044
rect 30377 8035 30435 8041
rect 30558 8032 30564 8044
rect 30616 8032 30622 8084
rect 31757 8075 31815 8081
rect 31757 8041 31769 8075
rect 31803 8072 31815 8075
rect 34146 8072 34152 8084
rect 31803 8044 34152 8072
rect 31803 8041 31815 8044
rect 31757 8035 31815 8041
rect 34146 8032 34152 8044
rect 34204 8032 34210 8084
rect 15749 8007 15807 8013
rect 15749 7973 15761 8007
rect 15795 8004 15807 8007
rect 18874 8004 18880 8016
rect 15795 7976 18880 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 18874 7964 18880 7976
rect 18932 7964 18938 8016
rect 33045 8007 33103 8013
rect 33045 7973 33057 8007
rect 33091 8004 33103 8007
rect 39022 8004 39028 8016
rect 33091 7976 39028 8004
rect 33091 7973 33103 7976
rect 33045 7967 33103 7973
rect 39022 7964 39028 7976
rect 39080 7964 39086 8016
rect 16758 7896 16764 7948
rect 16816 7896 16822 7948
rect 16942 7896 16948 7948
rect 17000 7896 17006 7948
rect 18049 7939 18107 7945
rect 18049 7905 18061 7939
rect 18095 7936 18107 7939
rect 18598 7936 18604 7948
rect 18095 7908 18604 7936
rect 18095 7905 18107 7908
rect 18049 7899 18107 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 19944 7908 20913 7936
rect 19944 7896 19950 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7936 22707 7939
rect 23658 7936 23664 7948
rect 22695 7908 23664 7936
rect 22695 7905 22707 7908
rect 22649 7899 22707 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 29914 7896 29920 7948
rect 29972 7896 29978 7948
rect 31205 7939 31263 7945
rect 31205 7905 31217 7939
rect 31251 7936 31263 7939
rect 32214 7936 32220 7948
rect 31251 7908 32220 7936
rect 31251 7905 31263 7908
rect 31205 7899 31263 7905
rect 32214 7896 32220 7908
rect 32272 7896 32278 7948
rect 32493 7939 32551 7945
rect 32493 7905 32505 7939
rect 32539 7936 32551 7939
rect 33413 7939 33471 7945
rect 33413 7936 33425 7939
rect 32539 7908 33425 7936
rect 32539 7905 32551 7908
rect 32493 7899 32551 7905
rect 33413 7905 33425 7908
rect 33459 7936 33471 7939
rect 34790 7936 34796 7948
rect 33459 7908 34796 7936
rect 33459 7905 33471 7908
rect 33413 7899 33471 7905
rect 34790 7896 34796 7908
rect 34848 7896 34854 7948
rect 49145 7939 49203 7945
rect 49145 7905 49157 7939
rect 49191 7936 49203 7939
rect 49234 7936 49240 7948
rect 49191 7908 49240 7936
rect 49191 7905 49203 7908
rect 49145 7899 49203 7905
rect 49234 7896 49240 7908
rect 49292 7896 49298 7948
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 1360 7840 1593 7868
rect 1360 7828 1366 7840
rect 1581 7837 1593 7840
rect 1627 7868 1639 7871
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1627 7840 2329 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 12434 7868 12440 7880
rect 2740 7840 12440 7868
rect 2740 7828 2746 7840
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 14976 7840 15577 7868
rect 14976 7828 14982 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 17034 7828 17040 7880
rect 17092 7828 17098 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 17236 7840 18153 7868
rect 13722 7800 13728 7812
rect 1780 7772 13728 7800
rect 1780 7741 1808 7772
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 16390 7760 16396 7812
rect 16448 7800 16454 7812
rect 17236 7800 17264 7840
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 21450 7868 21456 7880
rect 21223 7840 21456 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 16448 7772 17264 7800
rect 17420 7772 18245 7800
rect 16448 7760 16454 7772
rect 17420 7741 17448 7772
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 19610 7800 19616 7812
rect 18233 7763 18291 7769
rect 18616 7772 19616 7800
rect 18616 7741 18644 7772
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 20438 7760 20444 7812
rect 20496 7800 20502 7812
rect 20496 7772 20576 7800
rect 20496 7760 20502 7772
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7701 1823 7735
rect 1765 7695 1823 7701
rect 17405 7735 17463 7741
rect 17405 7701 17417 7735
rect 17451 7701 17463 7735
rect 17405 7695 17463 7701
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7701 18659 7735
rect 20548 7732 20576 7772
rect 20990 7760 20996 7812
rect 21048 7800 21054 7812
rect 21192 7800 21220 7831
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22244 7840 22385 7868
rect 22244 7828 22250 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 30558 7828 30564 7880
rect 30616 7868 30622 7880
rect 31297 7871 31355 7877
rect 31297 7868 31309 7871
rect 30616 7840 31309 7868
rect 30616 7828 30622 7840
rect 31297 7837 31309 7840
rect 31343 7837 31355 7871
rect 31297 7831 31355 7837
rect 32677 7871 32735 7877
rect 32677 7837 32689 7871
rect 32723 7868 32735 7871
rect 32766 7868 32772 7880
rect 32723 7840 32772 7868
rect 32723 7837 32735 7840
rect 32677 7831 32735 7837
rect 32766 7828 32772 7840
rect 32824 7828 32830 7880
rect 38746 7828 38752 7880
rect 38804 7868 38810 7880
rect 39209 7871 39267 7877
rect 39209 7868 39221 7871
rect 38804 7840 39221 7868
rect 38804 7828 38810 7840
rect 39209 7837 39221 7840
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 47118 7828 47124 7880
rect 47176 7868 47182 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 47176 7840 47961 7868
rect 47176 7828 47182 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 30466 7800 30472 7812
rect 21048 7772 21220 7800
rect 22388 7772 30472 7800
rect 21048 7760 21054 7772
rect 22388 7744 22416 7772
rect 30466 7760 30472 7772
rect 30524 7760 30530 7812
rect 37553 7803 37611 7809
rect 37553 7800 37565 7803
rect 30576 7772 37565 7800
rect 21450 7732 21456 7744
rect 20548 7704 21456 7732
rect 18601 7695 18659 7701
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 21634 7692 21640 7744
rect 21692 7692 21698 7744
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 23017 7735 23075 7741
rect 23017 7732 23029 7735
rect 22520 7704 23029 7732
rect 22520 7692 22526 7704
rect 23017 7701 23029 7704
rect 23063 7732 23075 7735
rect 25682 7732 25688 7744
rect 23063 7704 25688 7732
rect 23063 7701 23075 7704
rect 23017 7695 23075 7701
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 27246 7692 27252 7744
rect 27304 7732 27310 7744
rect 30576 7732 30604 7772
rect 37553 7769 37565 7772
rect 37599 7800 37611 7803
rect 38013 7803 38071 7809
rect 38013 7800 38025 7803
rect 37599 7772 38025 7800
rect 37599 7769 37611 7772
rect 37553 7763 37611 7769
rect 38013 7769 38025 7772
rect 38059 7769 38071 7803
rect 38013 7763 38071 7769
rect 38933 7803 38991 7809
rect 38933 7769 38945 7803
rect 38979 7800 38991 7803
rect 41322 7800 41328 7812
rect 38979 7772 41328 7800
rect 38979 7769 38991 7772
rect 38933 7763 38991 7769
rect 41322 7760 41328 7772
rect 41380 7760 41386 7812
rect 27304 7704 30604 7732
rect 27304 7692 27310 7704
rect 30650 7692 30656 7744
rect 30708 7692 30714 7744
rect 31386 7692 31392 7744
rect 31444 7692 31450 7744
rect 32582 7692 32588 7744
rect 32640 7692 32646 7744
rect 38105 7735 38163 7741
rect 38105 7701 38117 7735
rect 38151 7732 38163 7735
rect 38654 7732 38660 7744
rect 38151 7704 38660 7732
rect 38151 7701 38163 7704
rect 38105 7695 38163 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 17920 7500 18337 7528
rect 17920 7488 17926 7500
rect 18325 7497 18337 7500
rect 18371 7528 18383 7531
rect 18414 7528 18420 7540
rect 18371 7500 18420 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 18414 7488 18420 7500
rect 18472 7528 18478 7540
rect 18785 7531 18843 7537
rect 18785 7528 18797 7531
rect 18472 7500 18797 7528
rect 18472 7488 18478 7500
rect 18785 7497 18797 7500
rect 18831 7528 18843 7531
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 18831 7500 19073 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 19061 7497 19073 7500
rect 19107 7528 19119 7531
rect 20438 7528 20444 7540
rect 19107 7500 20444 7528
rect 19107 7497 19119 7500
rect 19061 7491 19119 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 20680 7500 22017 7528
rect 20680 7488 20686 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 22278 7488 22284 7540
rect 22336 7528 22342 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22336 7500 22477 7528
rect 22336 7488 22342 7500
rect 22465 7497 22477 7500
rect 22511 7528 22523 7531
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22511 7500 23029 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 31110 7488 31116 7540
rect 31168 7488 31174 7540
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 32309 7531 32367 7537
rect 32309 7528 32321 7531
rect 31444 7500 32321 7528
rect 31444 7488 31450 7500
rect 32309 7497 32321 7500
rect 32355 7497 32367 7531
rect 32309 7491 32367 7497
rect 38654 7488 38660 7540
rect 38712 7528 38718 7540
rect 47302 7528 47308 7540
rect 38712 7500 47308 7528
rect 38712 7488 38718 7500
rect 47302 7488 47308 7500
rect 47360 7488 47366 7540
rect 31938 7420 31944 7472
rect 31996 7420 32002 7472
rect 37369 7463 37427 7469
rect 37369 7460 37381 7463
rect 32048 7432 37381 7460
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1360 7364 1593 7392
rect 1360 7352 1366 7364
rect 1581 7361 1593 7364
rect 1627 7392 1639 7395
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1627 7364 2145 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 27614 7352 27620 7404
rect 27672 7392 27678 7404
rect 32048 7392 32076 7432
rect 37369 7429 37381 7432
rect 37415 7460 37427 7463
rect 37829 7463 37887 7469
rect 37829 7460 37841 7463
rect 37415 7432 37841 7460
rect 37415 7429 37427 7432
rect 37369 7423 37427 7429
rect 37829 7429 37841 7432
rect 37875 7429 37887 7463
rect 37829 7423 37887 7429
rect 44910 7420 44916 7472
rect 44968 7420 44974 7472
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 49326 7460 49332 7472
rect 49191 7432 49332 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 49326 7420 49332 7432
rect 49384 7420 49390 7472
rect 27672 7364 32076 7392
rect 27672 7352 27678 7364
rect 33318 7352 33324 7404
rect 33376 7392 33382 7404
rect 38565 7395 38623 7401
rect 38565 7392 38577 7395
rect 33376 7364 38577 7392
rect 33376 7352 33382 7364
rect 38565 7361 38577 7364
rect 38611 7392 38623 7395
rect 39025 7395 39083 7401
rect 39025 7392 39037 7395
rect 38611 7364 39037 7392
rect 38611 7361 38623 7364
rect 38565 7355 38623 7361
rect 39025 7361 39037 7364
rect 39071 7361 39083 7395
rect 39025 7355 39083 7361
rect 46934 7352 46940 7404
rect 46992 7392 46998 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 46992 7364 47961 7392
rect 46992 7352 46998 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 22554 7284 22560 7336
rect 22612 7284 22618 7336
rect 30466 7284 30472 7336
rect 30524 7324 30530 7336
rect 31294 7324 31300 7336
rect 30524 7296 31300 7324
rect 30524 7284 30530 7296
rect 31294 7284 31300 7296
rect 31352 7324 31358 7336
rect 38470 7324 38476 7336
rect 31352 7296 38476 7324
rect 31352 7284 31358 7296
rect 38470 7284 38476 7296
rect 38528 7284 38534 7336
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 18782 7256 18788 7268
rect 1811 7228 18788 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 20714 7216 20720 7268
rect 20772 7256 20778 7268
rect 21634 7256 21640 7268
rect 20772 7228 21640 7256
rect 20772 7216 20778 7228
rect 21634 7216 21640 7228
rect 21692 7256 21698 7268
rect 22646 7256 22652 7268
rect 21692 7228 22652 7256
rect 21692 7216 21698 7228
rect 22646 7216 22652 7228
rect 22704 7256 22710 7268
rect 32582 7256 32588 7268
rect 22704 7228 32588 7256
rect 22704 7216 22710 7228
rect 32582 7216 32588 7228
rect 32640 7256 32646 7268
rect 32769 7259 32827 7265
rect 32769 7256 32781 7259
rect 32640 7228 32781 7256
rect 32640 7216 32646 7228
rect 32769 7225 32781 7228
rect 32815 7256 32827 7259
rect 37274 7256 37280 7268
rect 32815 7228 37280 7256
rect 32815 7225 32827 7228
rect 32769 7219 32827 7225
rect 37274 7216 37280 7228
rect 37332 7216 37338 7268
rect 38749 7259 38807 7265
rect 38749 7225 38761 7259
rect 38795 7256 38807 7259
rect 45097 7259 45155 7265
rect 38795 7228 42104 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 21177 7191 21235 7197
rect 21177 7157 21189 7191
rect 21223 7188 21235 7191
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 21223 7160 21373 7188
rect 21223 7157 21235 7160
rect 21177 7151 21235 7157
rect 21361 7157 21373 7160
rect 21407 7188 21419 7191
rect 21450 7188 21456 7200
rect 21407 7160 21456 7188
rect 21407 7157 21419 7160
rect 21361 7151 21419 7157
rect 21450 7148 21456 7160
rect 21508 7188 21514 7200
rect 21545 7191 21603 7197
rect 21545 7188 21557 7191
rect 21508 7160 21557 7188
rect 21508 7148 21514 7160
rect 21545 7157 21557 7160
rect 21591 7188 21603 7191
rect 22002 7188 22008 7200
rect 21591 7160 22008 7188
rect 21591 7157 21603 7160
rect 21545 7151 21603 7157
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 37918 7148 37924 7200
rect 37976 7148 37982 7200
rect 42076 7188 42104 7228
rect 45097 7225 45109 7259
rect 45143 7256 45155 7259
rect 47762 7256 47768 7268
rect 45143 7228 47768 7256
rect 45143 7225 45155 7228
rect 45097 7219 45155 7225
rect 47762 7216 47768 7228
rect 47820 7216 47826 7268
rect 45830 7188 45836 7200
rect 42076 7160 45836 7188
rect 45830 7148 45836 7160
rect 45888 7148 45894 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 37918 6876 37924 6928
rect 37976 6916 37982 6928
rect 46934 6916 46940 6928
rect 37976 6888 46940 6916
rect 37976 6876 37982 6888
rect 46934 6876 46940 6888
rect 46992 6876 46998 6928
rect 15654 6808 15660 6860
rect 15712 6848 15718 6860
rect 21821 6851 21879 6857
rect 21821 6848 21833 6851
rect 15712 6820 21833 6848
rect 15712 6808 15718 6820
rect 21821 6817 21833 6820
rect 21867 6848 21879 6851
rect 22370 6848 22376 6860
rect 21867 6820 22376 6848
rect 21867 6817 21879 6820
rect 21821 6811 21879 6817
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 49142 6808 49148 6860
rect 49200 6808 49206 6860
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 2317 6783 2375 6789
rect 2317 6780 2329 6783
rect 1360 6752 2329 6780
rect 1360 6740 1366 6752
rect 2317 6749 2329 6752
rect 2363 6780 2375 6783
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2363 6752 2789 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 15988 6752 17693 6780
rect 15988 6740 15994 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 41322 6740 41328 6792
rect 41380 6780 41386 6792
rect 46109 6783 46167 6789
rect 46109 6780 46121 6783
rect 41380 6752 46121 6780
rect 41380 6740 41386 6752
rect 46109 6749 46121 6752
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 47854 6740 47860 6792
rect 47912 6780 47918 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47912 6752 47961 6780
rect 47912 6740 47918 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 1210 6672 1216 6724
rect 1268 6712 1274 6724
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 1268 6684 1685 6712
rect 1268 6672 1274 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 10594 6712 10600 6724
rect 1673 6675 1731 6681
rect 2516 6684 10600 6712
rect 1762 6604 1768 6656
rect 1820 6604 1826 6656
rect 2516 6653 2544 6684
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 47305 6715 47363 6721
rect 47305 6681 47317 6715
rect 47351 6712 47363 6715
rect 48682 6712 48688 6724
rect 47351 6684 48688 6712
rect 47351 6681 47363 6684
rect 47305 6675 47363 6681
rect 48682 6672 48688 6684
rect 48740 6672 48746 6724
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 17865 6647 17923 6653
rect 17865 6613 17877 6647
rect 17911 6644 17923 6647
rect 19242 6644 19248 6656
rect 17911 6616 19248 6644
rect 17911 6613 17923 6616
rect 17865 6607 17923 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19797 6647 19855 6653
rect 19797 6613 19809 6647
rect 19843 6644 19855 6647
rect 21726 6644 21732 6656
rect 19843 6616 21732 6644
rect 19843 6613 19855 6616
rect 19797 6607 19855 6613
rect 21726 6604 21732 6616
rect 21784 6604 21790 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1268 6412 2145 6440
rect 1268 6400 1274 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 27522 6332 27528 6384
rect 27580 6372 27586 6384
rect 36814 6372 36820 6384
rect 27580 6344 36820 6372
rect 27580 6332 27586 6344
rect 36814 6332 36820 6344
rect 36872 6332 36878 6384
rect 41414 6332 41420 6384
rect 41472 6372 41478 6384
rect 43993 6375 44051 6381
rect 43993 6372 44005 6375
rect 41472 6344 44005 6372
rect 41472 6332 41478 6344
rect 43993 6341 44005 6344
rect 44039 6341 44051 6375
rect 43993 6335 44051 6341
rect 49145 6375 49203 6381
rect 49145 6341 49157 6375
rect 49191 6372 49203 6375
rect 49418 6372 49424 6384
rect 49191 6344 49424 6372
rect 49191 6341 49203 6344
rect 49145 6335 49203 6341
rect 49418 6332 49424 6344
rect 49476 6332 49482 6384
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1596 6236 1624 6267
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 27798 6304 27804 6316
rect 1820 6276 27804 6304
rect 1820 6264 1826 6276
rect 27798 6264 27804 6276
rect 27856 6264 27862 6316
rect 30742 6264 30748 6316
rect 30800 6304 30806 6316
rect 37553 6307 37611 6313
rect 37553 6304 37565 6307
rect 30800 6276 37565 6304
rect 30800 6264 30806 6276
rect 37553 6273 37565 6276
rect 37599 6304 37611 6307
rect 38013 6307 38071 6313
rect 38013 6304 38025 6307
rect 37599 6276 38025 6304
rect 37599 6273 37611 6276
rect 37553 6267 37611 6273
rect 38013 6273 38025 6276
rect 38059 6273 38071 6307
rect 38013 6267 38071 6273
rect 47578 6264 47584 6316
rect 47636 6304 47642 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 47636 6276 47961 6304
rect 47636 6264 47642 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 1596 6208 2329 6236
rect 2317 6205 2329 6208
rect 2363 6205 2375 6239
rect 11146 6236 11152 6248
rect 2317 6199 2375 6205
rect 2746 6208 11152 6236
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 2746 6168 2774 6208
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 14516 6208 18061 6236
rect 14516 6196 14522 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18322 6236 18328 6248
rect 18279 6208 18328 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 26970 6196 26976 6248
rect 27028 6236 27034 6248
rect 37734 6236 37740 6248
rect 27028 6208 37740 6236
rect 27028 6196 27034 6208
rect 37734 6196 37740 6208
rect 37792 6196 37798 6248
rect 1811 6140 2774 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 23934 6168 23940 6180
rect 4120 6140 23940 6168
rect 4120 6128 4126 6140
rect 23934 6128 23940 6140
rect 23992 6128 23998 6180
rect 25682 6128 25688 6180
rect 25740 6168 25746 6180
rect 36446 6168 36452 6180
rect 25740 6140 36452 6168
rect 25740 6128 25746 6140
rect 36446 6128 36452 6140
rect 36504 6128 36510 6180
rect 44177 6171 44235 6177
rect 44177 6137 44189 6171
rect 44223 6168 44235 6171
rect 47026 6168 47032 6180
rect 44223 6140 47032 6168
rect 44223 6137 44235 6140
rect 44177 6131 44235 6137
rect 47026 6128 47032 6140
rect 47084 6128 47090 6180
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19426 6100 19432 6112
rect 18739 6072 19432 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 37642 6060 37648 6112
rect 37700 6060 37706 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 2501 5899 2559 5905
rect 2501 5865 2513 5899
rect 2547 5896 2559 5899
rect 2590 5896 2596 5908
rect 2547 5868 2596 5896
rect 2547 5865 2559 5868
rect 2501 5859 2559 5865
rect 2590 5856 2596 5868
rect 2648 5856 2654 5908
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 47210 5896 47216 5908
rect 37700 5868 47216 5896
rect 37700 5856 37706 5868
rect 47210 5856 47216 5868
rect 47268 5856 47274 5908
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 1596 5732 3065 5760
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1596 5701 1624 5732
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 49145 5763 49203 5769
rect 49145 5729 49157 5763
rect 49191 5760 49203 5763
rect 49234 5760 49240 5772
rect 49191 5732 49240 5760
rect 49191 5729 49203 5732
rect 49145 5723 49203 5729
rect 49234 5720 49240 5732
rect 49292 5720 49298 5772
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2774 5692 2780 5704
rect 2363 5664 2780 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 39942 5652 39948 5704
rect 40000 5692 40006 5704
rect 43717 5695 43775 5701
rect 43717 5692 43729 5695
rect 40000 5664 43729 5692
rect 40000 5652 40006 5664
rect 43717 5661 43729 5664
rect 43763 5661 43775 5695
rect 43717 5655 43775 5661
rect 47670 5652 47676 5704
rect 47728 5692 47734 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 47728 5664 47961 5692
rect 47728 5652 47734 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 16298 5624 16304 5636
rect 1780 5596 16304 5624
rect 1780 5565 1808 5596
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 43901 5627 43959 5633
rect 43901 5593 43913 5627
rect 43947 5624 43959 5627
rect 45738 5624 45744 5636
rect 43947 5596 45744 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 45738 5584 45744 5596
rect 45796 5584 45802 5636
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5525 1823 5559
rect 1765 5519 1823 5525
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 37274 5312 37280 5364
rect 37332 5352 37338 5364
rect 37332 5324 37780 5352
rect 37332 5312 37338 5324
rect 37752 5293 37780 5324
rect 37737 5287 37795 5293
rect 37737 5253 37749 5287
rect 37783 5253 37795 5287
rect 37737 5247 37795 5253
rect 38470 5244 38476 5296
rect 38528 5284 38534 5296
rect 38933 5287 38991 5293
rect 38933 5284 38945 5287
rect 38528 5256 38945 5284
rect 38528 5244 38534 5256
rect 38933 5253 38945 5256
rect 38979 5253 38991 5287
rect 38933 5247 38991 5253
rect 49142 5244 49148 5296
rect 49200 5244 49206 5296
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 12802 5216 12808 5228
rect 2179 5188 12808 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 18874 5176 18880 5228
rect 18932 5176 18938 5228
rect 28350 5176 28356 5228
rect 28408 5216 28414 5228
rect 33318 5216 33324 5228
rect 28408 5188 33324 5216
rect 28408 5176 28414 5188
rect 33318 5176 33324 5188
rect 33376 5176 33382 5228
rect 45830 5176 45836 5228
rect 45888 5176 45894 5228
rect 47762 5176 47768 5228
rect 47820 5216 47826 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47820 5188 47961 5216
rect 47820 5176 47826 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 1360 5120 2421 5148
rect 1360 5108 1366 5120
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 19058 5108 19064 5160
rect 19116 5108 19122 5160
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48314 5148 48320 5160
rect 46891 5120 48320 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 38657 5083 38715 5089
rect 38657 5049 38669 5083
rect 38703 5080 38715 5083
rect 41322 5080 41328 5092
rect 38703 5052 41328 5080
rect 38703 5049 38715 5052
rect 38657 5043 38715 5049
rect 41322 5040 41328 5052
rect 41380 5040 41386 5092
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 15654 5012 15660 5024
rect 4488 4984 15660 5012
rect 4488 4972 4494 4984
rect 15654 4972 15660 4984
rect 15712 4972 15718 5024
rect 19521 5015 19579 5021
rect 19521 4981 19533 5015
rect 19567 5012 19579 5015
rect 20622 5012 20628 5024
rect 19567 4984 20628 5012
rect 19567 4981 19579 4984
rect 19521 4975 19579 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 37826 4972 37832 5024
rect 37884 4972 37890 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1360 4780 2145 4808
rect 1360 4768 1366 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 2133 4771 2191 4777
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 20714 4808 20720 4820
rect 6880 4780 20720 4808
rect 6880 4768 6886 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 36814 4768 36820 4820
rect 36872 4768 36878 4820
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 47118 4808 47124 4820
rect 37884 4780 47124 4808
rect 37884 4768 37890 4780
rect 47118 4768 47124 4780
rect 47176 4768 47182 4820
rect 1765 4743 1823 4749
rect 1765 4709 1777 4743
rect 1811 4740 1823 4743
rect 4062 4740 4068 4752
rect 1811 4712 4068 4740
rect 1811 4709 1823 4712
rect 1765 4703 1823 4709
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 22557 4743 22615 4749
rect 22557 4709 22569 4743
rect 22603 4740 22615 4743
rect 26142 4740 26148 4752
rect 22603 4712 26148 4740
rect 22603 4709 22615 4712
rect 22557 4703 22615 4709
rect 26142 4700 26148 4712
rect 26200 4700 26206 4752
rect 38930 4700 38936 4752
rect 38988 4740 38994 4752
rect 46477 4743 46535 4749
rect 46477 4740 46489 4743
rect 38988 4712 46489 4740
rect 38988 4700 38994 4712
rect 46477 4709 46489 4712
rect 46523 4709 46535 4743
rect 46477 4703 46535 4709
rect 19242 4632 19248 4684
rect 19300 4672 19306 4684
rect 20441 4675 20499 4681
rect 20441 4672 20453 4675
rect 19300 4644 20453 4672
rect 19300 4632 19306 4644
rect 20441 4641 20453 4644
rect 20487 4641 20499 4675
rect 20441 4635 20499 4641
rect 21726 4632 21732 4684
rect 21784 4672 21790 4684
rect 21913 4675 21971 4681
rect 21913 4672 21925 4675
rect 21784 4644 21925 4672
rect 21784 4632 21790 4644
rect 21913 4641 21925 4644
rect 21959 4641 21971 4675
rect 22922 4672 22928 4684
rect 21913 4635 21971 4641
rect 22020 4644 22928 4672
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4604 1639 4607
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 1627 4576 2329 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 19978 4564 19984 4616
rect 20036 4604 20042 4616
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 20036 4576 20637 4604
rect 20036 4564 20042 4576
rect 20625 4573 20637 4576
rect 20671 4604 20683 4607
rect 22020 4604 22048 4644
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23198 4632 23204 4684
rect 23256 4672 23262 4684
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 23256 4644 26801 4672
rect 23256 4632 23262 4644
rect 26789 4641 26801 4644
rect 26835 4641 26847 4675
rect 26789 4635 26847 4641
rect 36998 4632 37004 4684
rect 37056 4672 37062 4684
rect 47213 4675 47271 4681
rect 47213 4672 47225 4675
rect 37056 4644 47225 4672
rect 37056 4632 37062 4644
rect 47213 4641 47225 4644
rect 47259 4641 47271 4675
rect 47213 4635 47271 4641
rect 49145 4675 49203 4681
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49418 4672 49424 4684
rect 49191 4644 49424 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 20671 4576 22048 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 23084 4607 23142 4613
rect 23084 4604 23096 4607
rect 22388 4576 23096 4604
rect 19058 4496 19064 4548
rect 19116 4536 19122 4548
rect 22388 4536 22416 4576
rect 23084 4573 23096 4576
rect 23130 4604 23142 4607
rect 23566 4604 23572 4616
rect 23130 4576 23572 4604
rect 23130 4573 23142 4576
rect 23084 4567 23142 4573
rect 23566 4564 23572 4576
rect 23624 4564 23630 4616
rect 26973 4607 27031 4613
rect 26973 4573 26985 4607
rect 27019 4604 27031 4607
rect 32766 4604 32772 4616
rect 27019 4576 32772 4604
rect 27019 4573 27031 4576
rect 26973 4567 27031 4573
rect 32766 4564 32772 4576
rect 32824 4564 32830 4616
rect 36814 4564 36820 4616
rect 36872 4604 36878 4616
rect 37277 4607 37335 4613
rect 37277 4604 37289 4607
rect 36872 4576 37289 4604
rect 36872 4564 36878 4576
rect 37277 4573 37289 4576
rect 37323 4573 37335 4607
rect 37277 4567 37335 4573
rect 37734 4564 37740 4616
rect 37792 4604 37798 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 37792 4576 38025 4604
rect 37792 4564 37798 4576
rect 38013 4573 38025 4576
rect 38059 4604 38071 4607
rect 38473 4607 38531 4613
rect 38473 4604 38485 4607
rect 38059 4576 38485 4604
rect 38059 4573 38071 4576
rect 38013 4567 38071 4573
rect 38473 4573 38485 4576
rect 38519 4573 38531 4607
rect 38473 4567 38531 4573
rect 47302 4564 47308 4616
rect 47360 4604 47366 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 47360 4576 47961 4604
rect 47360 4564 47366 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 25133 4539 25191 4545
rect 25133 4536 25145 4539
rect 19116 4508 22416 4536
rect 22480 4508 25145 4536
rect 19116 4496 19122 4508
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21266 4468 21272 4480
rect 21131 4440 21272 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 21818 4468 21824 4480
rect 21416 4440 21824 4468
rect 21416 4428 21422 4440
rect 21818 4428 21824 4440
rect 21876 4468 21882 4480
rect 22480 4468 22508 4508
rect 25133 4505 25145 4508
rect 25179 4505 25191 4539
rect 25133 4499 25191 4505
rect 38197 4539 38255 4545
rect 38197 4505 38209 4539
rect 38243 4536 38255 4539
rect 39942 4536 39948 4548
rect 38243 4508 39948 4536
rect 38243 4505 38255 4508
rect 38197 4499 38255 4505
rect 39942 4496 39948 4508
rect 40000 4496 40006 4548
rect 46661 4539 46719 4545
rect 46661 4505 46673 4539
rect 46707 4505 46719 4539
rect 46661 4499 46719 4505
rect 47397 4539 47455 4545
rect 47397 4505 47409 4539
rect 47443 4536 47455 4539
rect 47670 4536 47676 4548
rect 47443 4508 47676 4536
rect 47443 4505 47455 4508
rect 47397 4499 47455 4505
rect 21876 4440 22508 4468
rect 23155 4471 23213 4477
rect 21876 4428 21882 4440
rect 23155 4437 23167 4471
rect 23201 4468 23213 4471
rect 25866 4468 25872 4480
rect 23201 4440 25872 4468
rect 23201 4437 23213 4440
rect 23155 4431 23213 4437
rect 25866 4428 25872 4440
rect 25924 4428 25930 4480
rect 37366 4428 37372 4480
rect 37424 4428 37430 4480
rect 46201 4471 46259 4477
rect 46201 4437 46213 4471
rect 46247 4468 46259 4471
rect 46676 4468 46704 4499
rect 47670 4496 47676 4508
rect 47728 4496 47734 4548
rect 49786 4468 49792 4480
rect 46247 4440 49792 4468
rect 46247 4437 46259 4440
rect 46201 4431 46259 4437
rect 49786 4428 49792 4440
rect 49844 4428 49850 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 4798 4264 4804 4276
rect 1820 4236 4804 4264
rect 1820 4224 1826 4236
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 13722 4224 13728 4276
rect 13780 4264 13786 4276
rect 21358 4264 21364 4276
rect 13780 4236 21364 4264
rect 13780 4224 13786 4236
rect 21358 4224 21364 4236
rect 21416 4224 21422 4276
rect 37366 4224 37372 4276
rect 37424 4264 37430 4276
rect 45646 4264 45652 4276
rect 37424 4236 45652 4264
rect 37424 4224 37430 4236
rect 45646 4224 45652 4236
rect 45704 4224 45710 4276
rect 1394 4156 1400 4208
rect 1452 4196 1458 4208
rect 1673 4199 1731 4205
rect 1673 4196 1685 4199
rect 1452 4168 1685 4196
rect 1452 4156 1458 4168
rect 1673 4165 1685 4168
rect 1719 4196 1731 4199
rect 1719 4168 2728 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 1360 4100 2329 4128
rect 1360 4088 1366 4100
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2700 4128 2728 4168
rect 22094 4156 22100 4208
rect 22152 4196 22158 4208
rect 22152 4168 23336 4196
rect 22152 4156 22158 4168
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2700 4100 3065 4128
rect 2317 4091 2375 4097
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 22348 4130 22406 4136
rect 22348 4096 22360 4130
rect 22394 4127 22406 4130
rect 22394 4099 22462 4127
rect 22394 4096 22406 4099
rect 2332 4060 2360 4091
rect 22348 4090 22406 4096
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2332 4032 2881 4060
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 4430 3992 4436 4004
rect 2547 3964 4436 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 4430 3952 4436 3964
rect 4488 3952 4494 4004
rect 16574 3952 16580 4004
rect 16632 3992 16638 4004
rect 18322 3992 18328 4004
rect 16632 3964 18328 3992
rect 16632 3952 16638 3964
rect 18322 3952 18328 3964
rect 18380 3992 18386 4004
rect 22434 3992 22462 4099
rect 22922 4088 22928 4140
rect 22980 4137 22986 4140
rect 22980 4131 23018 4137
rect 23006 4097 23018 4131
rect 22980 4091 23018 4097
rect 23063 4131 23121 4137
rect 23063 4097 23075 4131
rect 23109 4128 23121 4131
rect 23198 4128 23204 4140
rect 23109 4100 23204 4128
rect 23109 4097 23121 4100
rect 23063 4091 23121 4097
rect 22980 4088 23003 4091
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23308 4128 23336 4168
rect 25866 4156 25872 4208
rect 25924 4156 25930 4208
rect 23604 4131 23662 4137
rect 23604 4128 23616 4131
rect 23308 4100 23616 4128
rect 23604 4097 23616 4100
rect 23650 4097 23662 4131
rect 23604 4091 23662 4097
rect 26053 4131 26111 4137
rect 26053 4097 26065 4131
rect 26099 4128 26111 4131
rect 27614 4128 27620 4140
rect 26099 4100 27620 4128
rect 26099 4097 26111 4100
rect 26053 4091 26111 4097
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 45830 4088 45836 4140
rect 45888 4088 45894 4140
rect 46934 4088 46940 4140
rect 46992 4128 46998 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 46992 4100 47961 4128
rect 46992 4088 46998 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4128 49203 4131
rect 49326 4128 49332 4140
rect 49191 4100 49332 4128
rect 49191 4097 49203 4100
rect 49145 4091 49203 4097
rect 49326 4088 49332 4100
rect 49384 4088 49390 4140
rect 22975 4060 23003 4088
rect 23290 4060 23296 4072
rect 22975 4032 23296 4060
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 24854 4020 24860 4072
rect 24912 4020 24918 4072
rect 25774 4020 25780 4072
rect 25832 4060 25838 4072
rect 27157 4063 27215 4069
rect 27157 4060 27169 4063
rect 25832 4032 27169 4060
rect 25832 4020 25838 4032
rect 27157 4029 27169 4032
rect 27203 4029 27215 4063
rect 27157 4023 27215 4029
rect 28813 4063 28871 4069
rect 28813 4029 28825 4063
rect 28859 4029 28871 4063
rect 28813 4023 28871 4029
rect 28997 4063 29055 4069
rect 28997 4029 29009 4063
rect 29043 4060 29055 4063
rect 32858 4060 32864 4072
rect 29043 4032 32864 4060
rect 29043 4029 29055 4032
rect 28997 4023 29055 4029
rect 23707 3995 23765 4001
rect 18380 3964 23003 3992
rect 18380 3952 18386 3964
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 6822 3924 6828 3936
rect 1811 3896 6828 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 22419 3927 22477 3933
rect 22419 3893 22431 3927
rect 22465 3924 22477 3927
rect 22830 3924 22836 3936
rect 22465 3896 22836 3924
rect 22465 3893 22477 3896
rect 22419 3887 22477 3893
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 22975 3924 23003 3964
rect 23707 3961 23719 3995
rect 23753 3992 23765 3995
rect 28828 3992 28856 4023
rect 32858 4020 32864 4032
rect 32916 4020 32922 4072
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 23753 3964 28856 3992
rect 23753 3961 23765 3964
rect 23707 3955 23765 3961
rect 27522 3924 27528 3936
rect 22975 3896 27528 3924
rect 27522 3884 27528 3896
rect 27580 3884 27586 3936
rect 47670 3884 47676 3936
rect 47728 3884 47734 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 22002 3680 22008 3732
rect 22060 3720 22066 3732
rect 23017 3723 23075 3729
rect 23017 3720 23029 3723
rect 22060 3692 23029 3720
rect 22060 3680 22066 3692
rect 23017 3689 23029 3692
rect 23063 3689 23075 3723
rect 23017 3683 23075 3689
rect 23566 3680 23572 3732
rect 23624 3680 23630 3732
rect 23937 3723 23995 3729
rect 23937 3689 23949 3723
rect 23983 3720 23995 3723
rect 25958 3720 25964 3732
rect 23983 3692 25964 3720
rect 23983 3689 23995 3692
rect 23937 3683 23995 3689
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 41322 3680 41328 3732
rect 41380 3720 41386 3732
rect 41380 3692 46152 3720
rect 41380 3680 41386 3692
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 7524 3624 17264 3652
rect 7524 3612 7530 3624
rect 2133 3587 2191 3593
rect 2133 3553 2145 3587
rect 2179 3584 2191 3587
rect 2682 3584 2688 3596
rect 2179 3556 2688 3584
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 13722 3584 13728 3596
rect 3384 3556 13728 3584
rect 3384 3544 3390 3556
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 10318 3516 10324 3528
rect 9723 3488 10324 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 2424 3448 2452 3479
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 16574 3476 16580 3528
rect 16632 3476 16638 3528
rect 1360 3420 2452 3448
rect 1360 3408 1366 3420
rect 14090 3408 14096 3460
rect 14148 3448 14154 3460
rect 16393 3451 16451 3457
rect 16393 3448 16405 3451
rect 14148 3420 16405 3448
rect 14148 3408 14154 3420
rect 16393 3417 16405 3420
rect 16439 3417 16451 3451
rect 16393 3411 16451 3417
rect 10321 3383 10379 3389
rect 10321 3349 10333 3383
rect 10367 3380 10379 3383
rect 10686 3380 10692 3392
rect 10367 3352 10692 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 17236 3380 17264 3624
rect 33410 3612 33416 3664
rect 33468 3652 33474 3664
rect 45373 3655 45431 3661
rect 45373 3652 45385 3655
rect 33468 3624 45385 3652
rect 33468 3612 33474 3624
rect 45373 3621 45385 3624
rect 45419 3621 45431 3655
rect 45373 3615 45431 3621
rect 22830 3544 22836 3596
rect 22888 3584 22894 3596
rect 26237 3587 26295 3593
rect 26237 3584 26249 3587
rect 22888 3556 26249 3584
rect 22888 3544 22894 3556
rect 26237 3553 26249 3556
rect 26283 3553 26295 3587
rect 26237 3547 26295 3553
rect 36633 3587 36691 3593
rect 36633 3553 36645 3587
rect 36679 3584 36691 3587
rect 36679 3556 41920 3584
rect 36679 3553 36691 3556
rect 36633 3547 36691 3553
rect 20990 3476 20996 3528
rect 21048 3476 21054 3528
rect 23293 3519 23351 3525
rect 23293 3485 23305 3519
rect 23339 3516 23351 3519
rect 24026 3516 24032 3528
rect 23339 3488 24032 3516
rect 23339 3485 23351 3488
rect 23293 3479 23351 3485
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 24118 3476 24124 3528
rect 24176 3516 24182 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24176 3488 24593 3516
rect 24176 3476 24182 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 26421 3519 26479 3525
rect 26421 3485 26433 3519
rect 26467 3516 26479 3519
rect 28994 3516 29000 3528
rect 26467 3488 29000 3516
rect 26467 3485 26479 3488
rect 26421 3479 26479 3485
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 33318 3476 33324 3528
rect 33376 3516 33382 3528
rect 39206 3516 39212 3528
rect 33376 3488 39212 3516
rect 33376 3476 33382 3488
rect 39206 3476 39212 3488
rect 39264 3476 39270 3528
rect 41892 3516 41920 3556
rect 45830 3516 45836 3528
rect 41892 3488 45836 3516
rect 45830 3476 45836 3488
rect 45888 3476 45894 3528
rect 46124 3525 46152 3692
rect 49142 3544 49148 3596
rect 49200 3544 49206 3596
rect 46109 3519 46167 3525
rect 46109 3485 46121 3519
rect 46155 3485 46167 3519
rect 46109 3479 46167 3485
rect 47026 3476 47032 3528
rect 47084 3516 47090 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 47084 3488 47961 3516
rect 47084 3476 47090 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 21269 3451 21327 3457
rect 21269 3448 21281 3451
rect 19392 3420 21281 3448
rect 19392 3408 19398 3420
rect 21269 3417 21281 3420
rect 21315 3448 21327 3451
rect 21358 3448 21364 3460
rect 21315 3420 21364 3448
rect 21315 3417 21327 3420
rect 21269 3411 21327 3417
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 24136 3448 24164 3476
rect 22664 3420 24164 3448
rect 22664 3380 22692 3420
rect 36446 3408 36452 3460
rect 36504 3448 36510 3460
rect 36909 3451 36967 3457
rect 36909 3448 36921 3451
rect 36504 3420 36921 3448
rect 36504 3408 36510 3420
rect 36909 3417 36921 3420
rect 36955 3417 36967 3451
rect 36909 3411 36967 3417
rect 45097 3451 45155 3457
rect 45097 3417 45109 3451
rect 45143 3448 45155 3451
rect 45554 3448 45560 3460
rect 45143 3420 45560 3448
rect 45143 3417 45155 3420
rect 45097 3411 45155 3417
rect 45554 3408 45560 3420
rect 45612 3448 45618 3460
rect 47305 3451 47363 3457
rect 45612 3420 45657 3448
rect 45612 3408 45618 3420
rect 47305 3417 47317 3451
rect 47351 3448 47363 3451
rect 48682 3448 48688 3460
rect 47351 3420 48688 3448
rect 47351 3417 47363 3420
rect 47305 3411 47363 3417
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 17236 3352 22692 3380
rect 22738 3340 22744 3392
rect 22796 3340 22802 3392
rect 26326 3340 26332 3392
rect 26384 3380 26390 3392
rect 29638 3380 29644 3392
rect 26384 3352 29644 3380
rect 26384 3340 26390 3352
rect 29638 3340 29644 3352
rect 29696 3340 29702 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1360 3148 2145 3176
rect 1360 3136 1366 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 15194 3176 15200 3188
rect 14568 3148 15200 3176
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3040 1639 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1627 3012 2513 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3040 9459 3043
rect 9582 3040 9588 3052
rect 9447 3012 9588 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 9582 3000 9588 3012
rect 9640 3040 9646 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9640 3012 9689 3040
rect 9640 3000 9646 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 14568 3049 14596 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 19334 3176 19340 3188
rect 16347 3148 19340 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19981 3179 20039 3185
rect 19981 3176 19993 3179
rect 19536 3148 19993 3176
rect 16761 3111 16819 3117
rect 16761 3108 16773 3111
rect 16054 3080 16773 3108
rect 16761 3077 16773 3080
rect 16807 3108 16819 3111
rect 17862 3108 17868 3120
rect 16807 3080 17868 3108
rect 16807 3077 16819 3080
rect 16761 3071 16819 3077
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 9824 3012 12357 3040
rect 9824 3000 9830 3012
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3040 17647 3043
rect 19058 3040 19064 3052
rect 17635 3012 19064 3040
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19536 3049 19564 3148
rect 19981 3145 19993 3148
rect 20027 3145 20039 3179
rect 19981 3139 20039 3145
rect 21453 3179 21511 3185
rect 21453 3145 21465 3179
rect 21499 3176 21511 3179
rect 24578 3176 24584 3188
rect 21499 3148 24584 3176
rect 21499 3145 21511 3148
rect 21453 3139 21511 3145
rect 24578 3136 24584 3148
rect 24636 3136 24642 3188
rect 28353 3179 28411 3185
rect 28353 3176 28365 3179
rect 24688 3148 28365 3176
rect 22094 3108 22100 3120
rect 20180 3080 22100 3108
rect 20180 3049 20208 3080
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 24026 3108 24032 3120
rect 23768 3080 24032 3108
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 21266 3000 21272 3052
rect 21324 3000 21330 3052
rect 23768 3049 23796 3080
rect 24026 3068 24032 3080
rect 24084 3108 24090 3120
rect 24688 3108 24716 3148
rect 28353 3145 28365 3148
rect 28399 3176 28411 3179
rect 37734 3176 37740 3188
rect 28399 3148 37740 3176
rect 28399 3145 28411 3148
rect 28353 3139 28411 3145
rect 26326 3108 26332 3120
rect 24084 3080 24716 3108
rect 25714 3080 26332 3108
rect 24084 3068 24090 3080
rect 26326 3068 26332 3080
rect 26384 3068 26390 3120
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3040 22707 3043
rect 23017 3043 23075 3049
rect 23017 3040 23029 3043
rect 22695 3012 23029 3040
rect 22695 3009 22707 3012
rect 22649 3003 22707 3009
rect 23017 3009 23029 3012
rect 23063 3040 23075 3043
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23063 3012 23765 3040
rect 23063 3009 23075 3012
rect 23017 3003 23075 3009
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 26142 3000 26148 3052
rect 26200 3040 26206 3052
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 26200 3012 26433 3040
rect 26200 3000 26206 3012
rect 26421 3009 26433 3012
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 27985 3043 28043 3049
rect 27985 3009 27997 3043
rect 28031 3040 28043 3043
rect 28368 3040 28396 3139
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 29638 3068 29644 3120
rect 29696 3068 29702 3120
rect 49145 3111 49203 3117
rect 49145 3077 49157 3111
rect 49191 3108 49203 3111
rect 49234 3108 49240 3120
rect 49191 3080 49240 3108
rect 49191 3077 49203 3080
rect 49145 3071 49203 3077
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 28031 3012 28396 3040
rect 28031 3009 28043 3012
rect 27985 3003 28043 3009
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28868 3012 28917 3040
rect 28868 3000 28874 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 39942 3000 39948 3052
rect 40000 3040 40006 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 40000 3012 44005 3040
rect 40000 3000 40006 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 45833 3043 45891 3049
rect 45833 3040 45845 3043
rect 45796 3012 45845 3040
rect 45796 3000 45802 3012
rect 45833 3009 45845 3012
rect 45879 3009 45891 3043
rect 45833 3003 45891 3009
rect 47210 3000 47216 3052
rect 47268 3040 47274 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47268 3012 47961 3040
rect 47268 3000 47274 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 13035 2944 14841 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 21048 2944 24225 2972
rect 21048 2932 21054 2944
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24489 2975 24547 2981
rect 24489 2972 24501 2975
rect 24213 2935 24271 2941
rect 24320 2944 24501 2972
rect 1762 2864 1768 2916
rect 1820 2864 1826 2916
rect 20809 2907 20867 2913
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 22094 2904 22100 2916
rect 20855 2876 22100 2904
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 22186 2864 22192 2916
rect 22244 2864 22250 2916
rect 22738 2864 22744 2916
rect 22796 2904 22802 2916
rect 24320 2904 24348 2944
rect 24489 2941 24501 2944
rect 24535 2941 24547 2975
rect 24489 2935 24547 2941
rect 25958 2932 25964 2984
rect 26016 2972 26022 2984
rect 29181 2975 29239 2981
rect 29181 2972 29193 2975
rect 26016 2944 29193 2972
rect 26016 2932 26022 2944
rect 29181 2941 29193 2944
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 29638 2932 29644 2984
rect 29696 2972 29702 2984
rect 30650 2972 30656 2984
rect 29696 2944 30656 2972
rect 29696 2932 29702 2944
rect 30650 2932 30656 2944
rect 30708 2972 30714 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30708 2944 31033 2972
rect 30708 2932 30714 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 46750 2972 46756 2984
rect 45235 2944 46756 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 46842 2932 46848 2984
rect 46900 2932 46906 2984
rect 22796 2876 24348 2904
rect 22796 2864 22802 2876
rect 2314 2796 2320 2848
rect 2372 2796 2378 2848
rect 2774 2796 2780 2848
rect 2832 2796 2838 2848
rect 17402 2796 17408 2848
rect 17460 2796 17466 2848
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 22373 2839 22431 2845
rect 22373 2836 22385 2839
rect 21416 2808 22385 2836
rect 21416 2796 21422 2808
rect 22373 2805 22385 2808
rect 22419 2805 22431 2839
rect 22373 2799 22431 2805
rect 23290 2796 23296 2848
rect 23348 2796 23354 2848
rect 23492 2845 23520 2876
rect 27522 2864 27528 2916
rect 27580 2864 27586 2916
rect 38286 2904 38292 2916
rect 27908 2876 29040 2904
rect 23477 2839 23535 2845
rect 23477 2805 23489 2839
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 26605 2839 26663 2845
rect 26605 2805 26617 2839
rect 26651 2836 26663 2839
rect 27154 2836 27160 2848
rect 26651 2808 27160 2836
rect 26651 2805 26663 2808
rect 26605 2799 26663 2805
rect 27154 2796 27160 2808
rect 27212 2796 27218 2848
rect 27908 2845 27936 2876
rect 27893 2839 27951 2845
rect 27893 2805 27905 2839
rect 27939 2805 27951 2839
rect 29012 2836 29040 2876
rect 30668 2876 38292 2904
rect 30668 2845 30696 2876
rect 38286 2864 38292 2876
rect 38344 2864 38350 2916
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 29012 2808 30665 2836
rect 27893 2799 27951 2805
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 2547 2604 16574 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 1765 2567 1823 2573
rect 1765 2533 1777 2567
rect 1811 2533 1823 2567
rect 1765 2527 1823 2533
rect 3237 2567 3295 2573
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 9585 2567 9643 2573
rect 3283 2536 6914 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 1780 2496 1808 2527
rect 6886 2496 6914 2536
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 9766 2564 9772 2576
rect 9631 2536 9772 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 16546 2564 16574 2604
rect 24026 2592 24032 2644
rect 24084 2592 24090 2644
rect 26326 2592 26332 2644
rect 26384 2592 26390 2644
rect 27614 2592 27620 2644
rect 27672 2592 27678 2644
rect 28994 2592 29000 2644
rect 29052 2592 29058 2644
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 32916 2604 35081 2632
rect 32916 2592 32922 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 22462 2564 22468 2576
rect 16546 2536 22468 2564
rect 22462 2524 22468 2536
rect 22520 2524 22526 2576
rect 27632 2564 27660 2592
rect 30837 2567 30895 2573
rect 30837 2564 30849 2567
rect 27632 2536 30849 2564
rect 30837 2533 30849 2536
rect 30883 2533 30895 2567
rect 30837 2527 30895 2533
rect 32766 2524 32772 2576
rect 32824 2564 32830 2576
rect 32953 2567 33011 2573
rect 32953 2564 32965 2567
rect 32824 2536 32965 2564
rect 32824 2524 32830 2536
rect 32953 2533 32965 2536
rect 32999 2533 33011 2567
rect 32953 2527 33011 2533
rect 34330 2524 34336 2576
rect 34388 2564 34394 2576
rect 34388 2536 43852 2564
rect 34388 2524 34394 2536
rect 12250 2496 12256 2508
rect 1780 2468 4384 2496
rect 6886 2468 12256 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2428 1639 2431
rect 2774 2428 2780 2440
rect 1627 2400 2780 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2884 2400 3065 2428
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2314 2360 2320 2372
rect 1268 2332 2320 2360
rect 1268 2320 1274 2332
rect 2314 2320 2320 2332
rect 2372 2360 2378 2372
rect 2409 2363 2467 2369
rect 2409 2360 2421 2363
rect 2372 2332 2421 2360
rect 2372 2320 2378 2332
rect 2409 2329 2421 2332
rect 2455 2329 2467 2363
rect 2409 2323 2467 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 2884 2292 2912 2400
rect 3053 2397 3065 2400
rect 3099 2428 3111 2431
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3099 2400 3525 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 4356 2360 4384 2468
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 19978 2496 19984 2508
rect 19306 2468 19984 2496
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2428 9459 2431
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 9447 2400 10057 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 10686 2388 10692 2440
rect 10744 2388 10750 2440
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 14090 2428 14096 2440
rect 13219 2400 14096 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 17402 2428 17408 2440
rect 15703 2400 17408 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18877 2431 18935 2437
rect 18279 2400 18736 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 4356 2332 6914 2360
rect 1360 2264 2912 2292
rect 6886 2292 6914 2332
rect 11698 2320 11704 2372
rect 11756 2360 11762 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11756 2332 11989 2360
rect 11756 2320 11762 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 13872 2332 14473 2360
rect 13872 2320 13878 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 14461 2323 14519 2329
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 17037 2363 17095 2369
rect 17037 2360 17049 2363
rect 15988 2332 17049 2360
rect 15988 2320 15994 2332
rect 17037 2329 17049 2332
rect 17083 2329 17095 2363
rect 17037 2323 17095 2329
rect 14734 2292 14740 2304
rect 6886 2264 14740 2292
rect 1360 2252 1366 2264
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 18708 2301 18736 2400
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19306 2428 19334 2468
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22336 2468 22845 2496
rect 22336 2456 22342 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 24394 2456 24400 2508
rect 24452 2496 24458 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24452 2468 25053 2496
rect 24452 2456 24458 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 37734 2456 37740 2508
rect 37792 2456 37798 2508
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 43824 2505 43852 2536
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 41380 2468 41429 2496
rect 41380 2456 41386 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 41417 2459 41475 2465
rect 43809 2499 43867 2505
rect 43809 2465 43821 2499
rect 43855 2465 43867 2499
rect 43809 2459 43867 2465
rect 49142 2456 49148 2508
rect 49200 2456 49206 2508
rect 18923 2400 19334 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 19628 2400 20085 2428
rect 19628 2301 19656 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22152 2400 22385 2428
rect 22152 2388 22158 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29181 2431 29239 2437
rect 29181 2428 29193 2431
rect 29052 2400 29193 2428
rect 29052 2388 29058 2400
rect 29181 2397 29193 2400
rect 29227 2428 29239 2431
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29227 2400 29561 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 33192 2400 33425 2428
rect 33192 2388 33198 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35032 2400 35265 2428
rect 35032 2388 35038 2400
rect 35253 2397 35265 2400
rect 35299 2428 35311 2431
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35299 2400 35541 2428
rect 35299 2397 35311 2400
rect 35253 2391 35311 2397
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35529 2391 35587 2397
rect 37108 2400 37473 2428
rect 37108 2304 37136 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38286 2388 38292 2440
rect 38344 2428 38350 2440
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 38344 2400 40693 2428
rect 38344 2388 38350 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 40681 2391 40739 2397
rect 43456 2400 43545 2428
rect 43456 2304 43484 2400
rect 43533 2397 43545 2400
rect 43579 2397 43591 2431
rect 43533 2391 43591 2397
rect 45646 2388 45652 2440
rect 45704 2428 45710 2440
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 45704 2400 45845 2428
rect 45704 2388 45710 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 47176 2400 47961 2428
rect 47176 2388 47182 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2360 47087 2363
rect 48498 2360 48504 2372
rect 47075 2332 48504 2360
rect 47075 2329 47087 2332
rect 47029 2323 47087 2329
rect 48498 2320 48504 2332
rect 48556 2320 48562 2372
rect 18693 2295 18751 2301
rect 18693 2261 18705 2295
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 37090 2252 37096 2304
rect 37148 2252 37154 2304
rect 43257 2295 43315 2301
rect 43257 2261 43269 2295
rect 43303 2292 43315 2295
rect 43438 2292 43444 2304
rect 43303 2264 43444 2292
rect 43303 2261 43315 2264
rect 43257 2255 43315 2261
rect 43438 2252 43444 2264
rect 43496 2252 43502 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 3148 25440 3200 25492
rect 9772 25440 9824 25492
rect 39580 24964 39632 25016
rect 45744 24964 45796 25016
rect 21548 24896 21600 24948
rect 25964 24896 26016 24948
rect 26056 24896 26108 24948
rect 40960 24896 41012 24948
rect 25872 24828 25924 24880
rect 40408 24828 40460 24880
rect 3884 24760 3936 24812
rect 5908 24760 5960 24812
rect 16028 24760 16080 24812
rect 21732 24760 21784 24812
rect 29920 24760 29972 24812
rect 32864 24760 32916 24812
rect 34888 24760 34940 24812
rect 44364 24760 44416 24812
rect 18880 24692 18932 24744
rect 27252 24692 27304 24744
rect 29552 24692 29604 24744
rect 30656 24692 30708 24744
rect 33968 24692 34020 24744
rect 35164 24692 35216 24744
rect 40592 24692 40644 24744
rect 16212 24624 16264 24676
rect 24032 24624 24084 24676
rect 26424 24624 26476 24676
rect 34980 24624 35032 24676
rect 37556 24624 37608 24676
rect 37648 24624 37700 24676
rect 41052 24624 41104 24676
rect 46296 24624 46348 24676
rect 47768 24624 47820 24676
rect 17868 24556 17920 24608
rect 21640 24556 21692 24608
rect 21732 24556 21784 24608
rect 24492 24556 24544 24608
rect 24768 24556 24820 24608
rect 30380 24556 30432 24608
rect 30656 24556 30708 24608
rect 31024 24556 31076 24608
rect 32496 24556 32548 24608
rect 33140 24556 33192 24608
rect 39856 24556 39908 24608
rect 40040 24556 40092 24608
rect 44548 24556 44600 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 3516 24216 3568 24268
rect 3884 24148 3936 24200
rect 10048 24352 10100 24404
rect 6736 24216 6788 24268
rect 8668 24216 8720 24268
rect 4620 24191 4672 24200
rect 4620 24157 4629 24191
rect 4629 24157 4663 24191
rect 4663 24157 4672 24191
rect 4620 24148 4672 24157
rect 7104 24148 7156 24200
rect 7472 24148 7524 24200
rect 15568 24284 15620 24336
rect 11796 24216 11848 24268
rect 13820 24216 13872 24268
rect 17684 24216 17736 24268
rect 9496 24080 9548 24132
rect 12624 24080 12676 24132
rect 14280 24148 14332 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 20720 24352 20772 24404
rect 22560 24352 22612 24404
rect 26332 24352 26384 24404
rect 26424 24395 26476 24404
rect 26424 24361 26433 24395
rect 26433 24361 26467 24395
rect 26467 24361 26476 24395
rect 26424 24352 26476 24361
rect 27252 24395 27304 24404
rect 27252 24361 27261 24395
rect 27261 24361 27295 24395
rect 27295 24361 27304 24395
rect 27252 24352 27304 24361
rect 19524 24216 19576 24268
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 20996 24216 21048 24268
rect 22192 24216 22244 24268
rect 22468 24259 22520 24268
rect 22468 24225 22477 24259
rect 22477 24225 22511 24259
rect 22511 24225 22520 24259
rect 22468 24216 22520 24225
rect 14924 24080 14976 24132
rect 18696 24080 18748 24132
rect 21456 24148 21508 24200
rect 6644 24012 6696 24064
rect 7472 24012 7524 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 11152 24012 11204 24064
rect 11796 24012 11848 24064
rect 18604 24012 18656 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 22652 24080 22704 24132
rect 25780 24327 25832 24336
rect 25780 24293 25789 24327
rect 25789 24293 25823 24327
rect 25823 24293 25832 24327
rect 25780 24284 25832 24293
rect 33048 24352 33100 24404
rect 28632 24284 28684 24336
rect 25228 24148 25280 24200
rect 26424 24216 26476 24268
rect 27344 24216 27396 24268
rect 26240 24148 26292 24200
rect 31576 24284 31628 24336
rect 34612 24352 34664 24404
rect 39488 24352 39540 24404
rect 41052 24395 41104 24404
rect 41052 24361 41061 24395
rect 41061 24361 41095 24395
rect 41095 24361 41104 24395
rect 41052 24352 41104 24361
rect 42524 24352 42576 24404
rect 36452 24284 36504 24336
rect 24492 24080 24544 24132
rect 24400 24012 24452 24064
rect 25320 24080 25372 24132
rect 26608 24123 26660 24132
rect 26608 24089 26617 24123
rect 26617 24089 26651 24123
rect 26651 24089 26660 24123
rect 26608 24080 26660 24089
rect 27252 24080 27304 24132
rect 27344 24123 27396 24132
rect 27344 24089 27353 24123
rect 27353 24089 27387 24123
rect 27387 24089 27396 24123
rect 27344 24080 27396 24089
rect 29920 24191 29972 24200
rect 29920 24157 29929 24191
rect 29929 24157 29963 24191
rect 29963 24157 29972 24191
rect 29920 24148 29972 24157
rect 30380 24191 30432 24200
rect 30380 24157 30389 24191
rect 30389 24157 30423 24191
rect 30423 24157 30432 24191
rect 30380 24148 30432 24157
rect 26976 24012 27028 24064
rect 27804 24012 27856 24064
rect 28540 24012 28592 24064
rect 28632 24012 28684 24064
rect 30564 24055 30616 24064
rect 30564 24021 30573 24055
rect 30573 24021 30607 24055
rect 30607 24021 30616 24055
rect 30564 24012 30616 24021
rect 34244 24259 34296 24268
rect 34244 24225 34253 24259
rect 34253 24225 34287 24259
rect 34287 24225 34296 24259
rect 34244 24216 34296 24225
rect 35164 24216 35216 24268
rect 37188 24216 37240 24268
rect 37372 24216 37424 24268
rect 39672 24284 39724 24336
rect 40316 24216 40368 24268
rect 40592 24259 40644 24268
rect 40592 24225 40601 24259
rect 40601 24225 40635 24259
rect 40635 24225 40644 24259
rect 40592 24216 40644 24225
rect 32496 24191 32548 24200
rect 32496 24157 32505 24191
rect 32505 24157 32539 24191
rect 32539 24157 32548 24191
rect 32496 24148 32548 24157
rect 32864 24148 32916 24200
rect 33876 24148 33928 24200
rect 35532 24080 35584 24132
rect 36820 24080 36872 24132
rect 37648 24080 37700 24132
rect 38844 24191 38896 24200
rect 38844 24157 38853 24191
rect 38853 24157 38887 24191
rect 38887 24157 38896 24191
rect 38844 24148 38896 24157
rect 39396 24148 39448 24200
rect 42800 24148 42852 24200
rect 43352 24148 43404 24200
rect 40132 24080 40184 24132
rect 31852 24055 31904 24064
rect 31852 24021 31861 24055
rect 31861 24021 31895 24055
rect 31895 24021 31904 24055
rect 31852 24012 31904 24021
rect 32036 24012 32088 24064
rect 32956 24055 33008 24064
rect 32956 24021 32965 24055
rect 32965 24021 32999 24055
rect 32999 24021 33008 24055
rect 32956 24012 33008 24021
rect 33600 24055 33652 24064
rect 33600 24021 33609 24055
rect 33609 24021 33643 24055
rect 33643 24021 33652 24055
rect 33600 24012 33652 24021
rect 34980 24012 35032 24064
rect 35440 24012 35492 24064
rect 35624 24055 35676 24064
rect 35624 24021 35633 24055
rect 35633 24021 35667 24055
rect 35667 24021 35676 24055
rect 35624 24012 35676 24021
rect 36084 24055 36136 24064
rect 36084 24021 36093 24055
rect 36093 24021 36127 24055
rect 36127 24021 36136 24055
rect 36084 24012 36136 24021
rect 37556 24012 37608 24064
rect 38568 24012 38620 24064
rect 38752 24012 38804 24064
rect 39304 24055 39356 24064
rect 39304 24021 39313 24055
rect 39313 24021 39347 24055
rect 39347 24021 39356 24055
rect 39304 24012 39356 24021
rect 40040 24055 40092 24064
rect 40040 24021 40049 24055
rect 40049 24021 40083 24055
rect 40083 24021 40092 24055
rect 40040 24012 40092 24021
rect 40776 24012 40828 24064
rect 41236 24080 41288 24132
rect 44548 24191 44600 24200
rect 44548 24157 44557 24191
rect 44557 24157 44591 24191
rect 44591 24157 44600 24191
rect 44548 24148 44600 24157
rect 46480 24284 46532 24336
rect 47124 24080 47176 24132
rect 47768 24080 47820 24132
rect 49056 24148 49108 24200
rect 43628 24012 43680 24064
rect 43720 24055 43772 24064
rect 43720 24021 43729 24055
rect 43729 24021 43763 24055
rect 43763 24021 43772 24055
rect 43720 24012 43772 24021
rect 44364 24055 44416 24064
rect 44364 24021 44373 24055
rect 44373 24021 44407 24055
rect 44407 24021 44416 24055
rect 44364 24012 44416 24021
rect 46020 24012 46072 24064
rect 46572 24055 46624 24064
rect 46572 24021 46581 24055
rect 46581 24021 46615 24055
rect 46615 24021 46624 24055
rect 46572 24012 46624 24021
rect 49148 24055 49200 24064
rect 49148 24021 49157 24055
rect 49157 24021 49191 24055
rect 49191 24021 49200 24055
rect 49148 24012 49200 24021
rect 49332 24012 49384 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 4620 23808 4672 23860
rect 10324 23808 10376 23860
rect 4068 23715 4120 23724
rect 4068 23681 4077 23715
rect 4077 23681 4111 23715
rect 4111 23681 4120 23715
rect 4068 23672 4120 23681
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 4712 23672 4764 23681
rect 4160 23604 4212 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 8300 23672 8352 23724
rect 11796 23740 11848 23792
rect 16212 23808 16264 23860
rect 8392 23604 8444 23656
rect 9220 23604 9272 23656
rect 10600 23647 10652 23656
rect 10600 23613 10609 23647
rect 10609 23613 10643 23647
rect 10643 23613 10652 23647
rect 10600 23604 10652 23613
rect 12716 23672 12768 23724
rect 14188 23740 14240 23792
rect 14372 23740 14424 23792
rect 19616 23808 19668 23860
rect 21548 23808 21600 23860
rect 21640 23808 21692 23860
rect 18880 23740 18932 23792
rect 20352 23740 20404 23792
rect 24308 23740 24360 23792
rect 25780 23740 25832 23792
rect 27620 23740 27672 23792
rect 3976 23536 4028 23588
rect 5816 23536 5868 23588
rect 16396 23604 16448 23656
rect 18328 23604 18380 23656
rect 2780 23468 2832 23520
rect 5724 23468 5776 23520
rect 6000 23468 6052 23520
rect 18788 23511 18840 23520
rect 18788 23477 18797 23511
rect 18797 23477 18831 23511
rect 18831 23477 18840 23511
rect 18788 23468 18840 23477
rect 21548 23672 21600 23724
rect 22100 23604 22152 23656
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 25044 23672 25096 23724
rect 22744 23536 22796 23588
rect 21088 23468 21140 23520
rect 21456 23511 21508 23520
rect 21456 23477 21465 23511
rect 21465 23477 21499 23511
rect 21499 23477 21508 23511
rect 21456 23468 21508 23477
rect 24216 23604 24268 23656
rect 23480 23468 23532 23520
rect 26608 23647 26660 23656
rect 26608 23613 26617 23647
rect 26617 23613 26651 23647
rect 26651 23613 26660 23647
rect 26608 23604 26660 23613
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 40040 23808 40092 23860
rect 41052 23808 41104 23860
rect 46756 23808 46808 23860
rect 47124 23851 47176 23860
rect 47124 23817 47133 23851
rect 47133 23817 47167 23851
rect 47167 23817 47176 23851
rect 47124 23808 47176 23817
rect 47308 23808 47360 23860
rect 48596 23808 48648 23860
rect 49332 23851 49384 23860
rect 49332 23817 49341 23851
rect 49341 23817 49375 23851
rect 49375 23817 49384 23851
rect 49332 23808 49384 23817
rect 32588 23740 32640 23792
rect 33048 23740 33100 23792
rect 35624 23740 35676 23792
rect 38844 23740 38896 23792
rect 39764 23740 39816 23792
rect 39856 23740 39908 23792
rect 28356 23604 28408 23656
rect 30380 23672 30432 23724
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 29184 23604 29236 23656
rect 29736 23536 29788 23588
rect 30196 23536 30248 23588
rect 31760 23647 31812 23656
rect 31760 23613 31769 23647
rect 31769 23613 31803 23647
rect 31803 23613 31812 23647
rect 31760 23604 31812 23613
rect 31852 23604 31904 23656
rect 34060 23672 34112 23724
rect 35440 23672 35492 23724
rect 34520 23604 34572 23656
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 24860 23511 24912 23520
rect 24860 23477 24869 23511
rect 24869 23477 24903 23511
rect 24903 23477 24912 23511
rect 24860 23468 24912 23477
rect 28356 23468 28408 23520
rect 29368 23468 29420 23520
rect 30288 23468 30340 23520
rect 32036 23536 32088 23588
rect 35348 23647 35400 23656
rect 35348 23613 35357 23647
rect 35357 23613 35391 23647
rect 35391 23613 35400 23647
rect 35348 23604 35400 23613
rect 35624 23604 35676 23656
rect 35992 23604 36044 23656
rect 36452 23647 36504 23656
rect 36452 23613 36461 23647
rect 36461 23613 36495 23647
rect 36495 23613 36504 23647
rect 36452 23604 36504 23613
rect 35440 23536 35492 23588
rect 39580 23672 39632 23724
rect 45560 23740 45612 23792
rect 43996 23672 44048 23724
rect 45928 23715 45980 23724
rect 45928 23681 45937 23715
rect 45937 23681 45971 23715
rect 45971 23681 45980 23715
rect 45928 23672 45980 23681
rect 47768 23740 47820 23792
rect 39212 23536 39264 23588
rect 39764 23604 39816 23656
rect 36268 23468 36320 23520
rect 38568 23511 38620 23520
rect 38568 23477 38577 23511
rect 38577 23477 38611 23511
rect 38611 23477 38620 23511
rect 38568 23468 38620 23477
rect 39120 23468 39172 23520
rect 39488 23536 39540 23588
rect 40684 23647 40736 23656
rect 40684 23613 40693 23647
rect 40693 23613 40727 23647
rect 40727 23613 40736 23647
rect 40684 23604 40736 23613
rect 40960 23647 41012 23656
rect 40960 23613 40969 23647
rect 40969 23613 41003 23647
rect 41003 23613 41012 23647
rect 40960 23604 41012 23613
rect 42800 23604 42852 23656
rect 44548 23604 44600 23656
rect 48780 23715 48832 23724
rect 48780 23681 48789 23715
rect 48789 23681 48823 23715
rect 48823 23681 48832 23715
rect 48780 23672 48832 23681
rect 42064 23536 42116 23588
rect 47400 23536 47452 23588
rect 39396 23468 39448 23520
rect 42432 23511 42484 23520
rect 42432 23477 42441 23511
rect 42441 23477 42475 23511
rect 42475 23477 42484 23511
rect 42432 23468 42484 23477
rect 43536 23468 43588 23520
rect 46112 23468 46164 23520
rect 47676 23468 47728 23520
rect 47952 23468 48004 23520
rect 49056 23468 49108 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 4712 23307 4764 23316
rect 4712 23273 4721 23307
rect 4721 23273 4755 23307
rect 4755 23273 4764 23307
rect 4712 23264 4764 23273
rect 5632 23264 5684 23316
rect 14188 23307 14240 23316
rect 14188 23273 14197 23307
rect 14197 23273 14231 23307
rect 14231 23273 14240 23307
rect 14188 23264 14240 23273
rect 4436 23060 4488 23112
rect 9220 23196 9272 23248
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 15660 23196 15712 23248
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 13360 23128 13412 23180
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 1768 23035 1820 23044
rect 1768 23001 1777 23035
rect 1777 23001 1811 23035
rect 1811 23001 1820 23035
rect 1768 22992 1820 23001
rect 3608 22992 3660 23044
rect 6644 23060 6696 23112
rect 9128 23060 9180 23112
rect 11888 23103 11940 23112
rect 11888 23069 11897 23103
rect 11897 23069 11931 23103
rect 11931 23069 11940 23103
rect 11888 23060 11940 23069
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 19064 23128 19116 23180
rect 20260 23264 20312 23316
rect 22468 23264 22520 23316
rect 23388 23264 23440 23316
rect 24216 23264 24268 23316
rect 19616 23239 19668 23248
rect 19616 23205 19625 23239
rect 19625 23205 19659 23239
rect 19659 23205 19668 23239
rect 19616 23196 19668 23205
rect 22744 23196 22796 23248
rect 17500 23060 17552 23112
rect 19340 23060 19392 23112
rect 4620 22924 4672 22976
rect 5356 22924 5408 22976
rect 14096 22924 14148 22976
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 17132 22967 17184 22976
rect 17132 22933 17141 22967
rect 17141 22933 17175 22967
rect 17175 22933 17184 22967
rect 17132 22924 17184 22933
rect 18696 22992 18748 23044
rect 19800 23035 19852 23044
rect 19800 23001 19809 23035
rect 19809 23001 19843 23035
rect 19843 23001 19852 23035
rect 19800 22992 19852 23001
rect 17776 22924 17828 22976
rect 18880 22924 18932 22976
rect 20352 22967 20404 22976
rect 20352 22933 20361 22967
rect 20361 22933 20395 22967
rect 20395 22933 20404 22967
rect 20352 22924 20404 22933
rect 21180 23128 21232 23180
rect 22192 23128 22244 23180
rect 24860 23264 24912 23316
rect 25044 23264 25096 23316
rect 29736 23307 29788 23316
rect 29736 23273 29745 23307
rect 29745 23273 29779 23307
rect 29779 23273 29788 23307
rect 29736 23264 29788 23273
rect 30840 23264 30892 23316
rect 33232 23264 33284 23316
rect 33876 23264 33928 23316
rect 34244 23264 34296 23316
rect 25228 23239 25280 23248
rect 25228 23205 25237 23239
rect 25237 23205 25271 23239
rect 25271 23205 25280 23239
rect 25228 23196 25280 23205
rect 27804 23196 27856 23248
rect 24860 23128 24912 23180
rect 26700 23128 26752 23180
rect 29276 23128 29328 23180
rect 22100 23103 22152 23112
rect 22100 23069 22109 23103
rect 22109 23069 22143 23103
rect 22143 23069 22152 23103
rect 22100 23060 22152 23069
rect 23756 23103 23808 23112
rect 23756 23069 23765 23103
rect 23765 23069 23799 23103
rect 23799 23069 23808 23103
rect 23756 23060 23808 23069
rect 24768 23103 24820 23112
rect 24768 23069 24777 23103
rect 24777 23069 24811 23103
rect 24811 23069 24820 23103
rect 24768 23060 24820 23069
rect 25688 23103 25740 23112
rect 25688 23069 25697 23103
rect 25697 23069 25731 23103
rect 25731 23069 25740 23103
rect 25688 23060 25740 23069
rect 31300 23196 31352 23248
rect 33968 23196 34020 23248
rect 34060 23196 34112 23248
rect 30196 23171 30248 23180
rect 30196 23137 30205 23171
rect 30205 23137 30239 23171
rect 30239 23137 30248 23171
rect 30196 23128 30248 23137
rect 30288 23171 30340 23180
rect 30288 23137 30297 23171
rect 30297 23137 30331 23171
rect 30331 23137 30340 23171
rect 30288 23128 30340 23137
rect 31024 23171 31076 23180
rect 31024 23137 31033 23171
rect 31033 23137 31067 23171
rect 31067 23137 31076 23171
rect 31024 23128 31076 23137
rect 29460 23060 29512 23112
rect 21088 22992 21140 23044
rect 21916 22992 21968 23044
rect 25136 22992 25188 23044
rect 22836 22924 22888 22976
rect 23296 22967 23348 22976
rect 23296 22933 23305 22967
rect 23305 22933 23339 22967
rect 23339 22933 23348 22967
rect 23296 22924 23348 22933
rect 26240 22992 26292 23044
rect 27252 22992 27304 23044
rect 25320 22967 25372 22976
rect 25320 22933 25329 22967
rect 25329 22933 25363 22967
rect 25363 22933 25372 22967
rect 25320 22924 25372 22933
rect 26332 22924 26384 22976
rect 29920 22992 29972 23044
rect 30012 22924 30064 22976
rect 30104 22967 30156 22976
rect 30104 22933 30113 22967
rect 30113 22933 30147 22967
rect 30147 22933 30156 22967
rect 30104 22924 30156 22933
rect 31760 23128 31812 23180
rect 34336 23128 34388 23180
rect 35348 23128 35400 23180
rect 37464 23264 37516 23316
rect 39028 23264 39080 23316
rect 39948 23264 40000 23316
rect 38292 23128 38344 23180
rect 38660 23128 38712 23180
rect 39488 23171 39540 23180
rect 39488 23137 39497 23171
rect 39497 23137 39531 23171
rect 39531 23137 39540 23171
rect 39488 23128 39540 23137
rect 40684 23171 40736 23180
rect 40684 23137 40693 23171
rect 40693 23137 40727 23171
rect 40727 23137 40736 23171
rect 40684 23128 40736 23137
rect 43996 23307 44048 23316
rect 43996 23273 44005 23307
rect 44005 23273 44039 23307
rect 44039 23273 44048 23307
rect 43996 23264 44048 23273
rect 48780 23264 48832 23316
rect 49240 23307 49292 23316
rect 49240 23273 49249 23307
rect 49249 23273 49283 23307
rect 49283 23273 49292 23307
rect 49240 23264 49292 23273
rect 46756 23239 46808 23248
rect 46756 23205 46765 23239
rect 46765 23205 46799 23239
rect 46799 23205 46808 23239
rect 46756 23196 46808 23205
rect 42800 23128 42852 23180
rect 43996 23128 44048 23180
rect 46572 23128 46624 23180
rect 31392 23103 31444 23112
rect 31392 23069 31401 23103
rect 31401 23069 31435 23103
rect 31435 23069 31444 23103
rect 31392 23060 31444 23069
rect 31760 22992 31812 23044
rect 30380 22924 30432 22976
rect 31208 22924 31260 22976
rect 34520 22992 34572 23044
rect 33784 22924 33836 22976
rect 34060 22924 34112 22976
rect 36268 22924 36320 22976
rect 37648 23060 37700 23112
rect 39948 23060 40000 23112
rect 40040 23060 40092 23112
rect 38660 22992 38712 23044
rect 39120 22992 39172 23044
rect 41328 23060 41380 23112
rect 46480 23060 46532 23112
rect 46664 23060 46716 23112
rect 47676 23060 47728 23112
rect 36636 22924 36688 22976
rect 37832 22924 37884 22976
rect 39948 22924 40000 22976
rect 40132 22924 40184 22976
rect 40500 22967 40552 22976
rect 40500 22933 40509 22967
rect 40509 22933 40543 22967
rect 40543 22933 40552 22967
rect 40500 22924 40552 22933
rect 40868 22924 40920 22976
rect 42708 22992 42760 23044
rect 43536 22992 43588 23044
rect 44732 22992 44784 23044
rect 45376 23035 45428 23044
rect 45376 23001 45385 23035
rect 45385 23001 45419 23035
rect 45419 23001 45428 23035
rect 45376 22992 45428 23001
rect 46020 23035 46072 23044
rect 46020 23001 46029 23035
rect 46029 23001 46063 23035
rect 46063 23001 46072 23035
rect 46020 22992 46072 23001
rect 47308 22992 47360 23044
rect 48596 22992 48648 23044
rect 43720 22924 43772 22976
rect 46940 22924 46992 22976
rect 47676 22924 47728 22976
rect 47952 22924 48004 22976
rect 49332 22924 49384 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 1584 22720 1636 22772
rect 3424 22720 3476 22772
rect 4804 22695 4856 22704
rect 4804 22661 4813 22695
rect 4813 22661 4847 22695
rect 4847 22661 4856 22695
rect 4804 22652 4856 22661
rect 7104 22695 7156 22704
rect 7104 22661 7113 22695
rect 7113 22661 7147 22695
rect 7147 22661 7156 22695
rect 7104 22652 7156 22661
rect 9956 22695 10008 22704
rect 9956 22661 9965 22695
rect 9965 22661 9999 22695
rect 9999 22661 10008 22695
rect 9956 22652 10008 22661
rect 12808 22695 12860 22704
rect 12808 22661 12817 22695
rect 12817 22661 12851 22695
rect 12851 22661 12860 22695
rect 12808 22652 12860 22661
rect 18696 22720 18748 22772
rect 19340 22720 19392 22772
rect 21180 22763 21232 22772
rect 21180 22729 21189 22763
rect 21189 22729 21223 22763
rect 21223 22729 21232 22763
rect 21180 22720 21232 22729
rect 22192 22720 22244 22772
rect 25044 22720 25096 22772
rect 26240 22720 26292 22772
rect 15016 22652 15068 22704
rect 15108 22695 15160 22704
rect 15108 22661 15117 22695
rect 15117 22661 15151 22695
rect 15151 22661 15160 22695
rect 15108 22652 15160 22661
rect 17592 22652 17644 22704
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 7196 22584 7248 22636
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 11152 22627 11204 22636
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 7288 22516 7340 22568
rect 7380 22516 7432 22568
rect 13636 22584 13688 22636
rect 14648 22584 14700 22636
rect 16580 22584 16632 22636
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 21088 22652 21140 22704
rect 24032 22652 24084 22704
rect 24584 22652 24636 22704
rect 25780 22652 25832 22704
rect 26332 22695 26384 22704
rect 26332 22661 26341 22695
rect 26341 22661 26375 22695
rect 26375 22661 26384 22695
rect 26332 22652 26384 22661
rect 26608 22720 26660 22772
rect 27804 22652 27856 22704
rect 29276 22652 29328 22704
rect 29460 22652 29512 22704
rect 30472 22720 30524 22772
rect 35256 22720 35308 22772
rect 35440 22763 35492 22772
rect 35440 22729 35449 22763
rect 35449 22729 35483 22763
rect 35483 22729 35492 22763
rect 35440 22720 35492 22729
rect 35532 22720 35584 22772
rect 36360 22720 36412 22772
rect 37280 22720 37332 22772
rect 37464 22763 37516 22772
rect 37464 22729 37473 22763
rect 37473 22729 37507 22763
rect 37507 22729 37516 22763
rect 37464 22720 37516 22729
rect 38292 22720 38344 22772
rect 38844 22720 38896 22772
rect 39488 22763 39540 22772
rect 39488 22729 39497 22763
rect 39497 22729 39531 22763
rect 39531 22729 39540 22763
rect 39488 22720 39540 22729
rect 39764 22763 39816 22772
rect 39764 22729 39773 22763
rect 39773 22729 39807 22763
rect 39807 22729 39816 22763
rect 39764 22720 39816 22729
rect 21640 22627 21692 22636
rect 21640 22593 21649 22627
rect 21649 22593 21683 22627
rect 21683 22593 21692 22627
rect 21640 22584 21692 22593
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 23572 22584 23624 22636
rect 24400 22627 24452 22636
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 15476 22516 15528 22568
rect 17500 22516 17552 22568
rect 18880 22559 18932 22568
rect 18880 22525 18889 22559
rect 18889 22525 18923 22559
rect 18923 22525 18932 22559
rect 18880 22516 18932 22525
rect 19064 22516 19116 22568
rect 19248 22516 19300 22568
rect 19708 22559 19760 22568
rect 19708 22525 19717 22559
rect 19717 22525 19751 22559
rect 19751 22525 19760 22559
rect 19708 22516 19760 22525
rect 2780 22448 2832 22500
rect 6368 22448 6420 22500
rect 9128 22448 9180 22500
rect 11244 22448 11296 22500
rect 2964 22380 3016 22432
rect 6000 22380 6052 22432
rect 11980 22448 12032 22500
rect 12348 22423 12400 22432
rect 12348 22389 12357 22423
rect 12357 22389 12391 22423
rect 12391 22389 12400 22423
rect 12348 22380 12400 22389
rect 14096 22380 14148 22432
rect 14556 22423 14608 22432
rect 14556 22389 14565 22423
rect 14565 22389 14599 22423
rect 14599 22389 14608 22423
rect 14556 22380 14608 22389
rect 20812 22448 20864 22500
rect 26608 22627 26660 22636
rect 26608 22593 26617 22627
rect 26617 22593 26651 22627
rect 26651 22593 26660 22627
rect 26608 22584 26660 22593
rect 27712 22584 27764 22636
rect 31392 22652 31444 22704
rect 30656 22627 30708 22636
rect 30656 22593 30665 22627
rect 30665 22593 30699 22627
rect 30699 22593 30708 22627
rect 30656 22584 30708 22593
rect 33600 22652 33652 22704
rect 31668 22627 31720 22636
rect 31668 22593 31677 22627
rect 31677 22593 31711 22627
rect 31711 22593 31720 22627
rect 31668 22584 31720 22593
rect 33416 22584 33468 22636
rect 34244 22652 34296 22704
rect 34520 22652 34572 22704
rect 36360 22584 36412 22636
rect 25780 22516 25832 22568
rect 27620 22516 27672 22568
rect 28080 22559 28132 22568
rect 28080 22525 28089 22559
rect 28089 22525 28123 22559
rect 28123 22525 28132 22559
rect 28080 22516 28132 22525
rect 29184 22516 29236 22568
rect 24216 22448 24268 22500
rect 27344 22491 27396 22500
rect 27344 22457 27353 22491
rect 27353 22457 27387 22491
rect 27387 22457 27396 22491
rect 27344 22448 27396 22457
rect 27436 22448 27488 22500
rect 29920 22516 29972 22568
rect 20996 22380 21048 22432
rect 24032 22380 24084 22432
rect 24584 22380 24636 22432
rect 24768 22380 24820 22432
rect 24860 22423 24912 22432
rect 24860 22389 24869 22423
rect 24869 22389 24903 22423
rect 24903 22389 24912 22423
rect 24860 22380 24912 22389
rect 25780 22380 25832 22432
rect 27252 22380 27304 22432
rect 27896 22380 27948 22432
rect 31024 22448 31076 22500
rect 33968 22559 34020 22568
rect 33968 22525 33977 22559
rect 33977 22525 34011 22559
rect 34011 22525 34020 22559
rect 33968 22516 34020 22525
rect 36268 22516 36320 22568
rect 37648 22652 37700 22704
rect 38660 22652 38712 22704
rect 40224 22584 40276 22636
rect 47032 22763 47084 22772
rect 47032 22729 47041 22763
rect 47041 22729 47075 22763
rect 47075 22729 47084 22763
rect 47032 22720 47084 22729
rect 40868 22652 40920 22704
rect 41328 22584 41380 22636
rect 42064 22627 42116 22636
rect 42064 22593 42073 22627
rect 42073 22593 42107 22627
rect 42107 22593 42116 22627
rect 42064 22584 42116 22593
rect 42616 22627 42668 22636
rect 42616 22593 42625 22627
rect 42625 22593 42659 22627
rect 42659 22593 42668 22627
rect 42616 22584 42668 22593
rect 43720 22695 43772 22704
rect 43720 22661 43729 22695
rect 43729 22661 43763 22695
rect 43763 22661 43772 22695
rect 43720 22652 43772 22661
rect 44088 22652 44140 22704
rect 44272 22652 44324 22704
rect 47768 22720 47820 22772
rect 48596 22720 48648 22772
rect 45192 22584 45244 22636
rect 45744 22627 45796 22636
rect 45744 22593 45753 22627
rect 45753 22593 45787 22627
rect 45787 22593 45796 22627
rect 45744 22584 45796 22593
rect 47216 22627 47268 22636
rect 47216 22593 47225 22627
rect 47225 22593 47259 22627
rect 47259 22593 47268 22627
rect 47216 22584 47268 22593
rect 49240 22584 49292 22636
rect 31484 22423 31536 22432
rect 31484 22389 31493 22423
rect 31493 22389 31527 22423
rect 31527 22389 31536 22423
rect 31484 22380 31536 22389
rect 33692 22448 33744 22500
rect 36636 22448 36688 22500
rect 36912 22448 36964 22500
rect 43720 22516 43772 22568
rect 47676 22516 47728 22568
rect 49424 22516 49476 22568
rect 35072 22380 35124 22432
rect 38568 22380 38620 22432
rect 38936 22380 38988 22432
rect 43444 22448 43496 22500
rect 45560 22491 45612 22500
rect 45560 22457 45569 22491
rect 45569 22457 45603 22491
rect 45603 22457 45612 22491
rect 45560 22448 45612 22457
rect 40040 22423 40092 22432
rect 40040 22389 40049 22423
rect 40049 22389 40083 22423
rect 40083 22389 40092 22423
rect 40040 22380 40092 22389
rect 40132 22380 40184 22432
rect 40868 22380 40920 22432
rect 41236 22423 41288 22432
rect 41236 22389 41245 22423
rect 41245 22389 41279 22423
rect 41279 22389 41288 22423
rect 41236 22380 41288 22389
rect 41880 22423 41932 22432
rect 41880 22389 41889 22423
rect 41889 22389 41923 22423
rect 41923 22389 41932 22423
rect 41880 22380 41932 22389
rect 43536 22380 43588 22432
rect 48412 22423 48464 22432
rect 48412 22389 48421 22423
rect 48421 22389 48455 22423
rect 48455 22389 48464 22423
rect 48412 22380 48464 22389
rect 48504 22380 48556 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 4252 22176 4304 22228
rect 11888 22176 11940 22228
rect 3976 22108 4028 22160
rect 1032 21904 1084 21956
rect 6828 21972 6880 22024
rect 9680 22040 9732 22092
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 11980 22040 12032 22092
rect 3240 21904 3292 21956
rect 5632 21904 5684 21956
rect 8484 21904 8536 21956
rect 6736 21836 6788 21888
rect 8392 21879 8444 21888
rect 8392 21845 8401 21879
rect 8401 21845 8435 21879
rect 8435 21845 8444 21879
rect 8392 21836 8444 21845
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 13268 22040 13320 22092
rect 15476 22176 15528 22228
rect 16580 22176 16632 22228
rect 17224 22176 17276 22228
rect 18788 22176 18840 22228
rect 20812 22176 20864 22228
rect 21640 22176 21692 22228
rect 23020 22176 23072 22228
rect 23572 22176 23624 22228
rect 17040 22108 17092 22160
rect 14280 22040 14332 22092
rect 19892 22108 19944 22160
rect 13544 21972 13596 22024
rect 16948 22015 17000 22024
rect 16948 21981 16957 22015
rect 16957 21981 16991 22015
rect 16991 21981 17000 22015
rect 16948 21972 17000 21981
rect 21916 22040 21968 22092
rect 24308 22108 24360 22160
rect 25136 22176 25188 22228
rect 26700 22176 26752 22228
rect 27160 22219 27212 22228
rect 27160 22185 27169 22219
rect 27169 22185 27203 22219
rect 27203 22185 27212 22219
rect 27160 22176 27212 22185
rect 27896 22176 27948 22228
rect 29000 22176 29052 22228
rect 29460 22176 29512 22228
rect 30012 22176 30064 22228
rect 30196 22176 30248 22228
rect 32128 22176 32180 22228
rect 33600 22176 33652 22228
rect 34704 22176 34756 22228
rect 37464 22176 37516 22228
rect 38660 22176 38712 22228
rect 22652 22040 22704 22092
rect 24860 22108 24912 22160
rect 24768 22040 24820 22092
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 22376 21972 22428 22024
rect 22836 21972 22888 22024
rect 13268 21904 13320 21956
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 13912 21836 13964 21888
rect 14096 21879 14148 21888
rect 14096 21845 14105 21879
rect 14105 21845 14139 21879
rect 14139 21845 14148 21879
rect 14096 21836 14148 21845
rect 14648 21947 14700 21956
rect 14648 21913 14657 21947
rect 14657 21913 14691 21947
rect 14691 21913 14700 21947
rect 14648 21904 14700 21913
rect 15292 21904 15344 21956
rect 16580 21904 16632 21956
rect 17132 21904 17184 21956
rect 18880 21904 18932 21956
rect 18972 21904 19024 21956
rect 20628 21904 20680 21956
rect 21088 21836 21140 21888
rect 23940 21972 23992 22024
rect 24952 21972 25004 22024
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 25228 22040 25280 22092
rect 28264 22108 28316 22160
rect 26608 22083 26660 22092
rect 26608 22049 26617 22083
rect 26617 22049 26651 22083
rect 26651 22049 26660 22083
rect 26608 22040 26660 22049
rect 27528 22040 27580 22092
rect 28080 22040 28132 22092
rect 28908 22083 28960 22092
rect 28908 22049 28917 22083
rect 28917 22049 28951 22083
rect 28951 22049 28960 22083
rect 28908 22040 28960 22049
rect 29184 22040 29236 22092
rect 29460 22040 29512 22092
rect 25872 21972 25924 22024
rect 27436 21972 27488 22024
rect 27620 22015 27672 22024
rect 27620 21981 27629 22015
rect 27629 21981 27663 22015
rect 27663 21981 27672 22015
rect 27620 21972 27672 21981
rect 30564 22040 30616 22092
rect 31484 22040 31536 22092
rect 35440 22108 35492 22160
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 30840 22015 30892 22024
rect 30840 21981 30849 22015
rect 30849 21981 30883 22015
rect 30883 21981 30892 22015
rect 30840 21972 30892 21981
rect 32404 21972 32456 22024
rect 34520 22040 34572 22092
rect 35072 22083 35124 22092
rect 35072 22049 35081 22083
rect 35081 22049 35115 22083
rect 35115 22049 35124 22083
rect 35072 22040 35124 22049
rect 37832 22108 37884 22160
rect 39488 22108 39540 22160
rect 40500 22176 40552 22228
rect 41420 22219 41472 22228
rect 41420 22185 41429 22219
rect 41429 22185 41463 22219
rect 41463 22185 41472 22219
rect 41420 22176 41472 22185
rect 43536 22176 43588 22228
rect 45192 22219 45244 22228
rect 45192 22185 45201 22219
rect 45201 22185 45235 22219
rect 45235 22185 45244 22219
rect 45192 22176 45244 22185
rect 45376 22219 45428 22228
rect 45376 22185 45385 22219
rect 45385 22185 45419 22219
rect 45419 22185 45428 22219
rect 45376 22176 45428 22185
rect 45744 22176 45796 22228
rect 46848 22176 46900 22228
rect 47584 22219 47636 22228
rect 47584 22185 47593 22219
rect 47593 22185 47627 22219
rect 47627 22185 47636 22219
rect 47584 22176 47636 22185
rect 34244 21972 34296 22024
rect 38476 22040 38528 22092
rect 38844 22083 38896 22092
rect 38844 22049 38853 22083
rect 38853 22049 38887 22083
rect 38887 22049 38896 22083
rect 38844 22040 38896 22049
rect 40500 22040 40552 22092
rect 40960 22040 41012 22092
rect 41144 22040 41196 22092
rect 37464 21972 37516 22024
rect 37740 21972 37792 22024
rect 41880 22040 41932 22092
rect 42064 22108 42116 22160
rect 42708 22108 42760 22160
rect 42156 22040 42208 22092
rect 43260 22040 43312 22092
rect 45100 22040 45152 22092
rect 24584 21904 24636 21956
rect 24768 21904 24820 21956
rect 22468 21836 22520 21888
rect 22560 21836 22612 21888
rect 22836 21836 22888 21888
rect 23756 21836 23808 21888
rect 24032 21836 24084 21888
rect 24676 21836 24728 21888
rect 24860 21836 24912 21888
rect 28356 21904 28408 21956
rect 27620 21836 27672 21888
rect 30472 21904 30524 21956
rect 30748 21904 30800 21956
rect 31392 21904 31444 21956
rect 32772 21904 32824 21956
rect 33876 21904 33928 21956
rect 37004 21904 37056 21956
rect 37280 21904 37332 21956
rect 29184 21836 29236 21888
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 30380 21879 30432 21888
rect 30380 21845 30389 21879
rect 30389 21845 30423 21879
rect 30423 21845 30432 21879
rect 30380 21836 30432 21845
rect 30564 21836 30616 21888
rect 31944 21836 31996 21888
rect 32036 21836 32088 21888
rect 32588 21879 32640 21888
rect 32588 21845 32597 21879
rect 32597 21845 32631 21879
rect 32631 21845 32640 21879
rect 32588 21836 32640 21845
rect 32680 21836 32732 21888
rect 33416 21879 33468 21888
rect 33416 21845 33425 21879
rect 33425 21845 33459 21879
rect 33459 21845 33468 21879
rect 33416 21836 33468 21845
rect 34336 21879 34388 21888
rect 34336 21845 34345 21879
rect 34345 21845 34379 21879
rect 34379 21845 34388 21879
rect 34336 21836 34388 21845
rect 35256 21879 35308 21888
rect 35256 21845 35265 21879
rect 35265 21845 35299 21879
rect 35299 21845 35308 21879
rect 35256 21836 35308 21845
rect 35992 21836 36044 21888
rect 36268 21836 36320 21888
rect 36820 21879 36872 21888
rect 36820 21845 36829 21879
rect 36829 21845 36863 21879
rect 36863 21845 36872 21879
rect 36820 21836 36872 21845
rect 37372 21879 37424 21888
rect 37372 21845 37381 21879
rect 37381 21845 37415 21879
rect 37415 21845 37424 21879
rect 37372 21836 37424 21845
rect 41512 21972 41564 22024
rect 42524 21972 42576 22024
rect 42984 21972 43036 22024
rect 43720 21972 43772 22024
rect 43812 22015 43864 22024
rect 43812 21981 43821 22015
rect 43821 21981 43855 22015
rect 43855 21981 43864 22015
rect 43812 21972 43864 21981
rect 44088 22015 44140 22024
rect 44088 21981 44097 22015
rect 44097 21981 44131 22015
rect 44131 21981 44140 22015
rect 44088 21972 44140 21981
rect 39580 21879 39632 21888
rect 39580 21845 39589 21879
rect 39589 21845 39623 21879
rect 39623 21845 39632 21879
rect 39856 21879 39908 21888
rect 39580 21836 39632 21845
rect 39856 21845 39865 21879
rect 39865 21845 39899 21879
rect 39899 21845 39908 21879
rect 39856 21836 39908 21845
rect 39948 21836 40000 21888
rect 40960 21904 41012 21956
rect 41512 21836 41564 21888
rect 42156 21836 42208 21888
rect 42248 21836 42300 21888
rect 43260 21836 43312 21888
rect 45100 21836 45152 21888
rect 46112 21972 46164 22024
rect 47492 21972 47544 22024
rect 47584 21904 47636 21956
rect 47860 21904 47912 21956
rect 49240 21947 49292 21956
rect 49240 21913 49249 21947
rect 49249 21913 49283 21947
rect 49283 21913 49292 21947
rect 49240 21904 49292 21913
rect 48780 21879 48832 21888
rect 48780 21845 48789 21879
rect 48789 21845 48823 21879
rect 48823 21845 48832 21879
rect 48780 21836 48832 21845
rect 48872 21836 48924 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 6736 21632 6788 21684
rect 3332 21564 3384 21616
rect 7196 21564 7248 21616
rect 9496 21632 9548 21684
rect 12532 21632 12584 21684
rect 13728 21632 13780 21684
rect 14096 21632 14148 21684
rect 1768 21471 1820 21480
rect 1768 21437 1777 21471
rect 1777 21437 1811 21471
rect 1811 21437 1820 21471
rect 1768 21428 1820 21437
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 6552 21496 6604 21548
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 5632 21428 5684 21480
rect 5816 21428 5868 21480
rect 11428 21564 11480 21616
rect 11704 21607 11756 21616
rect 11704 21573 11713 21607
rect 11713 21573 11747 21607
rect 11747 21573 11756 21607
rect 11704 21564 11756 21573
rect 9588 21496 9640 21548
rect 9956 21496 10008 21548
rect 10968 21496 11020 21548
rect 12348 21539 12400 21548
rect 12348 21505 12357 21539
rect 12357 21505 12391 21539
rect 12391 21505 12400 21539
rect 12348 21496 12400 21505
rect 12624 21564 12676 21616
rect 14188 21564 14240 21616
rect 14280 21564 14332 21616
rect 16672 21632 16724 21684
rect 17408 21675 17460 21684
rect 17408 21641 17417 21675
rect 17417 21641 17451 21675
rect 17451 21641 17460 21675
rect 17408 21632 17460 21641
rect 17868 21675 17920 21684
rect 17868 21641 17877 21675
rect 17877 21641 17911 21675
rect 17911 21641 17920 21675
rect 17868 21632 17920 21641
rect 15292 21564 15344 21616
rect 17224 21564 17276 21616
rect 19800 21632 19852 21684
rect 22468 21632 22520 21684
rect 25780 21632 25832 21684
rect 14004 21496 14056 21548
rect 14372 21496 14424 21548
rect 18328 21496 18380 21548
rect 3792 21292 3844 21344
rect 12440 21428 12492 21480
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 18788 21564 18840 21616
rect 20720 21564 20772 21616
rect 23020 21564 23072 21616
rect 23204 21564 23256 21616
rect 24032 21564 24084 21616
rect 27436 21632 27488 21684
rect 27804 21632 27856 21684
rect 28816 21675 28868 21684
rect 28816 21641 28825 21675
rect 28825 21641 28859 21675
rect 28859 21641 28868 21675
rect 28816 21632 28868 21641
rect 30012 21632 30064 21684
rect 31392 21632 31444 21684
rect 31760 21632 31812 21684
rect 32404 21632 32456 21684
rect 33416 21632 33468 21684
rect 29460 21564 29512 21616
rect 20904 21496 20956 21548
rect 21364 21539 21416 21548
rect 21364 21505 21373 21539
rect 21373 21505 21407 21539
rect 21407 21505 21416 21539
rect 21364 21496 21416 21505
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25136 21496 25188 21505
rect 26148 21496 26200 21548
rect 11796 21360 11848 21412
rect 11704 21292 11756 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 12808 21292 12860 21344
rect 16856 21360 16908 21412
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 18972 21428 19024 21480
rect 16580 21292 16632 21344
rect 21456 21360 21508 21412
rect 22192 21428 22244 21480
rect 24216 21428 24268 21480
rect 25320 21428 25372 21480
rect 25412 21471 25464 21480
rect 25412 21437 25421 21471
rect 25421 21437 25455 21471
rect 25455 21437 25464 21471
rect 25412 21428 25464 21437
rect 27896 21496 27948 21548
rect 30656 21564 30708 21616
rect 31208 21607 31260 21616
rect 31208 21573 31217 21607
rect 31217 21573 31251 21607
rect 31251 21573 31260 21607
rect 31208 21564 31260 21573
rect 29920 21539 29972 21548
rect 29920 21505 29929 21539
rect 29929 21505 29963 21539
rect 29963 21505 29972 21539
rect 29920 21496 29972 21505
rect 30932 21496 30984 21548
rect 28908 21471 28960 21480
rect 28908 21437 28917 21471
rect 28917 21437 28951 21471
rect 28951 21437 28960 21471
rect 28908 21428 28960 21437
rect 26424 21403 26476 21412
rect 26424 21369 26433 21403
rect 26433 21369 26467 21403
rect 26467 21369 26476 21403
rect 26424 21360 26476 21369
rect 26884 21360 26936 21412
rect 30472 21428 30524 21480
rect 29920 21360 29972 21412
rect 31116 21360 31168 21412
rect 19340 21292 19392 21344
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 21640 21292 21692 21344
rect 26148 21292 26200 21344
rect 26240 21292 26292 21344
rect 26976 21292 27028 21344
rect 29552 21335 29604 21344
rect 29552 21301 29561 21335
rect 29561 21301 29595 21335
rect 29595 21301 29604 21335
rect 29552 21292 29604 21301
rect 30748 21335 30800 21344
rect 30748 21301 30757 21335
rect 30757 21301 30791 21335
rect 30791 21301 30800 21335
rect 30748 21292 30800 21301
rect 31944 21496 31996 21548
rect 33416 21496 33468 21548
rect 33508 21539 33560 21548
rect 33508 21505 33517 21539
rect 33517 21505 33551 21539
rect 33551 21505 33560 21539
rect 33508 21496 33560 21505
rect 33324 21471 33376 21480
rect 33324 21437 33333 21471
rect 33333 21437 33367 21471
rect 33367 21437 33376 21471
rect 33324 21428 33376 21437
rect 34612 21632 34664 21684
rect 34704 21675 34756 21684
rect 34704 21641 34713 21675
rect 34713 21641 34747 21675
rect 34747 21641 34756 21675
rect 34704 21632 34756 21641
rect 34796 21675 34848 21684
rect 34796 21641 34805 21675
rect 34805 21641 34839 21675
rect 34839 21641 34848 21675
rect 34796 21632 34848 21641
rect 35256 21632 35308 21684
rect 37740 21632 37792 21684
rect 38384 21632 38436 21684
rect 38292 21564 38344 21616
rect 38568 21564 38620 21616
rect 36820 21496 36872 21548
rect 37004 21496 37056 21548
rect 37280 21539 37332 21548
rect 37280 21505 37289 21539
rect 37289 21505 37323 21539
rect 37323 21505 37332 21539
rect 37280 21496 37332 21505
rect 39856 21632 39908 21684
rect 42064 21632 42116 21684
rect 42524 21675 42576 21684
rect 42524 21641 42533 21675
rect 42533 21641 42567 21675
rect 42567 21641 42576 21675
rect 42524 21632 42576 21641
rect 43720 21675 43772 21684
rect 43720 21641 43729 21675
rect 43729 21641 43763 21675
rect 43763 21641 43772 21675
rect 43720 21632 43772 21641
rect 44272 21675 44324 21684
rect 44272 21641 44281 21675
rect 44281 21641 44315 21675
rect 44315 21641 44324 21675
rect 44272 21632 44324 21641
rect 44456 21675 44508 21684
rect 44456 21641 44465 21675
rect 44465 21641 44499 21675
rect 44499 21641 44508 21675
rect 44456 21632 44508 21641
rect 45928 21632 45980 21684
rect 47860 21675 47912 21684
rect 47860 21641 47869 21675
rect 47869 21641 47903 21675
rect 47903 21641 47912 21675
rect 47860 21632 47912 21641
rect 40592 21564 40644 21616
rect 40776 21564 40828 21616
rect 40868 21564 40920 21616
rect 47676 21564 47728 21616
rect 47400 21496 47452 21548
rect 48228 21496 48280 21548
rect 49332 21539 49384 21548
rect 49332 21505 49341 21539
rect 49341 21505 49375 21539
rect 49375 21505 49384 21539
rect 49332 21496 49384 21505
rect 36176 21471 36228 21480
rect 36176 21437 36185 21471
rect 36185 21437 36219 21471
rect 36219 21437 36228 21471
rect 36176 21428 36228 21437
rect 34428 21360 34480 21412
rect 36452 21428 36504 21480
rect 36912 21428 36964 21480
rect 37556 21428 37608 21480
rect 38292 21471 38344 21480
rect 37372 21360 37424 21412
rect 38292 21437 38301 21471
rect 38301 21437 38335 21471
rect 38335 21437 38344 21471
rect 38292 21428 38344 21437
rect 38384 21428 38436 21480
rect 40040 21428 40092 21480
rect 40868 21428 40920 21480
rect 41512 21471 41564 21480
rect 41512 21437 41521 21471
rect 41521 21437 41555 21471
rect 41555 21437 41564 21471
rect 41512 21428 41564 21437
rect 41880 21428 41932 21480
rect 43812 21428 43864 21480
rect 46112 21428 46164 21480
rect 49240 21428 49292 21480
rect 39304 21360 39356 21412
rect 40960 21360 41012 21412
rect 33968 21335 34020 21344
rect 33968 21301 33977 21335
rect 33977 21301 34011 21335
rect 34011 21301 34020 21335
rect 33968 21292 34020 21301
rect 35624 21292 35676 21344
rect 35716 21335 35768 21344
rect 35716 21301 35725 21335
rect 35725 21301 35759 21335
rect 35759 21301 35768 21335
rect 35716 21292 35768 21301
rect 37556 21335 37608 21344
rect 37556 21301 37565 21335
rect 37565 21301 37599 21335
rect 37599 21301 37608 21335
rect 37556 21292 37608 21301
rect 37832 21292 37884 21344
rect 40868 21292 40920 21344
rect 41420 21292 41472 21344
rect 43444 21292 43496 21344
rect 48320 21292 48372 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 7196 21088 7248 21140
rect 9220 21131 9272 21140
rect 9220 21097 9229 21131
rect 9229 21097 9263 21131
rect 9263 21097 9272 21131
rect 9220 21088 9272 21097
rect 12256 21088 12308 21140
rect 12440 21131 12492 21140
rect 12440 21097 12449 21131
rect 12449 21097 12483 21131
rect 12483 21097 12492 21131
rect 12440 21088 12492 21097
rect 13360 21088 13412 21140
rect 14280 21131 14332 21140
rect 14280 21097 14289 21131
rect 14289 21097 14323 21131
rect 14323 21097 14332 21131
rect 14280 21088 14332 21097
rect 14372 21088 14424 21140
rect 15752 21088 15804 21140
rect 16304 21088 16356 21140
rect 19708 21088 19760 21140
rect 19800 21088 19852 21140
rect 2872 20952 2924 21004
rect 4160 20995 4212 21004
rect 4160 20961 4169 20995
rect 4169 20961 4203 20995
rect 4203 20961 4212 20995
rect 4160 20952 4212 20961
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 9588 20952 9640 21004
rect 12716 21063 12768 21072
rect 12716 21029 12725 21063
rect 12725 21029 12759 21063
rect 12759 21029 12768 21063
rect 12716 21020 12768 21029
rect 13452 20952 13504 21004
rect 8392 20927 8444 20936
rect 8392 20893 8401 20927
rect 8401 20893 8435 20927
rect 8435 20893 8444 20927
rect 8392 20884 8444 20893
rect 11060 20884 11112 20936
rect 11336 20927 11388 20936
rect 11336 20893 11345 20927
rect 11345 20893 11379 20927
rect 11379 20893 11388 20927
rect 11336 20884 11388 20893
rect 11796 20884 11848 20936
rect 8484 20816 8536 20868
rect 10876 20748 10928 20800
rect 11152 20791 11204 20800
rect 11152 20757 11161 20791
rect 11161 20757 11195 20791
rect 11195 20757 11204 20791
rect 11152 20748 11204 20757
rect 12072 20884 12124 20936
rect 16672 21020 16724 21072
rect 17500 21020 17552 21072
rect 19064 21020 19116 21072
rect 24124 21088 24176 21140
rect 26056 21088 26108 21140
rect 29644 21088 29696 21140
rect 30012 21088 30064 21140
rect 23940 21020 23992 21072
rect 26516 21020 26568 21072
rect 29552 21020 29604 21072
rect 29828 21020 29880 21072
rect 16856 20884 16908 20936
rect 17500 20884 17552 20936
rect 19340 20884 19392 20936
rect 12624 20816 12676 20868
rect 13176 20816 13228 20868
rect 14096 20816 14148 20868
rect 16120 20816 16172 20868
rect 13820 20748 13872 20800
rect 13912 20748 13964 20800
rect 16764 20748 16816 20800
rect 19432 20816 19484 20868
rect 18512 20748 18564 20800
rect 19800 20884 19852 20936
rect 22560 20952 22612 21004
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 23296 20952 23348 21004
rect 24216 20995 24268 21004
rect 24216 20961 24225 20995
rect 24225 20961 24259 20995
rect 24259 20961 24268 20995
rect 24216 20952 24268 20961
rect 25596 20952 25648 21004
rect 26332 20952 26384 21004
rect 22928 20927 22980 20936
rect 22928 20893 22937 20927
rect 22937 20893 22971 20927
rect 22971 20893 22980 20927
rect 22928 20884 22980 20893
rect 24124 20884 24176 20936
rect 27436 20927 27488 20936
rect 27436 20893 27445 20927
rect 27445 20893 27479 20927
rect 27479 20893 27488 20927
rect 27436 20884 27488 20893
rect 27896 20995 27948 21004
rect 27896 20961 27905 20995
rect 27905 20961 27939 20995
rect 27939 20961 27948 20995
rect 27896 20952 27948 20961
rect 35716 21088 35768 21140
rect 36636 21088 36688 21140
rect 34244 21063 34296 21072
rect 34244 21029 34253 21063
rect 34253 21029 34287 21063
rect 34287 21029 34296 21063
rect 34244 21020 34296 21029
rect 40316 21088 40368 21140
rect 42248 21088 42300 21140
rect 42800 21088 42852 21140
rect 43352 21088 43404 21140
rect 47768 21088 47820 21140
rect 40684 21020 40736 21072
rect 42708 21020 42760 21072
rect 29552 20884 29604 20936
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 32312 20952 32364 21004
rect 32864 20952 32916 21004
rect 34336 20952 34388 21004
rect 32036 20884 32088 20936
rect 32496 20927 32548 20936
rect 32496 20893 32505 20927
rect 32505 20893 32539 20927
rect 32539 20893 32548 20927
rect 32496 20884 32548 20893
rect 34520 20884 34572 20936
rect 35072 20884 35124 20936
rect 37556 20952 37608 21004
rect 39488 20952 39540 21004
rect 39672 20952 39724 21004
rect 21364 20816 21416 20868
rect 23572 20859 23624 20868
rect 23572 20825 23581 20859
rect 23581 20825 23615 20859
rect 23615 20825 23624 20859
rect 23572 20816 23624 20825
rect 19616 20791 19668 20800
rect 19616 20757 19625 20791
rect 19625 20757 19659 20791
rect 19659 20757 19668 20791
rect 19616 20748 19668 20757
rect 25228 20816 25280 20868
rect 25780 20748 25832 20800
rect 26792 20816 26844 20868
rect 27712 20816 27764 20868
rect 26516 20748 26568 20800
rect 26976 20748 27028 20800
rect 27068 20748 27120 20800
rect 28724 20791 28776 20800
rect 28724 20757 28733 20791
rect 28733 20757 28767 20791
rect 28767 20757 28776 20791
rect 28724 20748 28776 20757
rect 30104 20748 30156 20800
rect 30932 20816 30984 20868
rect 31760 20816 31812 20868
rect 32404 20816 32456 20868
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 31300 20748 31352 20800
rect 34428 20748 34480 20800
rect 36452 20816 36504 20868
rect 36728 20816 36780 20868
rect 38384 20816 38436 20868
rect 40684 20884 40736 20936
rect 41328 20884 41380 20936
rect 41604 20884 41656 20936
rect 41972 20952 42024 21004
rect 47124 20884 47176 20936
rect 47860 20884 47912 20936
rect 48780 20884 48832 20936
rect 49332 20927 49384 20936
rect 49332 20893 49341 20927
rect 49341 20893 49375 20927
rect 49375 20893 49384 20927
rect 49332 20884 49384 20893
rect 36636 20748 36688 20800
rect 36912 20791 36964 20800
rect 36912 20757 36921 20791
rect 36921 20757 36955 20791
rect 36955 20757 36964 20791
rect 36912 20748 36964 20757
rect 37188 20748 37240 20800
rect 37648 20791 37700 20800
rect 37648 20757 37657 20791
rect 37657 20757 37691 20791
rect 37691 20757 37700 20791
rect 37648 20748 37700 20757
rect 37832 20748 37884 20800
rect 40224 20748 40276 20800
rect 40868 20748 40920 20800
rect 41788 20816 41840 20868
rect 42064 20816 42116 20868
rect 46020 20816 46072 20868
rect 41604 20791 41656 20800
rect 41604 20757 41613 20791
rect 41613 20757 41647 20791
rect 41647 20757 41656 20791
rect 41604 20748 41656 20757
rect 43628 20748 43680 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 6644 20544 6696 20596
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 11060 20544 11112 20596
rect 1308 20476 1360 20528
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 5264 20451 5316 20460
rect 5264 20417 5273 20451
rect 5273 20417 5307 20451
rect 5307 20417 5316 20451
rect 5264 20408 5316 20417
rect 6368 20408 6420 20460
rect 6828 20476 6880 20528
rect 5908 20340 5960 20392
rect 9772 20408 9824 20460
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 12532 20476 12584 20528
rect 12808 20476 12860 20528
rect 13452 20476 13504 20528
rect 14924 20587 14976 20596
rect 14924 20553 14933 20587
rect 14933 20553 14967 20587
rect 14967 20553 14976 20587
rect 14924 20544 14976 20553
rect 15568 20587 15620 20596
rect 15568 20553 15577 20587
rect 15577 20553 15611 20587
rect 15611 20553 15620 20587
rect 15568 20544 15620 20553
rect 15660 20544 15712 20596
rect 16028 20587 16080 20596
rect 16028 20553 16037 20587
rect 16037 20553 16071 20587
rect 16071 20553 16080 20587
rect 16028 20544 16080 20553
rect 17132 20544 17184 20596
rect 17500 20544 17552 20596
rect 18880 20544 18932 20596
rect 19432 20544 19484 20596
rect 19892 20544 19944 20596
rect 21364 20544 21416 20596
rect 22928 20544 22980 20596
rect 19064 20519 19116 20528
rect 11060 20340 11112 20392
rect 11888 20451 11940 20460
rect 11888 20417 11897 20451
rect 11897 20417 11931 20451
rect 11931 20417 11940 20451
rect 11888 20408 11940 20417
rect 2780 20272 2832 20324
rect 3332 20272 3384 20324
rect 10784 20272 10836 20324
rect 4160 20204 4212 20256
rect 12532 20340 12584 20392
rect 14280 20383 14332 20392
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 15936 20340 15988 20392
rect 19064 20485 19073 20519
rect 19073 20485 19107 20519
rect 19107 20485 19116 20519
rect 19064 20476 19116 20485
rect 20904 20476 20956 20528
rect 21548 20476 21600 20528
rect 23756 20476 23808 20528
rect 25688 20544 25740 20596
rect 25780 20544 25832 20596
rect 27068 20544 27120 20596
rect 16856 20408 16908 20460
rect 22192 20408 22244 20460
rect 23388 20451 23440 20460
rect 23388 20417 23397 20451
rect 23397 20417 23431 20451
rect 23431 20417 23440 20451
rect 23388 20408 23440 20417
rect 24216 20476 24268 20528
rect 20168 20340 20220 20392
rect 21548 20340 21600 20392
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 16856 20272 16908 20324
rect 11796 20204 11848 20256
rect 12808 20204 12860 20256
rect 13176 20247 13228 20256
rect 13176 20213 13185 20247
rect 13185 20213 13219 20247
rect 13219 20213 13228 20247
rect 13176 20204 13228 20213
rect 15476 20204 15528 20256
rect 17040 20204 17092 20256
rect 17132 20204 17184 20256
rect 19616 20204 19668 20256
rect 22284 20272 22336 20324
rect 24676 20340 24728 20392
rect 26884 20476 26936 20528
rect 26056 20451 26108 20460
rect 26056 20417 26065 20451
rect 26065 20417 26099 20451
rect 26099 20417 26108 20451
rect 26056 20408 26108 20417
rect 30840 20544 30892 20596
rect 31484 20544 31536 20596
rect 32496 20544 32548 20596
rect 34060 20544 34112 20596
rect 36176 20544 36228 20596
rect 36452 20544 36504 20596
rect 37464 20544 37516 20596
rect 47860 20544 47912 20596
rect 28908 20476 28960 20528
rect 29184 20476 29236 20528
rect 31024 20519 31076 20528
rect 31024 20485 31033 20519
rect 31033 20485 31067 20519
rect 31067 20485 31076 20519
rect 31024 20476 31076 20485
rect 31300 20476 31352 20528
rect 32128 20476 32180 20528
rect 32404 20476 32456 20528
rect 33692 20476 33744 20528
rect 34428 20476 34480 20528
rect 30196 20408 30248 20460
rect 26148 20340 26200 20392
rect 29276 20340 29328 20392
rect 29552 20383 29604 20392
rect 29552 20349 29561 20383
rect 29561 20349 29595 20383
rect 29595 20349 29604 20383
rect 29552 20340 29604 20349
rect 22744 20272 22796 20324
rect 26056 20272 26108 20324
rect 20628 20204 20680 20256
rect 21364 20204 21416 20256
rect 21548 20204 21600 20256
rect 24860 20204 24912 20256
rect 25596 20247 25648 20256
rect 25596 20213 25605 20247
rect 25605 20213 25639 20247
rect 25639 20213 25648 20247
rect 25596 20204 25648 20213
rect 26516 20204 26568 20256
rect 28908 20272 28960 20324
rect 30564 20340 30616 20392
rect 31116 20340 31168 20392
rect 32496 20408 32548 20460
rect 36728 20476 36780 20528
rect 37372 20476 37424 20528
rect 37924 20476 37976 20528
rect 39764 20476 39816 20528
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 34060 20383 34112 20392
rect 34060 20349 34069 20383
rect 34069 20349 34103 20383
rect 34103 20349 34112 20383
rect 34060 20340 34112 20349
rect 34888 20451 34940 20460
rect 34888 20417 34897 20451
rect 34897 20417 34931 20451
rect 34931 20417 34940 20451
rect 34888 20408 34940 20417
rect 35072 20408 35124 20460
rect 36452 20451 36504 20460
rect 36452 20417 36461 20451
rect 36461 20417 36495 20451
rect 36495 20417 36504 20451
rect 36452 20408 36504 20417
rect 37188 20408 37240 20460
rect 39488 20451 39540 20460
rect 39488 20417 39497 20451
rect 39497 20417 39531 20451
rect 39531 20417 39540 20451
rect 39488 20408 39540 20417
rect 39672 20408 39724 20460
rect 34980 20340 35032 20392
rect 31944 20315 31996 20324
rect 31944 20281 31953 20315
rect 31953 20281 31987 20315
rect 31987 20281 31996 20315
rect 31944 20272 31996 20281
rect 30564 20204 30616 20256
rect 30840 20204 30892 20256
rect 31392 20204 31444 20256
rect 35532 20315 35584 20324
rect 35532 20281 35541 20315
rect 35541 20281 35575 20315
rect 35575 20281 35584 20315
rect 35532 20272 35584 20281
rect 35992 20272 36044 20324
rect 37464 20340 37516 20392
rect 37648 20340 37700 20392
rect 40132 20383 40184 20392
rect 40132 20349 40141 20383
rect 40141 20349 40175 20383
rect 40175 20349 40184 20383
rect 40132 20340 40184 20349
rect 41052 20340 41104 20392
rect 37648 20204 37700 20256
rect 37740 20247 37792 20256
rect 37740 20213 37749 20247
rect 37749 20213 37783 20247
rect 37783 20213 37792 20247
rect 37740 20204 37792 20213
rect 39212 20204 39264 20256
rect 40684 20247 40736 20256
rect 40684 20213 40693 20247
rect 40693 20213 40727 20247
rect 40727 20213 40736 20247
rect 40684 20204 40736 20213
rect 48780 20408 48832 20460
rect 49424 20408 49476 20460
rect 48320 20204 48372 20256
rect 48412 20247 48464 20256
rect 48412 20213 48421 20247
rect 48421 20213 48455 20247
rect 48455 20213 48464 20247
rect 48412 20204 48464 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 4804 20000 4856 20052
rect 11980 20000 12032 20052
rect 12440 20000 12492 20052
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 5264 19932 5316 19984
rect 8300 19932 8352 19984
rect 9956 19975 10008 19984
rect 9956 19941 9965 19975
rect 9965 19941 9999 19975
rect 9999 19941 10008 19975
rect 9956 19932 10008 19941
rect 10784 19932 10836 19984
rect 18328 20000 18380 20052
rect 4252 19907 4304 19916
rect 4252 19873 4261 19907
rect 4261 19873 4295 19907
rect 4295 19873 4304 19907
rect 4252 19864 4304 19873
rect 5724 19864 5776 19916
rect 3332 19796 3384 19848
rect 5356 19839 5408 19848
rect 5356 19805 5365 19839
rect 5365 19805 5399 19839
rect 5399 19805 5408 19839
rect 5356 19796 5408 19805
rect 1492 19728 1544 19780
rect 9956 19796 10008 19848
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 14924 19975 14976 19984
rect 14924 19941 14933 19975
rect 14933 19941 14967 19975
rect 14967 19941 14976 19975
rect 14924 19932 14976 19941
rect 11428 19771 11480 19780
rect 11428 19737 11437 19771
rect 11437 19737 11471 19771
rect 11471 19737 11480 19771
rect 11428 19728 11480 19737
rect 10876 19660 10928 19712
rect 11704 19728 11756 19780
rect 12900 19728 12952 19780
rect 16304 19907 16356 19916
rect 16304 19873 16313 19907
rect 16313 19873 16347 19907
rect 16347 19873 16356 19907
rect 16304 19864 16356 19873
rect 18880 19932 18932 19984
rect 17592 19864 17644 19916
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 15476 19796 15528 19848
rect 16120 19796 16172 19848
rect 18604 19796 18656 19848
rect 20352 20000 20404 20052
rect 19248 19932 19300 19984
rect 22376 20000 22428 20052
rect 22468 20000 22520 20052
rect 20996 19864 21048 19916
rect 21456 19864 21508 19916
rect 21640 19864 21692 19916
rect 22836 19864 22888 19916
rect 18328 19728 18380 19780
rect 20352 19796 20404 19848
rect 20904 19796 20956 19848
rect 23020 19839 23072 19848
rect 23020 19805 23029 19839
rect 23029 19805 23063 19839
rect 23063 19805 23072 19839
rect 23020 19796 23072 19805
rect 17132 19660 17184 19712
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 17316 19703 17368 19712
rect 17316 19669 17325 19703
rect 17325 19669 17359 19703
rect 17359 19669 17368 19703
rect 17316 19660 17368 19669
rect 20720 19728 20772 19780
rect 22100 19728 22152 19780
rect 22376 19728 22428 19780
rect 23480 19864 23532 19916
rect 23848 19864 23900 19916
rect 25780 19932 25832 19984
rect 24308 19864 24360 19916
rect 24584 19907 24636 19916
rect 24584 19873 24593 19907
rect 24593 19873 24627 19907
rect 24627 19873 24636 19907
rect 24584 19864 24636 19873
rect 25228 19796 25280 19848
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 27068 20000 27120 20052
rect 30380 20000 30432 20052
rect 32772 20000 32824 20052
rect 26884 19864 26936 19916
rect 28908 19932 28960 19984
rect 28356 19864 28408 19916
rect 30012 19864 30064 19916
rect 30196 19907 30248 19916
rect 30196 19873 30205 19907
rect 30205 19873 30239 19907
rect 30239 19873 30248 19907
rect 30196 19864 30248 19873
rect 30288 19907 30340 19916
rect 30288 19873 30297 19907
rect 30297 19873 30331 19907
rect 30331 19873 30340 19907
rect 30288 19864 30340 19873
rect 34336 20000 34388 20052
rect 34888 20000 34940 20052
rect 36912 20000 36964 20052
rect 37832 20000 37884 20052
rect 39948 20000 40000 20052
rect 40500 20000 40552 20052
rect 48780 20043 48832 20052
rect 48780 20009 48789 20043
rect 48789 20009 48823 20043
rect 48823 20009 48832 20043
rect 48780 20000 48832 20009
rect 34704 19932 34756 19984
rect 28632 19796 28684 19848
rect 19064 19660 19116 19712
rect 19984 19660 20036 19712
rect 20260 19660 20312 19712
rect 22652 19703 22704 19712
rect 22652 19669 22661 19703
rect 22661 19669 22695 19703
rect 22695 19669 22704 19703
rect 22652 19660 22704 19669
rect 25044 19660 25096 19712
rect 25320 19703 25372 19712
rect 25320 19669 25329 19703
rect 25329 19669 25363 19703
rect 25363 19669 25372 19703
rect 25320 19660 25372 19669
rect 27804 19728 27856 19780
rect 30104 19796 30156 19848
rect 31576 19796 31628 19848
rect 26700 19660 26752 19712
rect 27068 19660 27120 19712
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27252 19660 27304 19669
rect 27620 19660 27672 19712
rect 31944 19728 31996 19780
rect 29184 19660 29236 19712
rect 29552 19660 29604 19712
rect 29736 19703 29788 19712
rect 29736 19669 29745 19703
rect 29745 19669 29779 19703
rect 29779 19669 29788 19703
rect 29736 19660 29788 19669
rect 30104 19703 30156 19712
rect 30104 19669 30113 19703
rect 30113 19669 30147 19703
rect 30147 19669 30156 19703
rect 30104 19660 30156 19669
rect 31300 19703 31352 19712
rect 31300 19669 31309 19703
rect 31309 19669 31343 19703
rect 31343 19669 31352 19703
rect 31300 19660 31352 19669
rect 32128 19703 32180 19712
rect 32128 19669 32137 19703
rect 32137 19669 32171 19703
rect 32171 19669 32180 19703
rect 32128 19660 32180 19669
rect 43444 19932 43496 19984
rect 33784 19839 33836 19848
rect 33784 19805 33793 19839
rect 33793 19805 33827 19839
rect 33827 19805 33836 19839
rect 33784 19796 33836 19805
rect 35072 19907 35124 19916
rect 35072 19873 35081 19907
rect 35081 19873 35115 19907
rect 35115 19873 35124 19907
rect 35072 19864 35124 19873
rect 36728 19907 36780 19916
rect 36728 19873 36737 19907
rect 36737 19873 36771 19907
rect 36771 19873 36780 19907
rect 36728 19864 36780 19873
rect 38384 19864 38436 19916
rect 39396 19864 39448 19916
rect 40500 19864 40552 19916
rect 35164 19796 35216 19848
rect 37832 19796 37884 19848
rect 38200 19839 38252 19848
rect 38200 19805 38209 19839
rect 38209 19805 38243 19839
rect 38243 19805 38252 19839
rect 38200 19796 38252 19805
rect 40224 19796 40276 19848
rect 40408 19839 40460 19848
rect 40408 19805 40417 19839
rect 40417 19805 40451 19839
rect 40451 19805 40460 19839
rect 40408 19796 40460 19805
rect 42708 19796 42760 19848
rect 34244 19728 34296 19780
rect 36268 19728 36320 19780
rect 40040 19728 40092 19780
rect 49332 19728 49384 19780
rect 33600 19660 33652 19712
rect 34336 19660 34388 19712
rect 35348 19660 35400 19712
rect 35808 19660 35860 19712
rect 35900 19660 35952 19712
rect 36544 19703 36596 19712
rect 36544 19669 36553 19703
rect 36553 19669 36587 19703
rect 36587 19669 36596 19703
rect 36544 19660 36596 19669
rect 37556 19703 37608 19712
rect 37556 19669 37565 19703
rect 37565 19669 37599 19703
rect 37599 19669 37608 19703
rect 37556 19660 37608 19669
rect 38476 19660 38528 19712
rect 39580 19703 39632 19712
rect 39580 19669 39589 19703
rect 39589 19669 39623 19703
rect 39623 19669 39632 19703
rect 39580 19660 39632 19669
rect 40868 19660 40920 19712
rect 49148 19703 49200 19712
rect 49148 19669 49157 19703
rect 49157 19669 49191 19703
rect 49191 19669 49200 19703
rect 49148 19660 49200 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 7288 19456 7340 19508
rect 7748 19456 7800 19508
rect 13452 19456 13504 19508
rect 3424 19388 3476 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 9220 19388 9272 19440
rect 12808 19388 12860 19440
rect 15016 19456 15068 19508
rect 15936 19456 15988 19508
rect 17316 19456 17368 19508
rect 19892 19456 19944 19508
rect 23940 19456 23992 19508
rect 24308 19456 24360 19508
rect 25228 19456 25280 19508
rect 26056 19456 26108 19508
rect 3884 19252 3936 19304
rect 5816 19320 5868 19372
rect 9588 19320 9640 19372
rect 6828 19252 6880 19304
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 11612 19320 11664 19372
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 12440 19320 12492 19372
rect 12900 19320 12952 19372
rect 16028 19388 16080 19440
rect 16948 19388 17000 19440
rect 17500 19388 17552 19440
rect 19708 19388 19760 19440
rect 20352 19388 20404 19440
rect 23480 19388 23532 19440
rect 24216 19388 24268 19440
rect 26516 19388 26568 19440
rect 12256 19184 12308 19236
rect 15200 19320 15252 19372
rect 15292 19252 15344 19304
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 17040 19320 17092 19372
rect 17592 19320 17644 19372
rect 22560 19320 22612 19372
rect 22652 19320 22704 19372
rect 23296 19320 23348 19372
rect 25688 19320 25740 19372
rect 28356 19456 28408 19508
rect 28724 19456 28776 19508
rect 28816 19456 28868 19508
rect 31392 19456 31444 19508
rect 31668 19456 31720 19508
rect 32864 19456 32916 19508
rect 26700 19388 26752 19440
rect 29644 19388 29696 19440
rect 31484 19431 31536 19440
rect 31484 19397 31493 19431
rect 31493 19397 31527 19431
rect 31527 19397 31536 19431
rect 31484 19388 31536 19397
rect 32496 19388 32548 19440
rect 34520 19456 34572 19508
rect 34888 19456 34940 19508
rect 36544 19456 36596 19508
rect 36912 19456 36964 19508
rect 37372 19456 37424 19508
rect 37924 19456 37976 19508
rect 33968 19388 34020 19440
rect 39580 19456 39632 19508
rect 40040 19456 40092 19508
rect 41052 19456 41104 19508
rect 39488 19388 39540 19440
rect 15568 19252 15620 19304
rect 16120 19252 16172 19304
rect 18604 19252 18656 19304
rect 19800 19295 19852 19304
rect 19800 19261 19809 19295
rect 19809 19261 19843 19295
rect 19843 19261 19852 19295
rect 19800 19252 19852 19261
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 8300 19116 8352 19168
rect 11888 19116 11940 19168
rect 12716 19159 12768 19168
rect 12716 19125 12725 19159
rect 12725 19125 12759 19159
rect 12759 19125 12768 19159
rect 12716 19116 12768 19125
rect 15936 19184 15988 19236
rect 14464 19116 14516 19168
rect 15292 19116 15344 19168
rect 19616 19116 19668 19168
rect 20904 19252 20956 19304
rect 20628 19184 20680 19236
rect 21548 19184 21600 19236
rect 20444 19116 20496 19168
rect 22192 19295 22244 19304
rect 22192 19261 22201 19295
rect 22201 19261 22235 19295
rect 22235 19261 22244 19295
rect 22192 19252 22244 19261
rect 24860 19252 24912 19304
rect 26976 19320 27028 19372
rect 27252 19320 27304 19372
rect 28172 19320 28224 19372
rect 28448 19320 28500 19372
rect 22652 19184 22704 19236
rect 23848 19116 23900 19168
rect 25872 19184 25924 19236
rect 27988 19252 28040 19304
rect 28356 19252 28408 19304
rect 29000 19295 29052 19304
rect 29000 19261 29009 19295
rect 29009 19261 29043 19295
rect 29043 19261 29052 19295
rect 29000 19252 29052 19261
rect 29092 19252 29144 19304
rect 30380 19320 30432 19372
rect 32588 19363 32640 19372
rect 32588 19329 32597 19363
rect 32597 19329 32631 19363
rect 32631 19329 32640 19363
rect 32588 19320 32640 19329
rect 34152 19320 34204 19372
rect 30472 19252 30524 19304
rect 32496 19295 32548 19304
rect 32496 19261 32505 19295
rect 32505 19261 32539 19295
rect 32539 19261 32548 19295
rect 32496 19252 32548 19261
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 28540 19184 28592 19236
rect 31024 19184 31076 19236
rect 34244 19227 34296 19236
rect 34244 19193 34253 19227
rect 34253 19193 34287 19227
rect 34287 19193 34296 19227
rect 34244 19184 34296 19193
rect 34980 19295 35032 19304
rect 34980 19261 34989 19295
rect 34989 19261 35023 19295
rect 35023 19261 35032 19295
rect 34980 19252 35032 19261
rect 35992 19295 36044 19304
rect 35992 19261 36001 19295
rect 36001 19261 36035 19295
rect 36035 19261 36044 19295
rect 35992 19252 36044 19261
rect 36268 19363 36320 19372
rect 36268 19329 36277 19363
rect 36277 19329 36311 19363
rect 36311 19329 36320 19363
rect 36268 19320 36320 19329
rect 48412 19388 48464 19440
rect 49240 19363 49292 19372
rect 49240 19329 49249 19363
rect 49249 19329 49283 19363
rect 49283 19329 49292 19363
rect 49240 19320 49292 19329
rect 37280 19252 37332 19304
rect 39396 19295 39448 19304
rect 39396 19261 39405 19295
rect 39405 19261 39439 19295
rect 39439 19261 39448 19295
rect 39396 19252 39448 19261
rect 37372 19184 37424 19236
rect 37740 19184 37792 19236
rect 29276 19116 29328 19168
rect 30104 19116 30156 19168
rect 30380 19159 30432 19168
rect 30380 19125 30389 19159
rect 30389 19125 30423 19159
rect 30423 19125 30432 19159
rect 30380 19116 30432 19125
rect 33968 19116 34020 19168
rect 35072 19116 35124 19168
rect 36636 19159 36688 19168
rect 36636 19125 36645 19159
rect 36645 19125 36679 19159
rect 36679 19125 36688 19159
rect 36636 19116 36688 19125
rect 36912 19159 36964 19168
rect 36912 19125 36921 19159
rect 36921 19125 36955 19159
rect 36955 19125 36964 19159
rect 36912 19116 36964 19125
rect 37832 19116 37884 19168
rect 41052 19252 41104 19304
rect 42064 19252 42116 19304
rect 40224 19184 40276 19236
rect 40040 19116 40092 19168
rect 41052 19116 41104 19168
rect 49424 19116 49476 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 6828 18912 6880 18964
rect 10968 18912 11020 18964
rect 11060 18912 11112 18964
rect 3516 18776 3568 18828
rect 11152 18844 11204 18896
rect 11888 18955 11940 18964
rect 11888 18921 11897 18955
rect 11897 18921 11931 18955
rect 11931 18921 11940 18955
rect 11888 18912 11940 18921
rect 12532 18844 12584 18896
rect 12716 18844 12768 18896
rect 13360 18844 13412 18896
rect 13636 18887 13688 18896
rect 13636 18853 13645 18887
rect 13645 18853 13679 18887
rect 13679 18853 13688 18887
rect 13636 18844 13688 18853
rect 1400 18640 1452 18692
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 13176 18776 13228 18828
rect 15936 18912 15988 18964
rect 16120 18912 16172 18964
rect 16672 18912 16724 18964
rect 16764 18912 16816 18964
rect 18328 18912 18380 18964
rect 19892 18955 19944 18964
rect 19892 18921 19901 18955
rect 19901 18921 19935 18955
rect 19935 18921 19944 18955
rect 19892 18912 19944 18921
rect 20996 18912 21048 18964
rect 22468 18912 22520 18964
rect 27160 18912 27212 18964
rect 29092 18912 29144 18964
rect 30288 18912 30340 18964
rect 30656 18912 30708 18964
rect 16304 18844 16356 18896
rect 16580 18844 16632 18896
rect 20812 18844 20864 18896
rect 19432 18776 19484 18828
rect 20168 18776 20220 18828
rect 21180 18776 21232 18828
rect 22100 18776 22152 18828
rect 25044 18819 25096 18828
rect 25044 18785 25053 18819
rect 25053 18785 25087 18819
rect 25087 18785 25096 18819
rect 25044 18776 25096 18785
rect 25688 18776 25740 18828
rect 27988 18844 28040 18896
rect 28908 18844 28960 18896
rect 29000 18887 29052 18896
rect 29000 18853 29009 18887
rect 29009 18853 29043 18887
rect 29043 18853 29052 18887
rect 29000 18844 29052 18853
rect 27528 18776 27580 18828
rect 27712 18776 27764 18828
rect 30104 18844 30156 18896
rect 30932 18887 30984 18896
rect 30932 18853 30941 18887
rect 30941 18853 30975 18887
rect 30975 18853 30984 18887
rect 30932 18844 30984 18853
rect 36084 18912 36136 18964
rect 39396 18912 39448 18964
rect 42064 18955 42116 18964
rect 42064 18921 42073 18955
rect 42073 18921 42107 18955
rect 42107 18921 42116 18955
rect 42064 18912 42116 18921
rect 33600 18844 33652 18896
rect 34244 18844 34296 18896
rect 34520 18887 34572 18896
rect 34520 18853 34529 18887
rect 34529 18853 34563 18887
rect 34563 18853 34572 18887
rect 34520 18844 34572 18853
rect 37188 18844 37240 18896
rect 37740 18844 37792 18896
rect 38016 18887 38068 18896
rect 38016 18853 38025 18887
rect 38025 18853 38059 18887
rect 38059 18853 38068 18887
rect 38016 18844 38068 18853
rect 42708 18844 42760 18896
rect 29552 18776 29604 18828
rect 29920 18776 29972 18828
rect 30656 18776 30708 18828
rect 4344 18640 4396 18692
rect 10232 18640 10284 18692
rect 7840 18572 7892 18624
rect 10692 18683 10744 18692
rect 10692 18649 10701 18683
rect 10701 18649 10735 18683
rect 10735 18649 10744 18683
rect 10692 18640 10744 18649
rect 11980 18572 12032 18624
rect 12348 18572 12400 18624
rect 13452 18708 13504 18760
rect 15660 18708 15712 18760
rect 16672 18708 16724 18760
rect 18512 18708 18564 18760
rect 22008 18708 22060 18760
rect 24124 18708 24176 18760
rect 28816 18708 28868 18760
rect 12808 18640 12860 18692
rect 13268 18572 13320 18624
rect 13912 18615 13964 18624
rect 13912 18581 13921 18615
rect 13921 18581 13955 18615
rect 13955 18581 13964 18615
rect 13912 18572 13964 18581
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 14556 18640 14608 18649
rect 17408 18683 17460 18692
rect 17408 18649 17417 18683
rect 17417 18649 17451 18683
rect 17451 18649 17460 18683
rect 17408 18640 17460 18649
rect 19340 18683 19392 18692
rect 19340 18649 19349 18683
rect 19349 18649 19383 18683
rect 19383 18649 19392 18683
rect 19340 18640 19392 18649
rect 15568 18572 15620 18624
rect 16764 18572 16816 18624
rect 18420 18572 18472 18624
rect 18604 18572 18656 18624
rect 19524 18572 19576 18624
rect 19616 18615 19668 18624
rect 19616 18581 19625 18615
rect 19625 18581 19659 18615
rect 19659 18581 19668 18615
rect 19616 18572 19668 18581
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 21916 18572 21968 18624
rect 22744 18640 22796 18692
rect 23480 18640 23532 18692
rect 23848 18640 23900 18692
rect 27436 18640 27488 18692
rect 27528 18640 27580 18692
rect 29460 18708 29512 18760
rect 32772 18819 32824 18828
rect 32772 18785 32781 18819
rect 32781 18785 32815 18819
rect 32815 18785 32824 18819
rect 32772 18776 32824 18785
rect 32956 18819 33008 18828
rect 32956 18785 32965 18819
rect 32965 18785 32999 18819
rect 32999 18785 33008 18819
rect 32956 18776 33008 18785
rect 33048 18776 33100 18828
rect 34060 18776 34112 18828
rect 37096 18776 37148 18828
rect 37924 18776 37976 18828
rect 38568 18819 38620 18828
rect 38568 18785 38577 18819
rect 38577 18785 38611 18819
rect 38611 18785 38620 18819
rect 38568 18776 38620 18785
rect 35348 18708 35400 18760
rect 24768 18572 24820 18624
rect 26792 18572 26844 18624
rect 27988 18572 28040 18624
rect 28172 18572 28224 18624
rect 28448 18572 28500 18624
rect 35532 18640 35584 18692
rect 37648 18708 37700 18760
rect 40040 18708 40092 18760
rect 48780 18708 48832 18760
rect 49424 18708 49476 18760
rect 29368 18572 29420 18624
rect 30472 18615 30524 18624
rect 30472 18581 30481 18615
rect 30481 18581 30515 18615
rect 30515 18581 30524 18615
rect 30472 18572 30524 18581
rect 30656 18572 30708 18624
rect 30932 18572 30984 18624
rect 31392 18572 31444 18624
rect 31668 18572 31720 18624
rect 31944 18615 31996 18624
rect 31944 18581 31953 18615
rect 31953 18581 31987 18615
rect 31987 18581 31996 18615
rect 31944 18572 31996 18581
rect 32036 18572 32088 18624
rect 34152 18572 34204 18624
rect 36268 18572 36320 18624
rect 37556 18572 37608 18624
rect 39764 18640 39816 18692
rect 39948 18572 40000 18624
rect 40132 18572 40184 18624
rect 40224 18572 40276 18624
rect 48412 18615 48464 18624
rect 48412 18581 48421 18615
rect 48421 18581 48455 18615
rect 48455 18581 48464 18615
rect 48412 18572 48464 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 4160 18300 4212 18352
rect 5632 18300 5684 18352
rect 9864 18368 9916 18420
rect 11796 18368 11848 18420
rect 10048 18300 10100 18352
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 4068 18232 4120 18284
rect 11244 18300 11296 18352
rect 12440 18300 12492 18352
rect 13176 18343 13228 18352
rect 13176 18309 13185 18343
rect 13185 18309 13219 18343
rect 13219 18309 13228 18343
rect 13176 18300 13228 18309
rect 13268 18300 13320 18352
rect 23296 18368 23348 18420
rect 4252 18164 4304 18216
rect 6828 18096 6880 18148
rect 11796 18232 11848 18284
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 13820 18232 13872 18284
rect 14188 18232 14240 18284
rect 18512 18300 18564 18352
rect 18236 18232 18288 18284
rect 10600 18164 10652 18216
rect 11704 18164 11756 18216
rect 12532 18164 12584 18216
rect 9772 18028 9824 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 14556 18207 14608 18216
rect 14556 18173 14565 18207
rect 14565 18173 14599 18207
rect 14599 18173 14608 18207
rect 14556 18164 14608 18173
rect 16488 18164 16540 18216
rect 16672 18207 16724 18216
rect 16672 18173 16681 18207
rect 16681 18173 16715 18207
rect 16715 18173 16724 18207
rect 16672 18164 16724 18173
rect 17500 18164 17552 18216
rect 13636 18028 13688 18080
rect 15108 18028 15160 18080
rect 15752 18096 15804 18148
rect 16304 18096 16356 18148
rect 18328 18096 18380 18148
rect 16580 18028 16632 18080
rect 19156 18300 19208 18352
rect 19984 18300 20036 18352
rect 21456 18300 21508 18352
rect 21732 18300 21784 18352
rect 25780 18368 25832 18420
rect 27252 18368 27304 18420
rect 27528 18411 27580 18420
rect 27528 18377 27537 18411
rect 27537 18377 27571 18411
rect 27571 18377 27580 18411
rect 27528 18368 27580 18377
rect 27712 18368 27764 18420
rect 29736 18368 29788 18420
rect 29828 18368 29880 18420
rect 31208 18368 31260 18420
rect 32312 18368 32364 18420
rect 32956 18368 33008 18420
rect 24124 18343 24176 18352
rect 24124 18309 24133 18343
rect 24133 18309 24167 18343
rect 24167 18309 24176 18343
rect 24124 18300 24176 18309
rect 19616 18207 19668 18216
rect 19616 18173 19625 18207
rect 19625 18173 19659 18207
rect 19659 18173 19668 18207
rect 19616 18164 19668 18173
rect 20352 18164 20404 18216
rect 22468 18164 22520 18216
rect 23296 18275 23348 18284
rect 23296 18241 23305 18275
rect 23305 18241 23339 18275
rect 23339 18241 23348 18275
rect 23296 18232 23348 18241
rect 32128 18300 32180 18352
rect 35348 18411 35400 18420
rect 35348 18377 35357 18411
rect 35357 18377 35391 18411
rect 35391 18377 35400 18411
rect 35348 18368 35400 18377
rect 35532 18368 35584 18420
rect 36820 18368 36872 18420
rect 37556 18368 37608 18420
rect 37740 18368 37792 18420
rect 40868 18411 40920 18420
rect 40868 18377 40877 18411
rect 40877 18377 40911 18411
rect 40911 18377 40920 18411
rect 40868 18368 40920 18377
rect 48780 18411 48832 18420
rect 48780 18377 48789 18411
rect 48789 18377 48823 18411
rect 48823 18377 48832 18411
rect 48780 18368 48832 18377
rect 36176 18300 36228 18352
rect 37464 18300 37516 18352
rect 38016 18300 38068 18352
rect 48412 18300 48464 18352
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 19432 18096 19484 18148
rect 21364 18071 21416 18080
rect 21364 18037 21373 18071
rect 21373 18037 21407 18071
rect 21407 18037 21416 18071
rect 21364 18028 21416 18037
rect 21456 18028 21508 18080
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 26424 18207 26476 18216
rect 26424 18173 26433 18207
rect 26433 18173 26467 18207
rect 26467 18173 26476 18207
rect 26424 18164 26476 18173
rect 27528 18232 27580 18284
rect 27712 18207 27764 18216
rect 27712 18173 27721 18207
rect 27721 18173 27755 18207
rect 27755 18173 27764 18207
rect 27712 18164 27764 18173
rect 23756 18096 23808 18148
rect 22836 18028 22888 18080
rect 25044 18028 25096 18080
rect 26056 18096 26108 18148
rect 27068 18028 27120 18080
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 27620 18028 27672 18080
rect 29736 18071 29788 18080
rect 29736 18037 29745 18071
rect 29745 18037 29779 18071
rect 29779 18037 29788 18071
rect 29736 18028 29788 18037
rect 33324 18232 33376 18284
rect 30564 18164 30616 18216
rect 30932 18164 30984 18216
rect 32404 18207 32456 18216
rect 32404 18173 32413 18207
rect 32413 18173 32447 18207
rect 32447 18173 32456 18207
rect 32404 18164 32456 18173
rect 30748 18028 30800 18080
rect 31024 18096 31076 18148
rect 33600 18207 33652 18216
rect 33600 18173 33609 18207
rect 33609 18173 33643 18207
rect 33643 18173 33652 18207
rect 33600 18164 33652 18173
rect 34520 18164 34572 18216
rect 36268 18275 36320 18284
rect 36268 18241 36277 18275
rect 36277 18241 36311 18275
rect 36311 18241 36320 18275
rect 36268 18232 36320 18241
rect 37188 18232 37240 18284
rect 37924 18232 37976 18284
rect 39764 18275 39816 18284
rect 39764 18241 39773 18275
rect 39773 18241 39807 18275
rect 39807 18241 39816 18275
rect 39764 18232 39816 18241
rect 49332 18275 49384 18284
rect 49332 18241 49341 18275
rect 49341 18241 49375 18275
rect 49375 18241 49384 18275
rect 49332 18232 49384 18241
rect 37740 18164 37792 18216
rect 37832 18164 37884 18216
rect 35716 18096 35768 18148
rect 36728 18096 36780 18148
rect 33692 18028 33744 18080
rect 34980 18028 35032 18080
rect 36544 18028 36596 18080
rect 37096 18096 37148 18148
rect 37924 18096 37976 18148
rect 38016 18139 38068 18148
rect 38016 18105 38025 18139
rect 38025 18105 38059 18139
rect 38059 18105 38068 18139
rect 38016 18096 38068 18105
rect 37004 18028 37056 18080
rect 37280 18028 37332 18080
rect 37464 18028 37516 18080
rect 40224 18096 40276 18148
rect 40040 18071 40092 18080
rect 40040 18037 40049 18071
rect 40049 18037 40083 18071
rect 40083 18037 40092 18071
rect 40040 18028 40092 18037
rect 49148 18071 49200 18080
rect 49148 18037 49157 18071
rect 49157 18037 49191 18071
rect 49191 18037 49200 18071
rect 49148 18028 49200 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 10232 17824 10284 17876
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 13544 17824 13596 17876
rect 14556 17824 14608 17876
rect 11428 17688 11480 17740
rect 12532 17688 12584 17740
rect 13452 17688 13504 17740
rect 16672 17824 16724 17876
rect 17224 17824 17276 17876
rect 19340 17824 19392 17876
rect 19616 17824 19668 17876
rect 10416 17620 10468 17672
rect 15384 17688 15436 17740
rect 16028 17731 16080 17740
rect 16028 17697 16037 17731
rect 16037 17697 16071 17731
rect 16071 17697 16080 17731
rect 16028 17688 16080 17697
rect 16304 17688 16356 17740
rect 19984 17756 20036 17808
rect 16856 17731 16908 17740
rect 16856 17697 16865 17731
rect 16865 17697 16899 17731
rect 16899 17697 16908 17731
rect 16856 17688 16908 17697
rect 18328 17688 18380 17740
rect 21088 17824 21140 17876
rect 21180 17824 21232 17876
rect 22284 17824 22336 17876
rect 22560 17824 22612 17876
rect 23572 17824 23624 17876
rect 26240 17867 26292 17876
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 22100 17756 22152 17808
rect 25228 17756 25280 17808
rect 28816 17824 28868 17876
rect 29644 17867 29696 17876
rect 29644 17833 29653 17867
rect 29653 17833 29687 17867
rect 29687 17833 29696 17867
rect 29644 17824 29696 17833
rect 31484 17824 31536 17876
rect 30012 17756 30064 17808
rect 20260 17688 20312 17740
rect 21180 17688 21232 17740
rect 21640 17688 21692 17740
rect 22192 17688 22244 17740
rect 24860 17688 24912 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 1032 17552 1084 17604
rect 11980 17552 12032 17604
rect 12072 17595 12124 17604
rect 12072 17561 12081 17595
rect 12081 17561 12115 17595
rect 12115 17561 12124 17595
rect 12072 17552 12124 17561
rect 11704 17484 11756 17536
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 16488 17620 16540 17672
rect 18880 17620 18932 17672
rect 15292 17552 15344 17604
rect 15660 17552 15712 17604
rect 20352 17552 20404 17604
rect 15936 17484 15988 17536
rect 16304 17484 16356 17536
rect 16488 17527 16540 17536
rect 16488 17493 16497 17527
rect 16497 17493 16531 17527
rect 16531 17493 16540 17527
rect 16488 17484 16540 17493
rect 17408 17484 17460 17536
rect 18604 17484 18656 17536
rect 20260 17527 20312 17536
rect 20260 17493 20269 17527
rect 20269 17493 20303 17527
rect 20303 17493 20312 17527
rect 20260 17484 20312 17493
rect 23480 17620 23532 17672
rect 28448 17688 28500 17740
rect 29092 17688 29144 17740
rect 29920 17688 29972 17740
rect 30288 17688 30340 17740
rect 31116 17688 31168 17740
rect 31484 17731 31536 17740
rect 31484 17697 31493 17731
rect 31493 17697 31527 17731
rect 31527 17697 31536 17731
rect 31484 17688 31536 17697
rect 38384 17824 38436 17876
rect 39948 17824 40000 17876
rect 40592 17824 40644 17876
rect 49148 17824 49200 17876
rect 33968 17756 34020 17808
rect 34244 17756 34296 17808
rect 34980 17756 35032 17808
rect 40868 17756 40920 17808
rect 33232 17688 33284 17740
rect 34520 17688 34572 17740
rect 35716 17688 35768 17740
rect 37280 17688 37332 17740
rect 40040 17688 40092 17740
rect 40684 17688 40736 17740
rect 27436 17620 27488 17672
rect 28908 17620 28960 17672
rect 31760 17620 31812 17672
rect 20996 17552 21048 17604
rect 21732 17552 21784 17604
rect 24768 17552 24820 17604
rect 27252 17552 27304 17604
rect 22100 17484 22152 17536
rect 23756 17527 23808 17536
rect 23756 17493 23765 17527
rect 23765 17493 23799 17527
rect 23799 17493 23808 17527
rect 23756 17484 23808 17493
rect 24860 17484 24912 17536
rect 27620 17484 27672 17536
rect 28816 17484 28868 17536
rect 30012 17552 30064 17604
rect 30748 17595 30800 17604
rect 30748 17561 30757 17595
rect 30757 17561 30791 17595
rect 30791 17561 30800 17595
rect 30748 17552 30800 17561
rect 37556 17663 37608 17672
rect 37556 17629 37565 17663
rect 37565 17629 37599 17663
rect 37599 17629 37608 17663
rect 37556 17620 37608 17629
rect 37924 17620 37976 17672
rect 38660 17620 38712 17672
rect 38844 17620 38896 17672
rect 49332 17663 49384 17672
rect 49332 17629 49341 17663
rect 49341 17629 49375 17663
rect 49375 17629 49384 17663
rect 49332 17620 49384 17629
rect 31944 17484 31996 17536
rect 32312 17527 32364 17536
rect 32312 17493 32321 17527
rect 32321 17493 32355 17527
rect 32355 17493 32364 17527
rect 32312 17484 32364 17493
rect 33416 17484 33468 17536
rect 35992 17552 36044 17604
rect 36544 17552 36596 17604
rect 37004 17552 37056 17604
rect 37372 17552 37424 17604
rect 48412 17552 48464 17604
rect 49240 17552 49292 17604
rect 35072 17527 35124 17536
rect 35072 17493 35081 17527
rect 35081 17493 35115 17527
rect 35115 17493 35124 17527
rect 35072 17484 35124 17493
rect 35532 17484 35584 17536
rect 36636 17484 36688 17536
rect 38936 17484 38988 17536
rect 49148 17527 49200 17536
rect 49148 17493 49157 17527
rect 49157 17493 49191 17527
rect 49191 17493 49200 17527
rect 49148 17484 49200 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 7840 17280 7892 17332
rect 13360 17280 13412 17332
rect 14004 17280 14056 17332
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 3332 17212 3384 17264
rect 4344 17144 4396 17196
rect 9496 17144 9548 17196
rect 10508 17144 10560 17196
rect 10784 17187 10836 17196
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 10784 17144 10836 17153
rect 11428 17212 11480 17264
rect 11888 17255 11940 17264
rect 11888 17221 11897 17255
rect 11897 17221 11931 17255
rect 11931 17221 11940 17255
rect 11888 17212 11940 17221
rect 12164 17212 12216 17264
rect 13912 17212 13964 17264
rect 14740 17212 14792 17264
rect 15752 17212 15804 17264
rect 16028 17212 16080 17264
rect 17960 17255 18012 17264
rect 17960 17221 17969 17255
rect 17969 17221 18003 17255
rect 18003 17221 18012 17255
rect 17960 17212 18012 17221
rect 19156 17323 19208 17332
rect 19156 17289 19165 17323
rect 19165 17289 19199 17323
rect 19199 17289 19208 17323
rect 19156 17280 19208 17289
rect 19708 17280 19760 17332
rect 20904 17280 20956 17332
rect 23480 17280 23532 17332
rect 24952 17280 25004 17332
rect 27712 17323 27764 17332
rect 27712 17289 27721 17323
rect 27721 17289 27755 17323
rect 27755 17289 27764 17323
rect 27712 17280 27764 17289
rect 27804 17280 27856 17332
rect 29276 17280 29328 17332
rect 20996 17212 21048 17264
rect 21456 17212 21508 17264
rect 21548 17212 21600 17264
rect 22836 17212 22888 17264
rect 24124 17212 24176 17264
rect 940 17076 992 17128
rect 5816 17076 5868 17128
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 12808 17119 12860 17128
rect 12808 17085 12817 17119
rect 12817 17085 12851 17119
rect 12851 17085 12860 17119
rect 12808 17076 12860 17085
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 15200 17144 15252 17196
rect 14648 17076 14700 17128
rect 16948 17144 17000 17196
rect 12624 17008 12676 17060
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 18880 17144 18932 17196
rect 22192 17144 22244 17196
rect 22744 17144 22796 17196
rect 25964 17255 26016 17264
rect 25964 17221 25973 17255
rect 25973 17221 26007 17255
rect 26007 17221 26016 17255
rect 25964 17212 26016 17221
rect 29644 17212 29696 17264
rect 30932 17280 30984 17332
rect 31576 17280 31628 17332
rect 30656 17212 30708 17264
rect 30748 17212 30800 17264
rect 33600 17280 33652 17332
rect 34060 17323 34112 17332
rect 34060 17289 34069 17323
rect 34069 17289 34103 17323
rect 34103 17289 34112 17323
rect 34060 17280 34112 17289
rect 35072 17280 35124 17332
rect 25596 17144 25648 17196
rect 19892 17076 19944 17128
rect 19984 17076 20036 17128
rect 21824 17076 21876 17128
rect 22008 17119 22060 17128
rect 22008 17085 22017 17119
rect 22017 17085 22051 17119
rect 22051 17085 22060 17119
rect 22008 17076 22060 17085
rect 25504 17119 25556 17128
rect 25504 17085 25513 17119
rect 25513 17085 25547 17119
rect 25547 17085 25556 17119
rect 25504 17076 25556 17085
rect 16488 17008 16540 17060
rect 12164 16940 12216 16992
rect 12440 16983 12492 16992
rect 12440 16949 12449 16983
rect 12449 16949 12483 16983
rect 12483 16949 12492 16983
rect 12440 16940 12492 16949
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 14096 16940 14148 16992
rect 16764 16940 16816 16992
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 20904 16940 20956 16992
rect 21548 16983 21600 16992
rect 21548 16949 21557 16983
rect 21557 16949 21591 16983
rect 21591 16949 21600 16983
rect 21548 16940 21600 16949
rect 24584 17008 24636 17060
rect 26424 17144 26476 17196
rect 27068 17144 27120 17196
rect 27804 17119 27856 17128
rect 27804 17085 27813 17119
rect 27813 17085 27847 17119
rect 27847 17085 27856 17119
rect 27804 17076 27856 17085
rect 28264 17144 28316 17196
rect 29184 17144 29236 17196
rect 26884 17008 26936 17060
rect 29920 17119 29972 17128
rect 29920 17085 29929 17119
rect 29929 17085 29963 17119
rect 29963 17085 29972 17119
rect 29920 17076 29972 17085
rect 30748 17076 30800 17128
rect 32220 17144 32272 17196
rect 33876 17212 33928 17264
rect 34980 17212 35032 17264
rect 35532 17255 35584 17264
rect 35532 17221 35541 17255
rect 35541 17221 35575 17255
rect 35575 17221 35584 17255
rect 35532 17212 35584 17221
rect 40592 17280 40644 17332
rect 48412 17323 48464 17332
rect 48412 17289 48421 17323
rect 48421 17289 48455 17323
rect 48455 17289 48464 17323
rect 48412 17280 48464 17289
rect 35624 17144 35676 17196
rect 36360 17187 36412 17196
rect 36360 17153 36369 17187
rect 36369 17153 36403 17187
rect 36403 17153 36412 17187
rect 36360 17144 36412 17153
rect 32588 17119 32640 17128
rect 32588 17085 32597 17119
rect 32597 17085 32631 17119
rect 32631 17085 32640 17119
rect 32588 17076 32640 17085
rect 34796 17119 34848 17128
rect 34796 17085 34805 17119
rect 34805 17085 34839 17119
rect 34839 17085 34848 17119
rect 34796 17076 34848 17085
rect 36176 17119 36228 17128
rect 36176 17085 36185 17119
rect 36185 17085 36219 17119
rect 36219 17085 36228 17119
rect 36176 17076 36228 17085
rect 38660 17212 38712 17264
rect 40132 17212 40184 17264
rect 38936 17144 38988 17196
rect 48780 17144 48832 17196
rect 49332 17144 49384 17196
rect 32128 17008 32180 17060
rect 32312 17008 32364 17060
rect 35440 17008 35492 17060
rect 37832 17076 37884 17128
rect 38384 17076 38436 17128
rect 36452 17008 36504 17060
rect 40684 17119 40736 17128
rect 40684 17085 40693 17119
rect 40693 17085 40727 17119
rect 40727 17085 40736 17119
rect 40684 17076 40736 17085
rect 49056 17119 49108 17128
rect 49056 17085 49065 17119
rect 49065 17085 49099 17119
rect 49099 17085 49108 17119
rect 49056 17076 49108 17085
rect 43904 17008 43956 17060
rect 26240 16940 26292 16992
rect 27988 16940 28040 16992
rect 28632 16940 28684 16992
rect 31300 16940 31352 16992
rect 31760 16983 31812 16992
rect 31760 16949 31769 16983
rect 31769 16949 31803 16983
rect 31803 16949 31812 16983
rect 31760 16940 31812 16949
rect 31852 16940 31904 16992
rect 35348 16940 35400 16992
rect 36728 16983 36780 16992
rect 36728 16949 36737 16983
rect 36737 16949 36771 16983
rect 36771 16949 36780 16983
rect 36728 16940 36780 16949
rect 38844 16940 38896 16992
rect 40040 16940 40092 16992
rect 41052 16940 41104 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 10324 16668 10376 16720
rect 14832 16736 14884 16788
rect 4436 16600 4488 16652
rect 5448 16600 5500 16652
rect 3332 16532 3384 16584
rect 1032 16464 1084 16516
rect 9036 16600 9088 16652
rect 10968 16600 11020 16652
rect 12440 16600 12492 16652
rect 14280 16668 14332 16720
rect 7748 16532 7800 16584
rect 12256 16532 12308 16584
rect 13820 16532 13872 16584
rect 9680 16464 9732 16516
rect 10508 16507 10560 16516
rect 10508 16473 10517 16507
rect 10517 16473 10551 16507
rect 10551 16473 10560 16507
rect 10508 16464 10560 16473
rect 12808 16464 12860 16516
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 11336 16439 11388 16448
rect 11336 16405 11345 16439
rect 11345 16405 11379 16439
rect 11379 16405 11388 16439
rect 11336 16396 11388 16405
rect 12440 16396 12492 16448
rect 12716 16396 12768 16448
rect 13268 16396 13320 16448
rect 14096 16600 14148 16652
rect 15568 16668 15620 16720
rect 17408 16736 17460 16788
rect 20720 16736 20772 16788
rect 20996 16779 21048 16788
rect 20996 16745 21005 16779
rect 21005 16745 21039 16779
rect 21039 16745 21048 16779
rect 20996 16736 21048 16745
rect 21732 16736 21784 16788
rect 21824 16736 21876 16788
rect 23296 16736 23348 16788
rect 28816 16736 28868 16788
rect 30104 16736 30156 16788
rect 14740 16575 14792 16584
rect 14740 16541 14749 16575
rect 14749 16541 14783 16575
rect 14783 16541 14792 16575
rect 14740 16532 14792 16541
rect 15844 16532 15896 16584
rect 16856 16600 16908 16652
rect 17960 16600 18012 16652
rect 19156 16600 19208 16652
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 17500 16532 17552 16584
rect 16948 16464 17000 16516
rect 14188 16396 14240 16448
rect 15476 16396 15528 16448
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 17132 16439 17184 16448
rect 17132 16405 17141 16439
rect 17141 16405 17175 16439
rect 17175 16405 17184 16439
rect 17132 16396 17184 16405
rect 18604 16507 18656 16516
rect 18604 16473 18613 16507
rect 18613 16473 18647 16507
rect 18647 16473 18656 16507
rect 18604 16464 18656 16473
rect 20904 16532 20956 16584
rect 26056 16668 26108 16720
rect 27344 16668 27396 16720
rect 25228 16532 25280 16584
rect 19064 16396 19116 16448
rect 20904 16396 20956 16448
rect 22560 16464 22612 16516
rect 22836 16396 22888 16448
rect 23296 16439 23348 16448
rect 23296 16405 23305 16439
rect 23305 16405 23339 16439
rect 23339 16405 23348 16439
rect 23296 16396 23348 16405
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 24952 16464 25004 16516
rect 25320 16396 25372 16448
rect 25688 16600 25740 16652
rect 27620 16600 27672 16652
rect 27804 16668 27856 16720
rect 31024 16668 31076 16720
rect 28080 16600 28132 16652
rect 28264 16643 28316 16652
rect 28264 16609 28273 16643
rect 28273 16609 28307 16643
rect 28307 16609 28316 16643
rect 28264 16600 28316 16609
rect 28540 16600 28592 16652
rect 28632 16643 28684 16652
rect 28632 16609 28641 16643
rect 28641 16609 28675 16643
rect 28675 16609 28684 16643
rect 28632 16600 28684 16609
rect 29276 16643 29328 16652
rect 29276 16609 29285 16643
rect 29285 16609 29319 16643
rect 29319 16609 29328 16643
rect 29276 16600 29328 16609
rect 29460 16600 29512 16652
rect 30104 16600 30156 16652
rect 34520 16736 34572 16788
rect 36360 16736 36412 16788
rect 40224 16736 40276 16788
rect 41052 16779 41104 16788
rect 41052 16745 41061 16779
rect 41061 16745 41095 16779
rect 41095 16745 41104 16779
rect 41052 16736 41104 16745
rect 41236 16779 41288 16788
rect 41236 16745 41245 16779
rect 41245 16745 41279 16779
rect 41279 16745 41288 16779
rect 41236 16736 41288 16745
rect 48780 16779 48832 16788
rect 48780 16745 48789 16779
rect 48789 16745 48823 16779
rect 48823 16745 48832 16779
rect 48780 16736 48832 16745
rect 31300 16668 31352 16720
rect 28908 16532 28960 16584
rect 26976 16464 27028 16516
rect 31024 16532 31076 16584
rect 32220 16643 32272 16652
rect 32220 16609 32229 16643
rect 32229 16609 32263 16643
rect 32263 16609 32272 16643
rect 32220 16600 32272 16609
rect 34980 16668 35032 16720
rect 37556 16668 37608 16720
rect 41972 16668 42024 16720
rect 31852 16532 31904 16584
rect 35532 16532 35584 16584
rect 36820 16643 36872 16652
rect 36820 16609 36829 16643
rect 36829 16609 36863 16643
rect 36863 16609 36872 16643
rect 36820 16600 36872 16609
rect 37832 16600 37884 16652
rect 38844 16600 38896 16652
rect 40316 16600 40368 16652
rect 41052 16600 41104 16652
rect 39488 16575 39540 16584
rect 39488 16541 39497 16575
rect 39497 16541 39531 16575
rect 39531 16541 39540 16575
rect 39488 16532 39540 16541
rect 40684 16532 40736 16584
rect 41604 16532 41656 16584
rect 49424 16532 49476 16584
rect 29368 16464 29420 16516
rect 26148 16396 26200 16448
rect 26240 16396 26292 16448
rect 26700 16396 26752 16448
rect 27436 16396 27488 16448
rect 28264 16396 28316 16448
rect 28632 16396 28684 16448
rect 32220 16464 32272 16516
rect 32404 16464 32456 16516
rect 33876 16464 33928 16516
rect 35900 16464 35952 16516
rect 38660 16464 38712 16516
rect 40224 16464 40276 16516
rect 41236 16464 41288 16516
rect 31300 16439 31352 16448
rect 31300 16405 31309 16439
rect 31309 16405 31343 16439
rect 31343 16405 31352 16439
rect 31300 16396 31352 16405
rect 31668 16439 31720 16448
rect 31668 16405 31677 16439
rect 31677 16405 31711 16439
rect 31711 16405 31720 16439
rect 31668 16396 31720 16405
rect 33968 16439 34020 16448
rect 33968 16405 33977 16439
rect 33977 16405 34011 16439
rect 34011 16405 34020 16439
rect 33968 16396 34020 16405
rect 34060 16396 34112 16448
rect 34336 16439 34388 16448
rect 34336 16405 34345 16439
rect 34345 16405 34379 16439
rect 34379 16405 34388 16439
rect 34336 16396 34388 16405
rect 36544 16396 36596 16448
rect 37004 16396 37056 16448
rect 37464 16396 37516 16448
rect 38568 16396 38620 16448
rect 40960 16396 41012 16448
rect 49148 16439 49200 16448
rect 49148 16405 49157 16439
rect 49157 16405 49191 16439
rect 49191 16405 49200 16439
rect 49148 16396 49200 16405
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 11336 16192 11388 16244
rect 10876 16124 10928 16176
rect 11428 16124 11480 16176
rect 14004 16124 14056 16176
rect 15108 16192 15160 16244
rect 16396 16192 16448 16244
rect 18328 16192 18380 16244
rect 19340 16192 19392 16244
rect 16304 16124 16356 16176
rect 16856 16124 16908 16176
rect 17132 16124 17184 16176
rect 4252 16056 4304 16108
rect 1032 15988 1084 16040
rect 9036 15988 9088 16040
rect 11704 16056 11756 16108
rect 13176 16056 13228 16108
rect 13268 16056 13320 16108
rect 10784 15988 10836 16040
rect 10968 15988 11020 16040
rect 13360 15988 13412 16040
rect 9772 15920 9824 15972
rect 13820 15988 13872 16040
rect 15016 16056 15068 16108
rect 17776 16056 17828 16108
rect 14832 15988 14884 16040
rect 15568 15988 15620 16040
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 17132 15988 17184 16040
rect 20904 16124 20956 16176
rect 21548 16124 21600 16176
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 24768 16124 24820 16176
rect 25780 16124 25832 16176
rect 26148 16124 26200 16176
rect 6828 15852 6880 15904
rect 10324 15852 10376 15904
rect 13912 15920 13964 15972
rect 14280 15920 14332 15972
rect 15292 15920 15344 15972
rect 17592 15920 17644 15972
rect 20628 15988 20680 16040
rect 11428 15852 11480 15904
rect 12716 15852 12768 15904
rect 12900 15852 12952 15904
rect 14004 15852 14056 15904
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 16948 15852 17000 15861
rect 17316 15852 17368 15904
rect 18880 15895 18932 15904
rect 18880 15861 18889 15895
rect 18889 15861 18923 15895
rect 18923 15861 18932 15895
rect 18880 15852 18932 15861
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 27804 16124 27856 16176
rect 26700 16099 26752 16108
rect 26700 16065 26709 16099
rect 26709 16065 26743 16099
rect 26743 16065 26752 16099
rect 26700 16056 26752 16065
rect 27344 16056 27396 16108
rect 28908 16124 28960 16176
rect 30656 16192 30708 16244
rect 31760 16192 31812 16244
rect 34796 16192 34848 16244
rect 31668 16124 31720 16176
rect 32036 16124 32088 16176
rect 20904 15963 20956 15972
rect 20904 15929 20913 15963
rect 20913 15929 20947 15963
rect 20947 15929 20956 15963
rect 20904 15920 20956 15929
rect 21364 15920 21416 15972
rect 23388 16031 23440 16040
rect 23388 15997 23397 16031
rect 23397 15997 23431 16031
rect 23431 15997 23440 16031
rect 23388 15988 23440 15997
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 26056 16031 26108 16040
rect 26056 15997 26065 16031
rect 26065 15997 26099 16031
rect 26099 15997 26108 16031
rect 26056 15988 26108 15997
rect 24860 15920 24912 15972
rect 27344 15920 27396 15972
rect 21548 15852 21600 15904
rect 21824 15852 21876 15904
rect 22468 15852 22520 15904
rect 26700 15852 26752 15904
rect 28632 16031 28684 16040
rect 28632 15997 28641 16031
rect 28641 15997 28675 16031
rect 28675 15997 28684 16031
rect 28632 15988 28684 15997
rect 29000 15988 29052 16040
rect 29368 15988 29420 16040
rect 30104 16056 30156 16108
rect 29828 15988 29880 16040
rect 30840 16099 30892 16108
rect 30840 16065 30849 16099
rect 30849 16065 30883 16099
rect 30883 16065 30892 16099
rect 30840 16056 30892 16065
rect 31024 16056 31076 16108
rect 34980 16124 35032 16176
rect 31392 15988 31444 16040
rect 32496 16031 32548 16040
rect 32496 15997 32505 16031
rect 32505 15997 32539 16031
rect 32539 15997 32548 16031
rect 32496 15988 32548 15997
rect 33324 16056 33376 16108
rect 37188 16192 37240 16244
rect 40960 16235 41012 16244
rect 40960 16201 40969 16235
rect 40969 16201 41003 16235
rect 41003 16201 41012 16235
rect 40960 16192 41012 16201
rect 38568 16124 38620 16176
rect 39948 16124 40000 16176
rect 37372 16056 37424 16108
rect 48688 16056 48740 16108
rect 49332 16099 49384 16108
rect 49332 16065 49341 16099
rect 49341 16065 49375 16099
rect 49375 16065 49384 16099
rect 49332 16056 49384 16065
rect 32772 15988 32824 16040
rect 36268 15988 36320 16040
rect 37280 15988 37332 16040
rect 37464 16031 37516 16040
rect 37464 15997 37473 16031
rect 37473 15997 37507 16031
rect 37507 15997 37516 16031
rect 37464 15988 37516 15997
rect 39212 15988 39264 16040
rect 41788 15988 41840 16040
rect 28632 15852 28684 15904
rect 30748 15852 30800 15904
rect 31392 15852 31444 15904
rect 33416 15920 33468 15972
rect 34336 15920 34388 15972
rect 35532 15920 35584 15972
rect 49148 15963 49200 15972
rect 49148 15929 49157 15963
rect 49157 15929 49191 15963
rect 49191 15929 49200 15963
rect 49148 15920 49200 15929
rect 31760 15852 31812 15904
rect 31852 15895 31904 15904
rect 31852 15861 31861 15895
rect 31861 15861 31895 15895
rect 31895 15861 31904 15895
rect 31852 15852 31904 15861
rect 32680 15852 32732 15904
rect 33692 15852 33744 15904
rect 34612 15852 34664 15904
rect 35164 15895 35216 15904
rect 35164 15861 35173 15895
rect 35173 15861 35207 15895
rect 35207 15861 35216 15895
rect 35164 15852 35216 15861
rect 36820 15852 36872 15904
rect 40316 15852 40368 15904
rect 41604 15895 41656 15904
rect 41604 15861 41613 15895
rect 41613 15861 41647 15895
rect 41647 15861 41656 15895
rect 41604 15852 41656 15861
rect 42064 15852 42116 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 10692 15648 10744 15700
rect 10968 15648 11020 15700
rect 12164 15648 12216 15700
rect 16580 15648 16632 15700
rect 17868 15691 17920 15700
rect 17868 15657 17877 15691
rect 17877 15657 17911 15691
rect 17911 15657 17920 15691
rect 17868 15648 17920 15657
rect 18788 15648 18840 15700
rect 18972 15691 19024 15700
rect 18972 15657 18981 15691
rect 18981 15657 19015 15691
rect 19015 15657 19024 15691
rect 18972 15648 19024 15657
rect 19524 15648 19576 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20812 15648 20864 15700
rect 21364 15648 21416 15700
rect 12900 15580 12952 15632
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 15108 15580 15160 15632
rect 15384 15580 15436 15632
rect 15844 15580 15896 15632
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 15568 15512 15620 15564
rect 16120 15555 16172 15564
rect 16120 15521 16129 15555
rect 16129 15521 16163 15555
rect 16163 15521 16172 15555
rect 16120 15512 16172 15521
rect 16396 15512 16448 15564
rect 18420 15623 18472 15632
rect 18420 15589 18429 15623
rect 18429 15589 18463 15623
rect 18463 15589 18472 15623
rect 18420 15580 18472 15589
rect 21916 15580 21968 15632
rect 22468 15623 22520 15632
rect 22468 15589 22477 15623
rect 22477 15589 22511 15623
rect 22511 15589 22520 15623
rect 22468 15580 22520 15589
rect 23848 15580 23900 15632
rect 26056 15648 26108 15700
rect 26792 15648 26844 15700
rect 30196 15648 30248 15700
rect 21364 15512 21416 15564
rect 21456 15512 21508 15564
rect 10232 15444 10284 15496
rect 12624 15444 12676 15496
rect 13452 15444 13504 15496
rect 13728 15444 13780 15496
rect 18420 15444 18472 15496
rect 23296 15512 23348 15564
rect 23940 15512 23992 15564
rect 24032 15512 24084 15564
rect 27528 15580 27580 15632
rect 32588 15580 32640 15632
rect 25320 15512 25372 15564
rect 26608 15512 26660 15564
rect 31116 15512 31168 15564
rect 31484 15512 31536 15564
rect 32404 15512 32456 15564
rect 34980 15648 35032 15700
rect 35624 15648 35676 15700
rect 34428 15580 34480 15632
rect 37280 15648 37332 15700
rect 37740 15691 37792 15700
rect 37740 15657 37749 15691
rect 37749 15657 37783 15691
rect 37783 15657 37792 15691
rect 37740 15648 37792 15657
rect 41788 15691 41840 15700
rect 41788 15657 41797 15691
rect 41797 15657 41831 15691
rect 41831 15657 41840 15691
rect 41788 15648 41840 15657
rect 42064 15691 42116 15700
rect 42064 15657 42073 15691
rect 42073 15657 42107 15691
rect 42107 15657 42116 15691
rect 42064 15648 42116 15657
rect 48688 15648 48740 15700
rect 37464 15580 37516 15632
rect 27160 15444 27212 15496
rect 27712 15444 27764 15496
rect 940 15376 992 15428
rect 4712 15376 4764 15428
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 10968 15376 11020 15428
rect 11980 15376 12032 15428
rect 12532 15376 12584 15428
rect 16764 15376 16816 15428
rect 17132 15419 17184 15428
rect 17132 15385 17141 15419
rect 17141 15385 17175 15419
rect 17175 15385 17184 15419
rect 17132 15376 17184 15385
rect 17868 15376 17920 15428
rect 21272 15376 21324 15428
rect 11888 15308 11940 15360
rect 13544 15308 13596 15360
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 16304 15308 16356 15360
rect 16396 15308 16448 15360
rect 18696 15308 18748 15360
rect 19984 15308 20036 15360
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 20352 15308 20404 15360
rect 20904 15308 20956 15360
rect 21456 15308 21508 15360
rect 21916 15376 21968 15428
rect 22192 15351 22244 15360
rect 22192 15317 22201 15351
rect 22201 15317 22235 15351
rect 22235 15317 22244 15351
rect 22192 15308 22244 15317
rect 25964 15376 26016 15428
rect 26332 15419 26384 15428
rect 26332 15385 26341 15419
rect 26341 15385 26375 15419
rect 26375 15385 26384 15419
rect 26332 15376 26384 15385
rect 27252 15376 27304 15428
rect 28356 15376 28408 15428
rect 30104 15376 30156 15428
rect 31852 15444 31904 15496
rect 34796 15512 34848 15564
rect 35900 15512 35952 15564
rect 37372 15512 37424 15564
rect 39488 15555 39540 15564
rect 39488 15521 39497 15555
rect 39497 15521 39531 15555
rect 39531 15521 39540 15555
rect 39488 15512 39540 15521
rect 40316 15555 40368 15564
rect 40316 15521 40325 15555
rect 40325 15521 40359 15555
rect 40359 15521 40368 15555
rect 40316 15512 40368 15521
rect 34060 15444 34112 15496
rect 49332 15487 49384 15496
rect 49332 15453 49341 15487
rect 49341 15453 49375 15487
rect 49375 15453 49384 15487
rect 49332 15444 49384 15453
rect 30656 15376 30708 15428
rect 30748 15419 30800 15428
rect 30748 15385 30757 15419
rect 30757 15385 30791 15419
rect 30791 15385 30800 15419
rect 30748 15376 30800 15385
rect 35072 15376 35124 15428
rect 38660 15376 38712 15428
rect 39212 15419 39264 15428
rect 39212 15385 39221 15419
rect 39221 15385 39255 15419
rect 39255 15385 39264 15419
rect 39212 15376 39264 15385
rect 39948 15376 40000 15428
rect 25228 15308 25280 15360
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 26424 15308 26476 15360
rect 26976 15351 27028 15360
rect 26976 15317 26985 15351
rect 26985 15317 27019 15351
rect 27019 15317 27028 15351
rect 26976 15308 27028 15317
rect 27436 15351 27488 15360
rect 27436 15317 27445 15351
rect 27445 15317 27479 15351
rect 27479 15317 27488 15351
rect 27436 15308 27488 15317
rect 29368 15351 29420 15360
rect 29368 15317 29377 15351
rect 29377 15317 29411 15351
rect 29411 15317 29420 15351
rect 29368 15308 29420 15317
rect 30840 15308 30892 15360
rect 32312 15308 32364 15360
rect 33508 15308 33560 15360
rect 33876 15351 33928 15360
rect 33876 15317 33885 15351
rect 33885 15317 33919 15351
rect 33919 15317 33928 15351
rect 33876 15308 33928 15317
rect 35348 15308 35400 15360
rect 36452 15308 36504 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 11796 15104 11848 15156
rect 11980 15104 12032 15156
rect 12348 15104 12400 15156
rect 12900 15104 12952 15156
rect 13912 15104 13964 15156
rect 10876 15079 10928 15088
rect 10876 15045 10885 15079
rect 10885 15045 10919 15079
rect 10919 15045 10928 15079
rect 10876 15036 10928 15045
rect 10968 15036 11020 15088
rect 11612 15036 11664 15088
rect 940 14968 992 15020
rect 4712 14968 4764 15020
rect 10600 14968 10652 15020
rect 13452 15036 13504 15088
rect 14280 15036 14332 15088
rect 14556 15104 14608 15156
rect 14740 15036 14792 15088
rect 16028 15036 16080 15088
rect 19432 15104 19484 15156
rect 21456 15104 21508 15156
rect 23756 15104 23808 15156
rect 24768 15104 24820 15156
rect 9772 14900 9824 14952
rect 11980 14832 12032 14884
rect 12072 14832 12124 14884
rect 14464 14900 14516 14952
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 18696 14968 18748 15020
rect 20812 15036 20864 15088
rect 21180 15036 21232 15088
rect 25872 15036 25924 15088
rect 14832 14900 14884 14909
rect 15660 14900 15712 14952
rect 15384 14832 15436 14884
rect 16948 14900 17000 14952
rect 18788 14943 18840 14952
rect 16304 14832 16356 14884
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 12532 14764 12584 14816
rect 14280 14764 14332 14816
rect 14740 14764 14792 14816
rect 15936 14764 15988 14816
rect 17224 14832 17276 14884
rect 18788 14909 18797 14943
rect 18797 14909 18831 14943
rect 18831 14909 18840 14943
rect 18788 14900 18840 14909
rect 19524 14968 19576 15020
rect 20904 14968 20956 15020
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 20536 14900 20588 14952
rect 20628 14900 20680 14952
rect 21272 14943 21324 14952
rect 21272 14909 21281 14943
rect 21281 14909 21315 14943
rect 21315 14909 21324 14943
rect 21272 14900 21324 14909
rect 21916 14900 21968 14952
rect 23940 14968 23992 15020
rect 24952 14968 25004 15020
rect 25228 14968 25280 15020
rect 25964 14968 26016 15020
rect 26240 15011 26292 15020
rect 26240 14977 26249 15011
rect 26249 14977 26283 15011
rect 26283 14977 26292 15011
rect 26240 14968 26292 14977
rect 23572 14943 23624 14952
rect 23572 14909 23581 14943
rect 23581 14909 23615 14943
rect 23615 14909 23624 14943
rect 23572 14900 23624 14909
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 24860 14900 24912 14952
rect 27252 15104 27304 15156
rect 27528 15147 27580 15156
rect 27528 15113 27537 15147
rect 27537 15113 27571 15147
rect 27571 15113 27580 15147
rect 27528 15104 27580 15113
rect 28448 15104 28500 15156
rect 29828 15104 29880 15156
rect 30656 15104 30708 15156
rect 31300 15104 31352 15156
rect 32036 15104 32088 15156
rect 33784 15104 33836 15156
rect 33876 15147 33928 15156
rect 33876 15113 33885 15147
rect 33885 15113 33919 15147
rect 33919 15113 33928 15147
rect 33876 15104 33928 15113
rect 35624 15104 35676 15156
rect 36084 15104 36136 15156
rect 38660 15104 38712 15156
rect 27252 15011 27304 15020
rect 27252 14977 27261 15011
rect 27261 14977 27295 15011
rect 27295 14977 27304 15011
rect 27252 14968 27304 14977
rect 27804 14968 27856 15020
rect 29368 14968 29420 15020
rect 29552 14968 29604 15020
rect 17500 14832 17552 14884
rect 21088 14832 21140 14884
rect 21456 14832 21508 14884
rect 22836 14832 22888 14884
rect 22376 14764 22428 14816
rect 22652 14764 22704 14816
rect 27160 14900 27212 14952
rect 30288 14900 30340 14952
rect 30380 14900 30432 14952
rect 32312 15036 32364 15088
rect 31760 14968 31812 15020
rect 34244 15036 34296 15088
rect 34888 15036 34940 15088
rect 35808 15036 35860 15088
rect 36360 15036 36412 15088
rect 37648 15036 37700 15088
rect 37740 15079 37792 15088
rect 37740 15045 37749 15079
rect 37749 15045 37783 15079
rect 37783 15045 37792 15079
rect 37740 15036 37792 15045
rect 38752 15036 38804 15088
rect 48412 15036 48464 15088
rect 33968 14968 34020 15020
rect 24952 14764 25004 14816
rect 25412 14764 25464 14816
rect 27988 14764 28040 14816
rect 31484 14832 31536 14884
rect 33784 14943 33836 14952
rect 33784 14909 33793 14943
rect 33793 14909 33827 14943
rect 33827 14909 33836 14943
rect 33784 14900 33836 14909
rect 35900 14900 35952 14952
rect 35992 14943 36044 14952
rect 35992 14909 36001 14943
rect 36001 14909 36035 14943
rect 36035 14909 36044 14943
rect 35992 14900 36044 14909
rect 36084 14900 36136 14952
rect 37096 14900 37148 14952
rect 37372 14968 37424 15020
rect 40868 15011 40920 15020
rect 40868 14977 40877 15011
rect 40877 14977 40911 15011
rect 40911 14977 40920 15011
rect 40868 14968 40920 14977
rect 49332 15011 49384 15020
rect 49332 14977 49341 15011
rect 49341 14977 49375 15011
rect 49375 14977 49384 15011
rect 49332 14968 49384 14977
rect 37832 14900 37884 14952
rect 38292 14900 38344 14952
rect 39396 14900 39448 14952
rect 30196 14807 30248 14816
rect 30196 14773 30205 14807
rect 30205 14773 30239 14807
rect 30239 14773 30248 14807
rect 30196 14764 30248 14773
rect 30380 14764 30432 14816
rect 34244 14807 34296 14816
rect 34244 14773 34253 14807
rect 34253 14773 34287 14807
rect 34287 14773 34296 14807
rect 34244 14764 34296 14773
rect 36360 14764 36412 14816
rect 36820 14764 36872 14816
rect 49148 14875 49200 14884
rect 49148 14841 49157 14875
rect 49157 14841 49191 14875
rect 49191 14841 49200 14875
rect 49148 14832 49200 14841
rect 45652 14764 45704 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 11244 14560 11296 14612
rect 12808 14560 12860 14612
rect 10232 14535 10284 14544
rect 10232 14501 10241 14535
rect 10241 14501 10275 14535
rect 10275 14501 10284 14535
rect 10232 14492 10284 14501
rect 14004 14560 14056 14612
rect 14188 14603 14240 14612
rect 14188 14569 14197 14603
rect 14197 14569 14231 14603
rect 14231 14569 14240 14603
rect 14188 14560 14240 14569
rect 14648 14560 14700 14612
rect 18420 14560 18472 14612
rect 940 14424 992 14476
rect 9956 14356 10008 14408
rect 13452 14492 13504 14544
rect 13268 14424 13320 14476
rect 13360 14424 13412 14476
rect 13636 14424 13688 14476
rect 14832 14424 14884 14476
rect 13820 14356 13872 14408
rect 15016 14356 15068 14408
rect 15384 14424 15436 14476
rect 17408 14356 17460 14408
rect 20076 14467 20128 14476
rect 20076 14433 20085 14467
rect 20085 14433 20119 14467
rect 20119 14433 20128 14467
rect 20076 14424 20128 14433
rect 21088 14467 21140 14476
rect 21088 14433 21097 14467
rect 21097 14433 21131 14467
rect 21131 14433 21140 14467
rect 21088 14424 21140 14433
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 21456 14424 21508 14476
rect 22744 14492 22796 14544
rect 23112 14560 23164 14612
rect 24584 14603 24636 14612
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 24860 14560 24912 14612
rect 25504 14560 25556 14612
rect 26332 14560 26384 14612
rect 26516 14560 26568 14612
rect 30380 14560 30432 14612
rect 33784 14560 33836 14612
rect 34244 14560 34296 14612
rect 29276 14492 29328 14544
rect 29736 14492 29788 14544
rect 33324 14492 33376 14544
rect 33508 14492 33560 14544
rect 36360 14560 36412 14612
rect 36820 14560 36872 14612
rect 38752 14560 38804 14612
rect 39948 14603 40000 14612
rect 39948 14569 39957 14603
rect 39957 14569 39991 14603
rect 39991 14569 40000 14603
rect 39948 14560 40000 14569
rect 27896 14424 27948 14476
rect 28724 14424 28776 14476
rect 30564 14424 30616 14476
rect 30748 14424 30800 14476
rect 32404 14424 32456 14476
rect 32588 14424 32640 14476
rect 34796 14424 34848 14476
rect 37556 14492 37608 14544
rect 49056 14535 49108 14544
rect 49056 14501 49065 14535
rect 49065 14501 49099 14535
rect 49099 14501 49108 14535
rect 49056 14492 49108 14501
rect 37280 14424 37332 14476
rect 37372 14424 37424 14476
rect 17684 14356 17736 14408
rect 19340 14356 19392 14408
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 27620 14356 27672 14408
rect 30012 14356 30064 14408
rect 30104 14399 30156 14408
rect 30104 14365 30113 14399
rect 30113 14365 30147 14399
rect 30147 14365 30156 14399
rect 30104 14356 30156 14365
rect 30840 14356 30892 14408
rect 32864 14356 32916 14408
rect 33692 14399 33744 14408
rect 33692 14365 33701 14399
rect 33701 14365 33735 14399
rect 33735 14365 33744 14399
rect 33692 14356 33744 14365
rect 39304 14399 39356 14408
rect 39304 14365 39313 14399
rect 39313 14365 39347 14399
rect 39347 14365 39356 14399
rect 39304 14356 39356 14365
rect 49240 14399 49292 14408
rect 49240 14365 49249 14399
rect 49249 14365 49283 14399
rect 49283 14365 49292 14399
rect 49240 14356 49292 14365
rect 10416 14331 10468 14340
rect 10416 14297 10425 14331
rect 10425 14297 10459 14331
rect 10459 14297 10468 14331
rect 10416 14288 10468 14297
rect 11244 14331 11296 14340
rect 11244 14297 11253 14331
rect 11253 14297 11287 14331
rect 11287 14297 11296 14331
rect 11244 14288 11296 14297
rect 12808 14288 12860 14340
rect 10508 14220 10560 14272
rect 12624 14220 12676 14272
rect 13912 14220 13964 14272
rect 14832 14263 14884 14272
rect 14832 14229 14841 14263
rect 14841 14229 14875 14263
rect 14875 14229 14884 14263
rect 14832 14220 14884 14229
rect 16580 14220 16632 14272
rect 16856 14263 16908 14272
rect 16856 14229 16865 14263
rect 16865 14229 16899 14263
rect 16899 14229 16908 14263
rect 16856 14220 16908 14229
rect 17224 14220 17276 14272
rect 19432 14288 19484 14340
rect 19984 14331 20036 14340
rect 19984 14297 19993 14331
rect 19993 14297 20027 14331
rect 20027 14297 20036 14331
rect 19984 14288 20036 14297
rect 21456 14288 21508 14340
rect 21824 14288 21876 14340
rect 25780 14288 25832 14340
rect 27068 14331 27120 14340
rect 27068 14297 27077 14331
rect 27077 14297 27111 14331
rect 27111 14297 27120 14331
rect 27068 14288 27120 14297
rect 27712 14288 27764 14340
rect 18420 14220 18472 14272
rect 18972 14220 19024 14272
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 20720 14263 20772 14272
rect 20720 14229 20729 14263
rect 20729 14229 20763 14263
rect 20763 14229 20772 14263
rect 20720 14220 20772 14229
rect 21548 14220 21600 14272
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 25136 14263 25188 14272
rect 25136 14229 25145 14263
rect 25145 14229 25179 14263
rect 25179 14229 25188 14263
rect 25136 14220 25188 14229
rect 27528 14220 27580 14272
rect 28448 14220 28500 14272
rect 31484 14288 31536 14340
rect 32036 14288 32088 14340
rect 35164 14331 35216 14340
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 35440 14288 35492 14340
rect 36636 14288 36688 14340
rect 38292 14288 38344 14340
rect 29000 14263 29052 14272
rect 29000 14229 29009 14263
rect 29009 14229 29043 14263
rect 29043 14229 29052 14263
rect 29000 14220 29052 14229
rect 29644 14220 29696 14272
rect 30380 14220 30432 14272
rect 32772 14220 32824 14272
rect 33692 14220 33744 14272
rect 35348 14220 35400 14272
rect 35808 14220 35860 14272
rect 35900 14220 35952 14272
rect 39396 14220 39448 14272
rect 39488 14263 39540 14272
rect 39488 14229 39497 14263
rect 39497 14229 39531 14263
rect 39531 14229 39540 14263
rect 39488 14220 39540 14229
rect 48320 14220 48372 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 12348 14016 12400 14068
rect 14280 14016 14332 14068
rect 1032 13948 1084 14000
rect 10508 13948 10560 14000
rect 11244 13948 11296 14000
rect 13268 13991 13320 14000
rect 13268 13957 13277 13991
rect 13277 13957 13311 13991
rect 13311 13957 13320 13991
rect 13268 13948 13320 13957
rect 15200 14016 15252 14068
rect 15936 14016 15988 14068
rect 16580 14016 16632 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 19064 14016 19116 14068
rect 19892 14016 19944 14068
rect 21364 14016 21416 14068
rect 25320 14016 25372 14068
rect 25504 14016 25556 14068
rect 14740 13948 14792 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 10324 13812 10376 13864
rect 9772 13676 9824 13728
rect 12072 13744 12124 13796
rect 13636 13812 13688 13864
rect 15844 13880 15896 13932
rect 19524 13948 19576 14000
rect 20628 13948 20680 14000
rect 21824 13948 21876 14000
rect 24032 13948 24084 14000
rect 25780 13948 25832 14000
rect 16764 13880 16816 13932
rect 17684 13880 17736 13932
rect 18420 13880 18472 13932
rect 18696 13880 18748 13932
rect 19432 13880 19484 13932
rect 27528 14016 27580 14068
rect 28816 14016 28868 14068
rect 30012 14016 30064 14068
rect 31116 14016 31168 14068
rect 31852 13948 31904 14000
rect 33324 13948 33376 14000
rect 34428 14016 34480 14068
rect 35716 14016 35768 14068
rect 35808 14016 35860 14068
rect 41328 14016 41380 14068
rect 47860 14016 47912 14068
rect 48412 14059 48464 14068
rect 48412 14025 48421 14059
rect 48421 14025 48455 14059
rect 48455 14025 48464 14059
rect 48412 14016 48464 14025
rect 48872 14016 48924 14068
rect 28908 13923 28960 13932
rect 28908 13889 28917 13923
rect 28917 13889 28951 13923
rect 28951 13889 28960 13923
rect 28908 13880 28960 13889
rect 31116 13923 31168 13932
rect 31116 13889 31125 13923
rect 31125 13889 31159 13923
rect 31159 13889 31168 13923
rect 31116 13880 31168 13889
rect 34704 13880 34756 13932
rect 15108 13812 15160 13864
rect 14464 13744 14516 13796
rect 18604 13812 18656 13864
rect 18972 13812 19024 13864
rect 20720 13812 20772 13864
rect 21916 13812 21968 13864
rect 12348 13676 12400 13728
rect 12716 13676 12768 13728
rect 16304 13676 16356 13728
rect 17960 13744 18012 13796
rect 23940 13812 23992 13864
rect 27068 13812 27120 13864
rect 32312 13855 32364 13864
rect 24584 13744 24636 13796
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 34060 13855 34112 13864
rect 34060 13821 34069 13855
rect 34069 13821 34103 13855
rect 34103 13821 34112 13855
rect 34060 13812 34112 13821
rect 36176 13880 36228 13932
rect 36360 13880 36412 13932
rect 36728 13948 36780 14000
rect 38660 13948 38712 14000
rect 38844 13948 38896 14000
rect 39488 13948 39540 14000
rect 49240 13991 49292 14000
rect 49240 13957 49249 13991
rect 49249 13957 49283 13991
rect 49283 13957 49292 13991
rect 49240 13948 49292 13957
rect 45652 13923 45704 13932
rect 45652 13889 45661 13923
rect 45661 13889 45695 13923
rect 45695 13889 45704 13923
rect 45652 13880 45704 13889
rect 48228 13880 48280 13932
rect 35992 13855 36044 13864
rect 35992 13821 36001 13855
rect 36001 13821 36035 13855
rect 36035 13821 36044 13855
rect 35992 13812 36044 13821
rect 36268 13812 36320 13864
rect 36636 13812 36688 13864
rect 34704 13744 34756 13796
rect 46572 13812 46624 13864
rect 38200 13744 38252 13796
rect 23112 13676 23164 13728
rect 24676 13676 24728 13728
rect 25688 13676 25740 13728
rect 30840 13676 30892 13728
rect 35900 13676 35952 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 13728 13515 13780 13524
rect 13728 13481 13737 13515
rect 13737 13481 13771 13515
rect 13771 13481 13780 13515
rect 13728 13472 13780 13481
rect 14004 13472 14056 13524
rect 15016 13472 15068 13524
rect 14740 13404 14792 13456
rect 10784 13379 10836 13388
rect 10784 13345 10793 13379
rect 10793 13345 10827 13379
rect 10827 13345 10836 13379
rect 10784 13336 10836 13345
rect 12072 13336 12124 13388
rect 12348 13336 12400 13388
rect 9036 13200 9088 13252
rect 10876 13132 10928 13184
rect 10968 13132 11020 13184
rect 12348 13200 12400 13252
rect 12808 13336 12860 13388
rect 13820 13336 13872 13388
rect 14004 13336 14056 13388
rect 15108 13336 15160 13388
rect 17960 13472 18012 13524
rect 18420 13472 18472 13524
rect 19156 13472 19208 13524
rect 20076 13472 20128 13524
rect 20260 13472 20312 13524
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 22100 13515 22152 13524
rect 22100 13481 22109 13515
rect 22109 13481 22143 13515
rect 22143 13481 22152 13515
rect 22100 13472 22152 13481
rect 16120 13404 16172 13456
rect 15476 13379 15528 13388
rect 15476 13345 15485 13379
rect 15485 13345 15519 13379
rect 15519 13345 15528 13379
rect 15476 13336 15528 13345
rect 15752 13336 15804 13388
rect 16304 13336 16356 13388
rect 18512 13404 18564 13456
rect 22468 13404 22520 13456
rect 20720 13336 20772 13388
rect 21364 13336 21416 13388
rect 22744 13472 22796 13524
rect 23664 13472 23716 13524
rect 25596 13515 25648 13524
rect 25596 13481 25605 13515
rect 25605 13481 25639 13515
rect 25639 13481 25648 13515
rect 25596 13472 25648 13481
rect 25780 13472 25832 13524
rect 27528 13472 27580 13524
rect 27712 13515 27764 13524
rect 27712 13481 27721 13515
rect 27721 13481 27755 13515
rect 27755 13481 27764 13515
rect 27712 13472 27764 13481
rect 27804 13515 27856 13524
rect 27804 13481 27813 13515
rect 27813 13481 27847 13515
rect 27847 13481 27856 13515
rect 27804 13472 27856 13481
rect 28356 13472 28408 13524
rect 28908 13472 28960 13524
rect 33784 13472 33836 13524
rect 35532 13472 35584 13524
rect 36268 13472 36320 13524
rect 24860 13404 24912 13456
rect 23020 13336 23072 13388
rect 14280 13268 14332 13320
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 24032 13336 24084 13388
rect 24400 13336 24452 13388
rect 27068 13336 27120 13388
rect 29920 13404 29972 13456
rect 30380 13404 30432 13456
rect 29828 13379 29880 13388
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 30472 13336 30524 13388
rect 31576 13336 31628 13388
rect 33692 13404 33744 13456
rect 38200 13515 38252 13524
rect 38200 13481 38209 13515
rect 38209 13481 38243 13515
rect 38243 13481 38252 13515
rect 38200 13472 38252 13481
rect 38844 13472 38896 13524
rect 33876 13379 33928 13388
rect 33876 13345 33885 13379
rect 33885 13345 33919 13379
rect 33919 13345 33928 13379
rect 33876 13336 33928 13345
rect 39212 13404 39264 13456
rect 36360 13336 36412 13388
rect 36820 13336 36872 13388
rect 39488 13336 39540 13388
rect 24676 13268 24728 13320
rect 25136 13268 25188 13320
rect 14924 13200 14976 13252
rect 13820 13132 13872 13184
rect 14096 13132 14148 13184
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 17132 13200 17184 13252
rect 21180 13200 21232 13252
rect 21640 13200 21692 13252
rect 22836 13200 22888 13252
rect 23664 13243 23716 13252
rect 23664 13209 23673 13243
rect 23673 13209 23707 13243
rect 23707 13209 23716 13243
rect 23664 13200 23716 13209
rect 27436 13268 27488 13320
rect 29000 13268 29052 13320
rect 30196 13268 30248 13320
rect 34060 13268 34112 13320
rect 34888 13268 34940 13320
rect 19892 13132 19944 13184
rect 20260 13132 20312 13184
rect 21272 13175 21324 13184
rect 21272 13141 21281 13175
rect 21281 13141 21315 13175
rect 21315 13141 21324 13175
rect 21272 13132 21324 13141
rect 21732 13132 21784 13184
rect 26056 13243 26108 13252
rect 26056 13209 26065 13243
rect 26065 13209 26099 13243
rect 26099 13209 26108 13243
rect 26056 13200 26108 13209
rect 23848 13132 23900 13184
rect 26516 13132 26568 13184
rect 28724 13175 28776 13184
rect 28724 13141 28733 13175
rect 28733 13141 28767 13175
rect 28767 13141 28776 13175
rect 28724 13132 28776 13141
rect 31668 13132 31720 13184
rect 31852 13132 31904 13184
rect 33968 13200 34020 13252
rect 35164 13243 35216 13252
rect 35164 13209 35173 13243
rect 35173 13209 35207 13243
rect 35207 13209 35216 13243
rect 35164 13200 35216 13209
rect 36360 13200 36412 13252
rect 41328 13311 41380 13320
rect 41328 13277 41337 13311
rect 41337 13277 41371 13311
rect 41371 13277 41380 13311
rect 41328 13268 41380 13277
rect 46572 13268 46624 13320
rect 49148 13311 49200 13320
rect 49148 13277 49157 13311
rect 49157 13277 49191 13311
rect 49191 13277 49200 13311
rect 49148 13268 49200 13277
rect 33324 13132 33376 13184
rect 33692 13175 33744 13184
rect 33692 13141 33701 13175
rect 33701 13141 33735 13175
rect 33735 13141 33744 13175
rect 33692 13132 33744 13141
rect 34336 13132 34388 13184
rect 36636 13200 36688 13252
rect 37464 13132 37516 13184
rect 37648 13132 37700 13184
rect 39304 13132 39356 13184
rect 45928 13132 45980 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 5448 12928 5500 12980
rect 10968 12971 11020 12980
rect 10968 12937 10977 12971
rect 10977 12937 11011 12971
rect 11011 12937 11020 12971
rect 10968 12928 11020 12937
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 12164 12928 12216 12980
rect 12532 12928 12584 12980
rect 13268 12928 13320 12980
rect 13636 12928 13688 12980
rect 1308 12860 1360 12912
rect 14648 12860 14700 12912
rect 15016 12928 15068 12980
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 15476 12860 15528 12912
rect 16212 12860 16264 12912
rect 16304 12860 16356 12912
rect 18972 12860 19024 12912
rect 20720 12971 20772 12980
rect 20720 12937 20729 12971
rect 20729 12937 20763 12971
rect 20763 12937 20772 12971
rect 20720 12928 20772 12937
rect 22652 12928 22704 12980
rect 22928 12971 22980 12980
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 23020 12928 23072 12980
rect 23664 12928 23716 12980
rect 24584 12928 24636 12980
rect 23848 12860 23900 12912
rect 24860 12860 24912 12912
rect 25320 12903 25372 12912
rect 25320 12869 25329 12903
rect 25329 12869 25363 12903
rect 25363 12869 25372 12903
rect 25320 12860 25372 12869
rect 1216 12792 1268 12844
rect 17040 12792 17092 12844
rect 18880 12792 18932 12844
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 21916 12792 21968 12844
rect 22192 12792 22244 12844
rect 22652 12792 22704 12844
rect 25780 12928 25832 12980
rect 26424 12928 26476 12980
rect 26516 12928 26568 12980
rect 27068 12928 27120 12980
rect 27896 12928 27948 12980
rect 27528 12860 27580 12912
rect 29644 12903 29696 12912
rect 29644 12869 29653 12903
rect 29653 12869 29687 12903
rect 29687 12869 29696 12903
rect 29644 12860 29696 12869
rect 30196 12860 30248 12912
rect 32404 12928 32456 12980
rect 32588 12928 32640 12980
rect 33692 12928 33744 12980
rect 34060 12928 34112 12980
rect 35164 12928 35216 12980
rect 40316 12928 40368 12980
rect 34888 12860 34940 12912
rect 35808 12903 35860 12912
rect 35808 12869 35817 12903
rect 35817 12869 35851 12903
rect 35851 12869 35860 12903
rect 35808 12860 35860 12869
rect 9496 12724 9548 12776
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 12440 12724 12492 12776
rect 13544 12724 13596 12776
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 15476 12724 15528 12776
rect 16120 12724 16172 12776
rect 19524 12724 19576 12776
rect 19708 12767 19760 12776
rect 19708 12733 19717 12767
rect 19717 12733 19751 12767
rect 19751 12733 19760 12767
rect 19708 12724 19760 12733
rect 20168 12724 20220 12776
rect 20444 12724 20496 12776
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 22100 12724 22152 12776
rect 12716 12656 12768 12708
rect 12900 12656 12952 12708
rect 15292 12656 15344 12708
rect 15844 12656 15896 12708
rect 11152 12588 11204 12640
rect 12532 12588 12584 12640
rect 12624 12588 12676 12640
rect 15568 12588 15620 12640
rect 17132 12656 17184 12708
rect 17776 12656 17828 12708
rect 16304 12631 16356 12640
rect 16304 12597 16313 12631
rect 16313 12597 16347 12631
rect 16347 12597 16356 12631
rect 16304 12588 16356 12597
rect 19340 12588 19392 12640
rect 21548 12656 21600 12708
rect 22928 12656 22980 12708
rect 23388 12699 23440 12708
rect 23388 12665 23397 12699
rect 23397 12665 23431 12699
rect 23431 12665 23440 12699
rect 23388 12656 23440 12665
rect 23572 12724 23624 12776
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 30012 12835 30064 12844
rect 30012 12801 30021 12835
rect 30021 12801 30055 12835
rect 30055 12801 30064 12835
rect 30012 12792 30064 12801
rect 31852 12792 31904 12844
rect 32128 12792 32180 12844
rect 34428 12792 34480 12844
rect 36084 12860 36136 12912
rect 36544 12860 36596 12912
rect 36912 12860 36964 12912
rect 37648 12860 37700 12912
rect 36820 12792 36872 12844
rect 37464 12835 37516 12844
rect 37464 12801 37473 12835
rect 37473 12801 37507 12835
rect 37507 12801 37516 12835
rect 37464 12792 37516 12801
rect 38844 12792 38896 12844
rect 40040 12835 40092 12844
rect 40040 12801 40049 12835
rect 40049 12801 40083 12835
rect 40083 12801 40092 12835
rect 40040 12792 40092 12801
rect 45928 12835 45980 12844
rect 45928 12801 45937 12835
rect 45937 12801 45971 12835
rect 45971 12801 45980 12835
rect 45928 12792 45980 12801
rect 47860 12792 47912 12844
rect 49148 12835 49200 12844
rect 49148 12801 49157 12835
rect 49157 12801 49191 12835
rect 49191 12801 49200 12835
rect 49148 12792 49200 12801
rect 26056 12724 26108 12776
rect 21272 12588 21324 12640
rect 24032 12588 24084 12640
rect 26792 12724 26844 12776
rect 28908 12767 28960 12776
rect 28908 12733 28917 12767
rect 28917 12733 28951 12767
rect 28951 12733 28960 12767
rect 28908 12724 28960 12733
rect 33876 12724 33928 12776
rect 34796 12724 34848 12776
rect 27804 12588 27856 12640
rect 34520 12656 34572 12708
rect 33324 12588 33376 12640
rect 34244 12588 34296 12640
rect 35440 12588 35492 12640
rect 37004 12724 37056 12776
rect 38292 12724 38344 12776
rect 39304 12724 39356 12776
rect 36912 12588 36964 12640
rect 37004 12631 37056 12640
rect 37004 12597 37013 12631
rect 37013 12597 37047 12631
rect 37047 12597 37056 12631
rect 37004 12588 37056 12597
rect 46756 12656 46808 12708
rect 39120 12588 39172 12640
rect 47952 12588 48004 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 11796 12384 11848 12436
rect 11980 12384 12032 12436
rect 1308 12248 1360 12300
rect 10784 12248 10836 12300
rect 12348 12248 12400 12300
rect 5816 12180 5868 12232
rect 10876 12180 10928 12232
rect 14832 12248 14884 12300
rect 15476 12248 15528 12300
rect 15752 12248 15804 12300
rect 14740 12180 14792 12232
rect 16672 12384 16724 12436
rect 21548 12384 21600 12436
rect 22468 12384 22520 12436
rect 23480 12316 23532 12368
rect 17408 12291 17460 12300
rect 17408 12257 17417 12291
rect 17417 12257 17451 12291
rect 17451 12257 17460 12291
rect 17408 12248 17460 12257
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 9772 12155 9824 12164
rect 9772 12121 9781 12155
rect 9781 12121 9815 12155
rect 9815 12121 9824 12155
rect 9772 12112 9824 12121
rect 11060 12112 11112 12164
rect 13452 12112 13504 12164
rect 14188 12044 14240 12096
rect 15568 12112 15620 12164
rect 18604 12112 18656 12164
rect 18880 12155 18932 12164
rect 18880 12121 18889 12155
rect 18889 12121 18923 12155
rect 18923 12121 18932 12155
rect 18880 12112 18932 12121
rect 19248 12112 19300 12164
rect 19892 12248 19944 12300
rect 22100 12248 22152 12300
rect 19524 12180 19576 12232
rect 20996 12180 21048 12232
rect 21732 12180 21784 12232
rect 26700 12384 26752 12436
rect 27896 12384 27948 12436
rect 31852 12427 31904 12436
rect 31852 12393 31861 12427
rect 31861 12393 31895 12427
rect 31895 12393 31904 12427
rect 31852 12384 31904 12393
rect 33876 12427 33928 12436
rect 33876 12393 33885 12427
rect 33885 12393 33919 12427
rect 33919 12393 33928 12427
rect 33876 12384 33928 12393
rect 26332 12359 26384 12368
rect 26332 12325 26341 12359
rect 26341 12325 26375 12359
rect 26375 12325 26384 12359
rect 26332 12316 26384 12325
rect 27344 12316 27396 12368
rect 34244 12359 34296 12368
rect 34244 12325 34253 12359
rect 34253 12325 34287 12359
rect 34287 12325 34296 12359
rect 34244 12316 34296 12325
rect 24860 12248 24912 12300
rect 26884 12248 26936 12300
rect 27068 12291 27120 12300
rect 27068 12257 27077 12291
rect 27077 12257 27111 12291
rect 27111 12257 27120 12291
rect 27068 12248 27120 12257
rect 30012 12248 30064 12300
rect 32404 12291 32456 12300
rect 32404 12257 32413 12291
rect 32413 12257 32447 12291
rect 32447 12257 32456 12291
rect 32404 12248 32456 12257
rect 16672 12044 16724 12096
rect 16764 12087 16816 12096
rect 16764 12053 16773 12087
rect 16773 12053 16807 12087
rect 16807 12053 16816 12087
rect 16764 12044 16816 12053
rect 20628 12044 20680 12096
rect 22376 12155 22428 12164
rect 22376 12121 22385 12155
rect 22385 12121 22419 12155
rect 22419 12121 22428 12155
rect 22376 12112 22428 12121
rect 22468 12155 22520 12164
rect 22468 12121 22477 12155
rect 22477 12121 22511 12155
rect 22511 12121 22520 12155
rect 22468 12112 22520 12121
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 25872 12180 25924 12232
rect 27528 12180 27580 12232
rect 32128 12223 32180 12232
rect 32128 12189 32137 12223
rect 32137 12189 32171 12223
rect 32171 12189 32180 12223
rect 32128 12180 32180 12189
rect 33508 12180 33560 12232
rect 34796 12248 34848 12300
rect 38844 12384 38896 12436
rect 39304 12427 39356 12436
rect 39304 12393 39313 12427
rect 39313 12393 39347 12427
rect 39347 12393 39356 12427
rect 39304 12384 39356 12393
rect 37372 12291 37424 12300
rect 37372 12257 37381 12291
rect 37381 12257 37415 12291
rect 37415 12257 37424 12291
rect 37372 12248 37424 12257
rect 38384 12291 38436 12300
rect 38384 12257 38393 12291
rect 38393 12257 38427 12291
rect 38427 12257 38436 12291
rect 38384 12248 38436 12257
rect 38752 12248 38804 12300
rect 47216 12316 47268 12368
rect 34888 12223 34940 12232
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 49148 12291 49200 12300
rect 49148 12257 49157 12291
rect 49157 12257 49191 12291
rect 49191 12257 49200 12291
rect 49148 12248 49200 12257
rect 23848 12112 23900 12164
rect 28816 12112 28868 12164
rect 29920 12112 29972 12164
rect 31852 12112 31904 12164
rect 35440 12112 35492 12164
rect 24216 12044 24268 12096
rect 26332 12044 26384 12096
rect 26976 12044 27028 12096
rect 27252 12087 27304 12096
rect 27252 12053 27261 12087
rect 27261 12053 27295 12087
rect 27295 12053 27304 12087
rect 27252 12044 27304 12053
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 31392 12044 31444 12096
rect 34336 12087 34388 12096
rect 34336 12053 34345 12087
rect 34345 12053 34379 12087
rect 34379 12053 34388 12087
rect 34336 12044 34388 12053
rect 36728 12044 36780 12096
rect 37556 12044 37608 12096
rect 40408 12112 40460 12164
rect 38660 12087 38712 12096
rect 38660 12053 38669 12087
rect 38669 12053 38703 12087
rect 38703 12053 38712 12087
rect 38660 12044 38712 12053
rect 40960 12087 41012 12096
rect 40960 12053 40969 12087
rect 40969 12053 41003 12087
rect 41003 12053 41012 12087
rect 40960 12044 41012 12053
rect 47952 12223 48004 12232
rect 47952 12189 47961 12223
rect 47961 12189 47995 12223
rect 47995 12189 48004 12223
rect 47952 12180 48004 12189
rect 46112 12087 46164 12096
rect 46112 12053 46121 12087
rect 46121 12053 46155 12087
rect 46155 12053 46164 12087
rect 46112 12044 46164 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 4252 11840 4304 11892
rect 10876 11840 10928 11892
rect 12348 11840 12400 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 13360 11883 13412 11892
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 13636 11840 13688 11892
rect 15200 11840 15252 11892
rect 15844 11840 15896 11892
rect 16396 11840 16448 11892
rect 17040 11840 17092 11892
rect 19248 11840 19300 11892
rect 2136 11772 2188 11824
rect 14004 11772 14056 11824
rect 14832 11772 14884 11824
rect 1216 11704 1268 11756
rect 1308 11636 1360 11688
rect 11796 11704 11848 11756
rect 14740 11704 14792 11756
rect 11428 11568 11480 11620
rect 12256 11568 12308 11620
rect 12716 11568 12768 11620
rect 13268 11636 13320 11688
rect 13636 11636 13688 11688
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 14004 11636 14056 11645
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 19340 11704 19392 11756
rect 16120 11636 16172 11688
rect 14372 11568 14424 11620
rect 15476 11568 15528 11620
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 14832 11500 14884 11552
rect 15384 11500 15436 11552
rect 16948 11568 17000 11620
rect 16212 11500 16264 11552
rect 17960 11500 18012 11552
rect 18604 11679 18656 11688
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 18880 11636 18932 11688
rect 20352 11772 20404 11824
rect 20996 11772 21048 11824
rect 21272 11772 21324 11824
rect 20076 11704 20128 11756
rect 20536 11704 20588 11756
rect 22008 11704 22060 11756
rect 27344 11840 27396 11892
rect 28724 11840 28776 11892
rect 31760 11840 31812 11892
rect 31852 11883 31904 11892
rect 31852 11849 31861 11883
rect 31861 11849 31895 11883
rect 31895 11849 31904 11883
rect 31852 11840 31904 11849
rect 31944 11840 31996 11892
rect 32772 11840 32824 11892
rect 35440 11840 35492 11892
rect 24216 11815 24268 11824
rect 24216 11781 24225 11815
rect 24225 11781 24259 11815
rect 24259 11781 24268 11815
rect 24216 11772 24268 11781
rect 25872 11772 25924 11824
rect 26148 11815 26200 11824
rect 26148 11781 26157 11815
rect 26157 11781 26191 11815
rect 26191 11781 26200 11815
rect 26148 11772 26200 11781
rect 26976 11772 27028 11824
rect 27620 11772 27672 11824
rect 31392 11772 31444 11824
rect 31576 11772 31628 11824
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 31116 11747 31168 11756
rect 31116 11713 31125 11747
rect 31125 11713 31159 11747
rect 31159 11713 31168 11747
rect 31116 11704 31168 11713
rect 20260 11611 20312 11620
rect 20260 11577 20269 11611
rect 20269 11577 20303 11611
rect 20303 11577 20312 11611
rect 20260 11568 20312 11577
rect 20812 11568 20864 11620
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 22376 11636 22428 11688
rect 22652 11568 22704 11620
rect 20444 11500 20496 11552
rect 21640 11500 21692 11552
rect 22008 11500 22060 11552
rect 24860 11636 24912 11688
rect 27160 11636 27212 11688
rect 27436 11679 27488 11688
rect 27436 11645 27445 11679
rect 27445 11645 27479 11679
rect 27479 11645 27488 11679
rect 27436 11636 27488 11645
rect 27344 11568 27396 11620
rect 29552 11636 29604 11688
rect 29644 11636 29696 11688
rect 30840 11679 30892 11688
rect 30840 11645 30849 11679
rect 30849 11645 30883 11679
rect 30883 11645 30892 11679
rect 30840 11636 30892 11645
rect 31944 11636 31996 11688
rect 32680 11636 32732 11688
rect 33876 11747 33928 11756
rect 33876 11713 33885 11747
rect 33885 11713 33919 11747
rect 33919 11713 33928 11747
rect 33876 11704 33928 11713
rect 24584 11500 24636 11552
rect 29276 11500 29328 11552
rect 30472 11500 30524 11552
rect 31392 11500 31444 11552
rect 31576 11568 31628 11620
rect 35532 11772 35584 11824
rect 35808 11840 35860 11892
rect 38660 11883 38712 11892
rect 38660 11849 38669 11883
rect 38669 11849 38703 11883
rect 38703 11849 38712 11883
rect 38660 11840 38712 11849
rect 39120 11883 39172 11892
rect 39120 11849 39129 11883
rect 39129 11849 39163 11883
rect 39163 11849 39172 11883
rect 39120 11840 39172 11849
rect 35900 11772 35952 11824
rect 37372 11772 37424 11824
rect 40960 11772 41012 11824
rect 49148 11815 49200 11824
rect 49148 11781 49157 11815
rect 49157 11781 49191 11815
rect 49191 11781 49200 11815
rect 49148 11772 49200 11781
rect 36820 11704 36872 11756
rect 39028 11747 39080 11756
rect 39028 11713 39037 11747
rect 39037 11713 39071 11747
rect 39071 11713 39080 11747
rect 39028 11704 39080 11713
rect 40408 11747 40460 11756
rect 40408 11713 40417 11747
rect 40417 11713 40451 11747
rect 40451 11713 40460 11747
rect 40408 11704 40460 11713
rect 46112 11704 46164 11756
rect 34428 11636 34480 11688
rect 34888 11636 34940 11688
rect 35072 11568 35124 11620
rect 32864 11500 32916 11552
rect 34612 11500 34664 11552
rect 36176 11636 36228 11688
rect 36636 11636 36688 11688
rect 37188 11568 37240 11620
rect 35624 11500 35676 11552
rect 35808 11500 35860 11552
rect 35992 11500 36044 11552
rect 36728 11500 36780 11552
rect 40224 11500 40276 11552
rect 46572 11568 46624 11620
rect 47032 11500 47084 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 1216 11296 1268 11348
rect 11060 11160 11112 11212
rect 11796 11160 11848 11212
rect 13912 11296 13964 11348
rect 14556 11296 14608 11348
rect 16120 11296 16172 11348
rect 16396 11296 16448 11348
rect 16856 11296 16908 11348
rect 17132 11296 17184 11348
rect 12716 11228 12768 11280
rect 14464 11160 14516 11212
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15292 11160 15344 11212
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 15936 11160 15988 11212
rect 16120 11160 16172 11212
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19432 11296 19484 11348
rect 20076 11296 20128 11348
rect 20444 11339 20496 11348
rect 20444 11305 20453 11339
rect 20453 11305 20487 11339
rect 20487 11305 20496 11339
rect 20444 11296 20496 11305
rect 19156 11228 19208 11280
rect 23296 11339 23348 11348
rect 23296 11305 23305 11339
rect 23305 11305 23339 11339
rect 23339 11305 23348 11339
rect 23296 11296 23348 11305
rect 23756 11228 23808 11280
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 17040 11092 17092 11144
rect 18328 11092 18380 11144
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 19524 11092 19576 11144
rect 12900 11024 12952 11076
rect 15568 11024 15620 11076
rect 16580 11024 16632 11076
rect 17776 11024 17828 11076
rect 17960 11024 18012 11076
rect 12532 10956 12584 11008
rect 14648 10956 14700 11008
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 18512 11024 18564 11076
rect 18604 11024 18656 11076
rect 23848 11160 23900 11212
rect 25228 11296 25280 11348
rect 26608 11296 26660 11348
rect 28816 11296 28868 11348
rect 33324 11296 33376 11348
rect 34428 11296 34480 11348
rect 35072 11296 35124 11348
rect 28908 11228 28960 11280
rect 30472 11271 30524 11280
rect 30472 11237 30481 11271
rect 30481 11237 30515 11271
rect 30515 11237 30524 11271
rect 30472 11228 30524 11237
rect 32680 11228 32732 11280
rect 32956 11228 33008 11280
rect 24860 11203 24912 11212
rect 24860 11169 24869 11203
rect 24869 11169 24903 11203
rect 24903 11169 24912 11203
rect 24860 11160 24912 11169
rect 20812 11092 20864 11144
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 28908 11092 28960 11144
rect 31484 11160 31536 11212
rect 32128 11160 32180 11212
rect 34888 11160 34940 11212
rect 37372 11160 37424 11212
rect 37464 11160 37516 11212
rect 29644 11092 29696 11144
rect 33232 11092 33284 11144
rect 33324 11135 33376 11144
rect 33324 11101 33333 11135
rect 33333 11101 33367 11135
rect 33367 11101 33376 11135
rect 33324 11092 33376 11101
rect 35900 11092 35952 11144
rect 36452 11092 36504 11144
rect 44364 11296 44416 11348
rect 38844 11228 38896 11280
rect 39488 11228 39540 11280
rect 40224 11092 40276 11144
rect 49148 11203 49200 11212
rect 49148 11169 49157 11203
rect 49157 11169 49191 11203
rect 49191 11169 49200 11203
rect 49148 11160 49200 11169
rect 46756 11092 46808 11144
rect 21640 11024 21692 11076
rect 19432 10956 19484 11008
rect 22008 10956 22060 11008
rect 22652 10999 22704 11008
rect 22652 10965 22661 10999
rect 22661 10965 22695 10999
rect 22695 10965 22704 10999
rect 22652 10956 22704 10965
rect 23940 11024 23992 11076
rect 25872 11024 25924 11076
rect 27160 11067 27212 11076
rect 27160 11033 27169 11067
rect 27169 11033 27203 11067
rect 27203 11033 27212 11067
rect 27160 11024 27212 11033
rect 27620 11024 27672 11076
rect 23572 10956 23624 11008
rect 23848 10956 23900 11008
rect 24492 10956 24544 11008
rect 29276 11024 29328 11076
rect 31392 11067 31444 11076
rect 31392 11033 31401 11067
rect 31401 11033 31435 11067
rect 31435 11033 31444 11067
rect 31392 11024 31444 11033
rect 31484 11024 31536 11076
rect 30748 10999 30800 11008
rect 30748 10965 30757 10999
rect 30757 10965 30791 10999
rect 30791 10965 30800 10999
rect 30748 10956 30800 10965
rect 35164 11024 35216 11076
rect 36084 11024 36136 11076
rect 37188 11024 37240 11076
rect 38384 11024 38436 11076
rect 33692 10956 33744 11008
rect 33968 10956 34020 11008
rect 38568 10956 38620 11008
rect 46940 11024 46992 11076
rect 46112 10956 46164 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 1216 10684 1268 10736
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 12808 10752 12860 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 17592 10752 17644 10804
rect 19432 10752 19484 10804
rect 19708 10752 19760 10804
rect 22652 10752 22704 10804
rect 22928 10752 22980 10804
rect 25872 10795 25924 10804
rect 25872 10761 25881 10795
rect 25881 10761 25915 10795
rect 25915 10761 25924 10795
rect 25872 10752 25924 10761
rect 26700 10752 26752 10804
rect 27068 10752 27120 10804
rect 30196 10752 30248 10804
rect 30840 10752 30892 10804
rect 31116 10752 31168 10804
rect 32312 10752 32364 10804
rect 32496 10752 32548 10804
rect 1308 10616 1360 10668
rect 14096 10684 14148 10736
rect 16764 10684 16816 10736
rect 17040 10684 17092 10736
rect 12256 10616 12308 10668
rect 13268 10548 13320 10600
rect 13452 10480 13504 10532
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 12532 10412 12584 10464
rect 16212 10616 16264 10668
rect 17316 10616 17368 10668
rect 18420 10616 18472 10668
rect 14556 10548 14608 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 15016 10548 15068 10600
rect 14004 10480 14056 10532
rect 16672 10548 16724 10600
rect 17592 10591 17644 10600
rect 17592 10557 17601 10591
rect 17601 10557 17635 10591
rect 17635 10557 17644 10591
rect 17592 10548 17644 10557
rect 17684 10591 17736 10600
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 18972 10616 19024 10668
rect 20996 10684 21048 10736
rect 22284 10684 22336 10736
rect 23572 10684 23624 10736
rect 26148 10684 26200 10736
rect 27436 10684 27488 10736
rect 20260 10616 20312 10668
rect 19984 10548 20036 10600
rect 21088 10548 21140 10600
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 15660 10412 15712 10464
rect 17040 10412 17092 10464
rect 21272 10480 21324 10532
rect 23388 10616 23440 10668
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 27528 10659 27580 10668
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 28816 10727 28868 10736
rect 28816 10693 28825 10727
rect 28825 10693 28859 10727
rect 28859 10693 28868 10727
rect 28816 10684 28868 10693
rect 29920 10616 29972 10668
rect 30656 10616 30708 10668
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 23940 10548 23992 10600
rect 24492 10548 24544 10600
rect 26608 10548 26660 10600
rect 27068 10548 27120 10600
rect 23572 10480 23624 10532
rect 29552 10591 29604 10600
rect 29552 10557 29561 10591
rect 29561 10557 29595 10591
rect 29595 10557 29604 10591
rect 29552 10548 29604 10557
rect 29828 10548 29880 10600
rect 30472 10591 30524 10600
rect 30472 10557 30481 10591
rect 30481 10557 30515 10591
rect 30515 10557 30524 10591
rect 30472 10548 30524 10557
rect 30840 10548 30892 10600
rect 32312 10548 32364 10600
rect 32404 10591 32456 10600
rect 32404 10557 32413 10591
rect 32413 10557 32447 10591
rect 32447 10557 32456 10591
rect 32404 10548 32456 10557
rect 33232 10684 33284 10736
rect 33508 10684 33560 10736
rect 35256 10684 35308 10736
rect 35624 10659 35676 10668
rect 35624 10625 35633 10659
rect 35633 10625 35667 10659
rect 35667 10625 35676 10659
rect 35624 10616 35676 10625
rect 35716 10616 35768 10668
rect 22100 10412 22152 10464
rect 23756 10455 23808 10464
rect 23756 10421 23765 10455
rect 23765 10421 23799 10455
rect 23799 10421 23808 10455
rect 23756 10412 23808 10421
rect 24768 10412 24820 10464
rect 35256 10548 35308 10600
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 36820 10795 36872 10804
rect 36820 10761 36829 10795
rect 36829 10761 36863 10795
rect 36863 10761 36872 10795
rect 36820 10752 36872 10761
rect 38568 10684 38620 10736
rect 49240 10684 49292 10736
rect 38936 10616 38988 10668
rect 46940 10616 46992 10668
rect 36360 10591 36412 10600
rect 36360 10557 36369 10591
rect 36369 10557 36403 10591
rect 36403 10557 36412 10591
rect 36360 10548 36412 10557
rect 36544 10548 36596 10600
rect 36912 10548 36964 10600
rect 30840 10412 30892 10464
rect 31760 10412 31812 10464
rect 31944 10455 31996 10464
rect 31944 10421 31953 10455
rect 31953 10421 31987 10455
rect 31987 10421 31996 10455
rect 31944 10412 31996 10421
rect 32864 10412 32916 10464
rect 36636 10480 36688 10532
rect 37556 10480 37608 10532
rect 47124 10480 47176 10532
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 15016 10208 15068 10260
rect 4804 10140 4856 10192
rect 12532 10140 12584 10192
rect 14740 10140 14792 10192
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 16120 10208 16172 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 18328 10208 18380 10260
rect 20168 10208 20220 10260
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 14280 10004 14332 10056
rect 14648 10004 14700 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 14188 9936 14240 9988
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 13084 9868 13136 9920
rect 13912 9868 13964 9920
rect 17684 10140 17736 10192
rect 16304 10072 16356 10124
rect 17868 10072 17920 10124
rect 18420 10072 18472 10124
rect 18604 10115 18656 10124
rect 18604 10081 18613 10115
rect 18613 10081 18647 10115
rect 18647 10081 18656 10115
rect 18604 10072 18656 10081
rect 19432 10072 19484 10124
rect 19616 10072 19668 10124
rect 16212 10004 16264 10056
rect 23664 10208 23716 10260
rect 24492 10208 24544 10260
rect 26332 10208 26384 10260
rect 27436 10208 27488 10260
rect 29092 10208 29144 10260
rect 29828 10208 29880 10260
rect 31392 10208 31444 10260
rect 20444 10072 20496 10124
rect 20720 10072 20772 10124
rect 21088 10072 21140 10124
rect 23848 10072 23900 10124
rect 26608 10140 26660 10192
rect 26700 10183 26752 10192
rect 26700 10149 26709 10183
rect 26709 10149 26743 10183
rect 26743 10149 26752 10183
rect 26700 10140 26752 10149
rect 29276 10183 29328 10192
rect 29276 10149 29285 10183
rect 29285 10149 29319 10183
rect 29319 10149 29328 10183
rect 29276 10140 29328 10149
rect 26884 10072 26936 10124
rect 29552 10072 29604 10124
rect 30656 10072 30708 10124
rect 30840 10072 30892 10124
rect 32588 10208 32640 10260
rect 35716 10208 35768 10260
rect 36636 10251 36688 10260
rect 36636 10217 36645 10251
rect 36645 10217 36679 10251
rect 36679 10217 36688 10251
rect 36636 10208 36688 10217
rect 36912 10251 36964 10260
rect 36912 10217 36921 10251
rect 36921 10217 36955 10251
rect 36955 10217 36964 10251
rect 36912 10208 36964 10217
rect 32220 10140 32272 10192
rect 32128 10115 32180 10124
rect 32128 10081 32137 10115
rect 32137 10081 32171 10115
rect 32171 10081 32180 10115
rect 32128 10072 32180 10081
rect 32588 10072 32640 10124
rect 34704 10072 34756 10124
rect 35624 10072 35676 10124
rect 35716 10072 35768 10124
rect 16764 9936 16816 9988
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 24032 10004 24084 10056
rect 32772 10004 32824 10056
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 36544 10004 36596 10056
rect 38936 10004 38988 10056
rect 49148 10115 49200 10124
rect 49148 10081 49157 10115
rect 49157 10081 49191 10115
rect 49191 10081 49200 10115
rect 49148 10072 49200 10081
rect 45836 10004 45888 10056
rect 46112 10047 46164 10056
rect 46112 10013 46121 10047
rect 46121 10013 46155 10047
rect 46155 10013 46164 10047
rect 46112 10004 46164 10013
rect 46572 10004 46624 10056
rect 16580 9911 16632 9920
rect 16580 9877 16589 9911
rect 16589 9877 16623 9911
rect 16623 9877 16632 9911
rect 16580 9868 16632 9877
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17316 9911 17368 9920
rect 17316 9877 17325 9911
rect 17325 9877 17359 9911
rect 17359 9877 17368 9911
rect 17316 9868 17368 9877
rect 22560 9936 22612 9988
rect 23388 9936 23440 9988
rect 24400 9936 24452 9988
rect 25596 9936 25648 9988
rect 25780 9936 25832 9988
rect 27344 9936 27396 9988
rect 23572 9868 23624 9920
rect 23940 9868 23992 9920
rect 26700 9868 26752 9920
rect 30840 9936 30892 9988
rect 31852 9979 31904 9988
rect 31852 9945 31861 9979
rect 31861 9945 31895 9979
rect 31895 9945 31904 9979
rect 31852 9936 31904 9945
rect 31944 9936 31996 9988
rect 28908 9868 28960 9920
rect 30104 9868 30156 9920
rect 33232 9868 33284 9920
rect 37464 9936 37516 9988
rect 44364 9979 44416 9988
rect 44364 9945 44373 9979
rect 44373 9945 44407 9979
rect 44407 9945 44416 9979
rect 44364 9936 44416 9945
rect 46756 9936 46808 9988
rect 47308 9979 47360 9988
rect 47308 9945 47317 9979
rect 47317 9945 47351 9979
rect 47351 9945 47360 9979
rect 47308 9936 47360 9945
rect 38384 9911 38436 9920
rect 38384 9877 38393 9911
rect 38393 9877 38427 9911
rect 38427 9877 38436 9911
rect 38384 9868 38436 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 1308 9664 1360 9716
rect 2412 9664 2464 9716
rect 14740 9664 14792 9716
rect 16580 9664 16632 9716
rect 19984 9664 20036 9716
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 22284 9707 22336 9716
rect 22284 9673 22293 9707
rect 22293 9673 22327 9707
rect 22327 9673 22336 9707
rect 22284 9664 22336 9673
rect 22560 9664 22612 9716
rect 24584 9664 24636 9716
rect 28816 9664 28868 9716
rect 28908 9664 28960 9716
rect 30656 9664 30708 9716
rect 30840 9664 30892 9716
rect 31484 9664 31536 9716
rect 12624 9596 12676 9648
rect 13728 9596 13780 9648
rect 15108 9596 15160 9648
rect 15200 9596 15252 9648
rect 1308 9528 1360 9580
rect 12348 9528 12400 9580
rect 16028 9596 16080 9648
rect 16212 9596 16264 9648
rect 16672 9596 16724 9648
rect 16856 9639 16908 9648
rect 16856 9605 16865 9639
rect 16865 9605 16899 9639
rect 16899 9605 16908 9639
rect 16856 9596 16908 9605
rect 18328 9596 18380 9648
rect 19524 9596 19576 9648
rect 20352 9596 20404 9648
rect 21272 9596 21324 9648
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 11060 9460 11112 9512
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 18604 9503 18656 9512
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 18880 9503 18932 9512
rect 18880 9469 18889 9503
rect 18889 9469 18923 9503
rect 18923 9469 18932 9503
rect 18880 9460 18932 9469
rect 24400 9596 24452 9648
rect 24676 9596 24728 9648
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 27344 9596 27396 9648
rect 30104 9596 30156 9648
rect 31668 9596 31720 9648
rect 33508 9664 33560 9716
rect 34428 9664 34480 9716
rect 35624 9707 35676 9716
rect 35624 9673 35633 9707
rect 35633 9673 35667 9707
rect 35667 9673 35676 9707
rect 35624 9664 35676 9673
rect 36544 9664 36596 9716
rect 38384 9664 38436 9716
rect 46940 9664 46992 9716
rect 32128 9596 32180 9648
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 17316 9392 17368 9444
rect 14924 9324 14976 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 16304 9324 16356 9376
rect 18420 9324 18472 9376
rect 21548 9367 21600 9376
rect 21548 9333 21557 9367
rect 21557 9333 21591 9367
rect 21591 9333 21600 9367
rect 21548 9324 21600 9333
rect 21824 9367 21876 9376
rect 21824 9333 21833 9367
rect 21833 9333 21867 9367
rect 21867 9333 21876 9367
rect 21824 9324 21876 9333
rect 23756 9324 23808 9376
rect 24492 9460 24544 9512
rect 25964 9503 26016 9512
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 25688 9392 25740 9444
rect 31116 9528 31168 9580
rect 31760 9528 31812 9580
rect 34704 9596 34756 9648
rect 49240 9596 49292 9648
rect 47216 9528 47268 9580
rect 27160 9460 27212 9512
rect 29276 9503 29328 9512
rect 29276 9469 29285 9503
rect 29285 9469 29319 9503
rect 29319 9469 29328 9503
rect 29276 9460 29328 9469
rect 29552 9460 29604 9512
rect 30012 9503 30064 9512
rect 25872 9324 25924 9376
rect 29460 9392 29512 9444
rect 30012 9469 30021 9503
rect 30021 9469 30055 9503
rect 30055 9469 30064 9503
rect 30012 9460 30064 9469
rect 30104 9460 30156 9512
rect 31852 9460 31904 9512
rect 34244 9460 34296 9512
rect 36084 9460 36136 9512
rect 32588 9392 32640 9444
rect 30472 9324 30524 9376
rect 31116 9324 31168 9376
rect 35164 9324 35216 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 2136 9052 2188 9104
rect 15384 9052 15436 9104
rect 15752 9120 15804 9172
rect 17132 9120 17184 9172
rect 17868 9163 17920 9172
rect 17868 9129 17889 9163
rect 17889 9129 17920 9163
rect 17868 9120 17920 9129
rect 19524 9120 19576 9172
rect 22100 9120 22152 9172
rect 16764 9052 16816 9104
rect 1216 8916 1268 8968
rect 3148 8984 3200 9036
rect 13360 8984 13412 9036
rect 15108 8984 15160 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 16488 8984 16540 9036
rect 18880 8984 18932 9036
rect 19432 8984 19484 9036
rect 1308 8848 1360 8900
rect 13544 8916 13596 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 21456 8916 21508 8968
rect 22008 8916 22060 8968
rect 2596 8780 2648 8832
rect 3148 8780 3200 8832
rect 13728 8848 13780 8900
rect 13820 8780 13872 8832
rect 14464 8823 14516 8832
rect 14464 8789 14473 8823
rect 14473 8789 14507 8823
rect 14507 8789 14516 8823
rect 14464 8780 14516 8789
rect 15292 8780 15344 8832
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 17408 8848 17460 8900
rect 18420 8848 18472 8900
rect 20444 8848 20496 8900
rect 24584 9120 24636 9172
rect 25964 9120 26016 9172
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 24032 9027 24084 9036
rect 24032 8993 24041 9027
rect 24041 8993 24075 9027
rect 24075 8993 24084 9027
rect 24032 8984 24084 8993
rect 24400 8984 24452 9036
rect 25596 8984 25648 9036
rect 30012 9052 30064 9104
rect 33508 9120 33560 9172
rect 36360 9120 36412 9172
rect 37096 9120 37148 9172
rect 39948 9052 40000 9104
rect 24400 8848 24452 8900
rect 22192 8780 22244 8832
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 27804 8823 27856 8832
rect 27804 8789 27813 8823
rect 27813 8789 27847 8823
rect 27847 8789 27856 8823
rect 31760 8984 31812 9036
rect 32128 8984 32180 9036
rect 30656 8916 30708 8968
rect 31116 8916 31168 8968
rect 32588 8916 32640 8968
rect 33600 9027 33652 9036
rect 33600 8993 33609 9027
rect 33609 8993 33643 9027
rect 33643 8993 33652 9027
rect 33600 8984 33652 8993
rect 34060 8984 34112 9036
rect 35164 8984 35216 9036
rect 34244 8916 34296 8968
rect 34520 8916 34572 8968
rect 49332 8984 49384 9036
rect 27804 8780 27856 8789
rect 30656 8780 30708 8832
rect 34060 8848 34112 8900
rect 34152 8848 34204 8900
rect 37096 8848 37148 8900
rect 47032 8916 47084 8968
rect 47584 8848 47636 8900
rect 31944 8780 31996 8832
rect 33692 8823 33744 8832
rect 33692 8789 33701 8823
rect 33701 8789 33735 8823
rect 33735 8789 33744 8823
rect 33692 8780 33744 8789
rect 34612 8780 34664 8832
rect 35624 8823 35676 8832
rect 35624 8789 35633 8823
rect 35633 8789 35667 8823
rect 35667 8789 35676 8823
rect 35624 8780 35676 8789
rect 39764 8780 39816 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 12716 8576 12768 8628
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 15200 8576 15252 8628
rect 13912 8551 13964 8560
rect 13912 8517 13921 8551
rect 13921 8517 13955 8551
rect 13955 8517 13964 8551
rect 13912 8508 13964 8517
rect 15292 8508 15344 8560
rect 17408 8576 17460 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 19892 8576 19944 8628
rect 16764 8508 16816 8560
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 18420 8508 18472 8560
rect 20444 8508 20496 8560
rect 15200 8440 15252 8492
rect 16488 8440 16540 8492
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 15108 8372 15160 8424
rect 17776 8372 17828 8424
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 22008 8440 22060 8492
rect 24400 8576 24452 8628
rect 31116 8576 31168 8628
rect 33876 8576 33928 8628
rect 34060 8619 34112 8628
rect 34060 8585 34069 8619
rect 34069 8585 34103 8619
rect 34103 8585 34112 8619
rect 34060 8576 34112 8585
rect 34244 8576 34296 8628
rect 41420 8576 41472 8628
rect 29092 8551 29144 8560
rect 29092 8517 29101 8551
rect 29101 8517 29135 8551
rect 29135 8517 29144 8551
rect 29092 8508 29144 8517
rect 30656 8508 30708 8560
rect 24032 8440 24084 8492
rect 31944 8508 31996 8560
rect 32588 8508 32640 8560
rect 34704 8551 34756 8560
rect 34704 8517 34713 8551
rect 34713 8517 34747 8551
rect 34747 8517 34756 8551
rect 34704 8508 34756 8517
rect 35624 8508 35676 8560
rect 22100 8372 22152 8424
rect 28816 8415 28868 8424
rect 28816 8381 28825 8415
rect 28825 8381 28859 8415
rect 28859 8381 28868 8415
rect 28816 8372 28868 8381
rect 29184 8372 29236 8424
rect 31760 8440 31812 8492
rect 32036 8440 32088 8492
rect 32128 8440 32180 8492
rect 31300 8415 31352 8424
rect 31300 8381 31309 8415
rect 31309 8381 31343 8415
rect 31343 8381 31352 8415
rect 31300 8372 31352 8381
rect 32220 8372 32272 8424
rect 32680 8372 32732 8424
rect 32956 8372 33008 8424
rect 33876 8372 33928 8424
rect 36452 8372 36504 8424
rect 37464 8483 37516 8492
rect 37464 8449 37473 8483
rect 37473 8449 37507 8483
rect 37507 8449 37516 8483
rect 37464 8440 37516 8449
rect 39764 8508 39816 8560
rect 47860 8508 47912 8560
rect 49148 8551 49200 8560
rect 49148 8517 49157 8551
rect 49157 8517 49191 8551
rect 49191 8517 49200 8551
rect 49148 8508 49200 8517
rect 40316 8483 40368 8492
rect 40316 8449 40325 8483
rect 40325 8449 40359 8483
rect 40359 8449 40368 8483
rect 40316 8440 40368 8449
rect 45836 8483 45888 8492
rect 45836 8449 45845 8483
rect 45845 8449 45879 8483
rect 45879 8449 45888 8483
rect 45836 8440 45888 8449
rect 46756 8440 46808 8492
rect 38752 8372 38804 8424
rect 22468 8304 22520 8356
rect 31852 8304 31904 8356
rect 33600 8304 33652 8356
rect 38936 8304 38988 8356
rect 44916 8304 44968 8356
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 47676 8304 47728 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 1308 8032 1360 8084
rect 2412 8032 2464 8084
rect 18512 8032 18564 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 21916 8032 21968 8084
rect 30564 8032 30616 8084
rect 34152 8032 34204 8084
rect 18880 7964 18932 8016
rect 39028 7964 39080 8016
rect 16764 7939 16816 7948
rect 16764 7905 16773 7939
rect 16773 7905 16807 7939
rect 16807 7905 16816 7939
rect 16764 7896 16816 7905
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 18604 7896 18656 7948
rect 19892 7896 19944 7948
rect 23664 7896 23716 7948
rect 29920 7939 29972 7948
rect 29920 7905 29929 7939
rect 29929 7905 29963 7939
rect 29963 7905 29972 7939
rect 29920 7896 29972 7905
rect 32220 7896 32272 7948
rect 34796 7896 34848 7948
rect 49240 7896 49292 7948
rect 1308 7828 1360 7880
rect 2688 7828 2740 7880
rect 12440 7828 12492 7880
rect 14924 7828 14976 7880
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 13728 7760 13780 7812
rect 16396 7760 16448 7812
rect 19616 7760 19668 7812
rect 20444 7760 20496 7812
rect 20996 7760 21048 7812
rect 21456 7828 21508 7880
rect 22192 7828 22244 7880
rect 30564 7828 30616 7880
rect 32772 7828 32824 7880
rect 38752 7871 38804 7880
rect 38752 7837 38761 7871
rect 38761 7837 38795 7871
rect 38795 7837 38804 7871
rect 38752 7828 38804 7837
rect 47124 7828 47176 7880
rect 30472 7803 30524 7812
rect 30472 7769 30481 7803
rect 30481 7769 30515 7803
rect 30515 7769 30524 7803
rect 30472 7760 30524 7769
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 21640 7735 21692 7744
rect 21640 7701 21649 7735
rect 21649 7701 21683 7735
rect 21683 7701 21692 7735
rect 21640 7692 21692 7701
rect 22376 7692 22428 7744
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 25688 7692 25740 7744
rect 27252 7692 27304 7744
rect 41328 7760 41380 7812
rect 30656 7735 30708 7744
rect 30656 7701 30665 7735
rect 30665 7701 30699 7735
rect 30699 7701 30708 7735
rect 30656 7692 30708 7701
rect 31392 7735 31444 7744
rect 31392 7701 31401 7735
rect 31401 7701 31435 7735
rect 31435 7701 31444 7735
rect 31392 7692 31444 7701
rect 32588 7735 32640 7744
rect 32588 7701 32597 7735
rect 32597 7701 32631 7735
rect 32631 7701 32640 7735
rect 32588 7692 32640 7701
rect 38660 7692 38712 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 17868 7488 17920 7540
rect 18420 7488 18472 7540
rect 20444 7488 20496 7540
rect 20628 7488 20680 7540
rect 22284 7488 22336 7540
rect 31116 7531 31168 7540
rect 31116 7497 31125 7531
rect 31125 7497 31159 7531
rect 31159 7497 31168 7531
rect 31116 7488 31168 7497
rect 31392 7488 31444 7540
rect 38660 7488 38712 7540
rect 47308 7488 47360 7540
rect 31944 7463 31996 7472
rect 31944 7429 31953 7463
rect 31953 7429 31987 7463
rect 31987 7429 31996 7463
rect 31944 7420 31996 7429
rect 1308 7352 1360 7404
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 27620 7352 27672 7404
rect 44916 7463 44968 7472
rect 44916 7429 44925 7463
rect 44925 7429 44959 7463
rect 44959 7429 44968 7463
rect 44916 7420 44968 7429
rect 49332 7420 49384 7472
rect 33324 7352 33376 7404
rect 46940 7352 46992 7404
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 30472 7284 30524 7336
rect 31300 7284 31352 7336
rect 38476 7284 38528 7336
rect 18788 7216 18840 7268
rect 20720 7216 20772 7268
rect 21640 7216 21692 7268
rect 22652 7216 22704 7268
rect 32588 7216 32640 7268
rect 37280 7216 37332 7268
rect 21456 7148 21508 7200
rect 22008 7148 22060 7200
rect 37924 7191 37976 7200
rect 37924 7157 37933 7191
rect 37933 7157 37967 7191
rect 37967 7157 37976 7191
rect 37924 7148 37976 7157
rect 47768 7216 47820 7268
rect 45836 7148 45888 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 37924 6876 37976 6928
rect 46940 6876 46992 6928
rect 15660 6808 15712 6860
rect 22376 6808 22428 6860
rect 49148 6851 49200 6860
rect 49148 6817 49157 6851
rect 49157 6817 49191 6851
rect 49191 6817 49200 6851
rect 49148 6808 49200 6817
rect 1308 6740 1360 6792
rect 15936 6740 15988 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 41328 6740 41380 6792
rect 47860 6740 47912 6792
rect 1216 6672 1268 6724
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 10600 6672 10652 6724
rect 48688 6672 48740 6724
rect 19248 6604 19300 6656
rect 21732 6604 21784 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 1216 6400 1268 6452
rect 27528 6332 27580 6384
rect 36820 6332 36872 6384
rect 41420 6332 41472 6384
rect 49424 6332 49476 6384
rect 1308 6264 1360 6316
rect 1768 6264 1820 6316
rect 27804 6264 27856 6316
rect 30748 6264 30800 6316
rect 47584 6264 47636 6316
rect 11152 6196 11204 6248
rect 14464 6196 14516 6248
rect 18328 6196 18380 6248
rect 26976 6196 27028 6248
rect 37740 6196 37792 6248
rect 4068 6128 4120 6180
rect 23940 6128 23992 6180
rect 25688 6128 25740 6180
rect 36452 6128 36504 6180
rect 47032 6128 47084 6180
rect 19432 6060 19484 6112
rect 37648 6103 37700 6112
rect 37648 6069 37657 6103
rect 37657 6069 37691 6103
rect 37691 6069 37700 6103
rect 37648 6060 37700 6069
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 2596 5856 2648 5908
rect 37648 5856 37700 5908
rect 47216 5856 47268 5908
rect 1308 5652 1360 5704
rect 49240 5720 49292 5772
rect 2780 5652 2832 5704
rect 39948 5652 40000 5704
rect 47676 5652 47728 5704
rect 16304 5584 16356 5636
rect 45744 5584 45796 5636
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 37280 5355 37332 5364
rect 37280 5321 37289 5355
rect 37289 5321 37323 5355
rect 37323 5321 37332 5355
rect 37280 5312 37332 5321
rect 38476 5287 38528 5296
rect 38476 5253 38485 5287
rect 38485 5253 38519 5287
rect 38519 5253 38528 5287
rect 38476 5244 38528 5253
rect 49148 5287 49200 5296
rect 49148 5253 49157 5287
rect 49157 5253 49191 5287
rect 49191 5253 49200 5287
rect 49148 5244 49200 5253
rect 12808 5176 12860 5228
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 28356 5176 28408 5228
rect 33324 5176 33376 5228
rect 45836 5219 45888 5228
rect 45836 5185 45845 5219
rect 45845 5185 45879 5219
rect 45879 5185 45888 5219
rect 45836 5176 45888 5185
rect 47768 5176 47820 5228
rect 1308 5108 1360 5160
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 48320 5108 48372 5160
rect 41328 5040 41380 5092
rect 4436 4972 4488 5024
rect 15660 4972 15712 5024
rect 20628 4972 20680 5024
rect 37832 5015 37884 5024
rect 37832 4981 37841 5015
rect 37841 4981 37875 5015
rect 37875 4981 37884 5015
rect 37832 4972 37884 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 1308 4768 1360 4820
rect 6828 4768 6880 4820
rect 20720 4768 20772 4820
rect 36820 4811 36872 4820
rect 36820 4777 36829 4811
rect 36829 4777 36863 4811
rect 36863 4777 36872 4811
rect 36820 4768 36872 4777
rect 37832 4768 37884 4820
rect 47124 4768 47176 4820
rect 4068 4700 4120 4752
rect 26148 4700 26200 4752
rect 38936 4700 38988 4752
rect 19248 4632 19300 4684
rect 21732 4632 21784 4684
rect 1308 4564 1360 4616
rect 19984 4564 20036 4616
rect 22928 4632 22980 4684
rect 23204 4632 23256 4684
rect 37004 4632 37056 4684
rect 49424 4632 49476 4684
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 19064 4496 19116 4548
rect 23572 4564 23624 4616
rect 32772 4564 32824 4616
rect 36820 4564 36872 4616
rect 37740 4564 37792 4616
rect 47308 4564 47360 4616
rect 21272 4428 21324 4480
rect 21364 4428 21416 4480
rect 21824 4428 21876 4480
rect 39948 4496 40000 4548
rect 25872 4428 25924 4480
rect 37372 4471 37424 4480
rect 37372 4437 37381 4471
rect 37381 4437 37415 4471
rect 37415 4437 37424 4471
rect 37372 4428 37424 4437
rect 47676 4496 47728 4548
rect 49792 4428 49844 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1768 4224 1820 4276
rect 4804 4224 4856 4276
rect 13728 4224 13780 4276
rect 21364 4224 21416 4276
rect 37372 4224 37424 4276
rect 45652 4224 45704 4276
rect 1400 4156 1452 4208
rect 1308 4088 1360 4140
rect 22100 4156 22152 4208
rect 4436 3952 4488 4004
rect 16580 3952 16632 4004
rect 18328 3952 18380 4004
rect 22928 4131 22980 4140
rect 22928 4097 22972 4131
rect 22972 4097 22980 4131
rect 22928 4088 22980 4097
rect 23204 4088 23256 4140
rect 25872 4199 25924 4208
rect 25872 4165 25881 4199
rect 25881 4165 25915 4199
rect 25915 4165 25924 4199
rect 25872 4156 25924 4165
rect 27620 4088 27672 4140
rect 45836 4131 45888 4140
rect 45836 4097 45845 4131
rect 45845 4097 45879 4131
rect 45879 4097 45888 4131
rect 45836 4088 45888 4097
rect 46940 4088 46992 4140
rect 49332 4088 49384 4140
rect 23296 4020 23348 4072
rect 24860 4063 24912 4072
rect 24860 4029 24869 4063
rect 24869 4029 24903 4063
rect 24903 4029 24912 4063
rect 24860 4020 24912 4029
rect 25780 4020 25832 4072
rect 6828 3884 6880 3936
rect 22836 3884 22888 3936
rect 32864 4020 32916 4072
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 27528 3884 27580 3936
rect 47676 3927 47728 3936
rect 47676 3893 47685 3927
rect 47685 3893 47719 3927
rect 47719 3893 47728 3927
rect 47676 3884 47728 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 22008 3680 22060 3732
rect 23572 3723 23624 3732
rect 23572 3689 23581 3723
rect 23581 3689 23615 3723
rect 23615 3689 23624 3723
rect 23572 3680 23624 3689
rect 25964 3680 26016 3732
rect 41328 3680 41380 3732
rect 7472 3612 7524 3664
rect 2688 3544 2740 3596
rect 3332 3544 3384 3596
rect 13728 3544 13780 3596
rect 1308 3408 1360 3460
rect 10324 3476 10376 3528
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 14096 3408 14148 3460
rect 10692 3340 10744 3392
rect 33416 3612 33468 3664
rect 22836 3544 22888 3596
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 24124 3476 24176 3528
rect 29000 3476 29052 3528
rect 33324 3476 33376 3528
rect 39212 3476 39264 3528
rect 45836 3476 45888 3528
rect 49148 3587 49200 3596
rect 49148 3553 49157 3587
rect 49157 3553 49191 3587
rect 49191 3553 49200 3587
rect 49148 3544 49200 3553
rect 47032 3476 47084 3528
rect 19340 3408 19392 3460
rect 21364 3408 21416 3460
rect 22008 3408 22060 3460
rect 36452 3451 36504 3460
rect 36452 3417 36461 3451
rect 36461 3417 36495 3451
rect 36495 3417 36504 3451
rect 36452 3408 36504 3417
rect 45560 3451 45612 3460
rect 45560 3417 45569 3451
rect 45569 3417 45603 3451
rect 45603 3417 45612 3451
rect 45560 3408 45612 3417
rect 48688 3408 48740 3460
rect 22744 3383 22796 3392
rect 22744 3349 22753 3383
rect 22753 3349 22787 3383
rect 22787 3349 22796 3383
rect 22744 3340 22796 3349
rect 26332 3340 26384 3392
rect 29644 3340 29696 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 1308 3136 1360 3188
rect 10324 3179 10376 3188
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 1308 3000 1360 3052
rect 9588 3000 9640 3052
rect 9772 3000 9824 3052
rect 15200 3136 15252 3188
rect 19340 3136 19392 3188
rect 17868 3068 17920 3120
rect 19064 3000 19116 3052
rect 24584 3136 24636 3188
rect 22100 3068 22152 3120
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 24032 3068 24084 3120
rect 26332 3068 26384 3120
rect 26148 3000 26200 3052
rect 37740 3136 37792 3188
rect 29644 3068 29696 3120
rect 49240 3068 49292 3120
rect 28816 3000 28868 3052
rect 39948 3000 40000 3052
rect 45744 3000 45796 3052
rect 47216 3000 47268 3052
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 20996 2932 21048 2984
rect 1768 2907 1820 2916
rect 1768 2873 1777 2907
rect 1777 2873 1811 2907
rect 1811 2873 1820 2907
rect 1768 2864 1820 2873
rect 22100 2864 22152 2916
rect 22192 2907 22244 2916
rect 22192 2873 22201 2907
rect 22201 2873 22235 2907
rect 22235 2873 22244 2907
rect 22192 2864 22244 2873
rect 22744 2864 22796 2916
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 29644 2932 29696 2984
rect 30656 2932 30708 2984
rect 46756 2932 46808 2984
rect 46848 2975 46900 2984
rect 46848 2941 46857 2975
rect 46857 2941 46891 2975
rect 46891 2941 46900 2975
rect 46848 2932 46900 2941
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 17408 2796 17460 2805
rect 21364 2796 21416 2848
rect 23296 2839 23348 2848
rect 23296 2805 23305 2839
rect 23305 2805 23339 2839
rect 23339 2805 23348 2839
rect 23296 2796 23348 2805
rect 27528 2907 27580 2916
rect 27528 2873 27537 2907
rect 27537 2873 27571 2907
rect 27571 2873 27580 2907
rect 27528 2864 27580 2873
rect 27160 2796 27212 2848
rect 38292 2864 38344 2916
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 9772 2524 9824 2576
rect 24032 2635 24084 2644
rect 24032 2601 24041 2635
rect 24041 2601 24075 2635
rect 24075 2601 24084 2635
rect 24032 2592 24084 2601
rect 26332 2635 26384 2644
rect 26332 2601 26341 2635
rect 26341 2601 26375 2635
rect 26375 2601 26384 2635
rect 26332 2592 26384 2601
rect 27620 2592 27672 2644
rect 29000 2635 29052 2644
rect 29000 2601 29009 2635
rect 29009 2601 29043 2635
rect 29043 2601 29052 2635
rect 29000 2592 29052 2601
rect 32864 2592 32916 2644
rect 22468 2524 22520 2576
rect 32772 2524 32824 2576
rect 34336 2524 34388 2576
rect 1308 2388 1360 2440
rect 2780 2388 2832 2440
rect 1216 2320 1268 2372
rect 2320 2320 2372 2372
rect 1308 2252 1360 2304
rect 12256 2456 12308 2508
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 14096 2388 14148 2440
rect 17408 2388 17460 2440
rect 11704 2320 11756 2372
rect 13820 2320 13872 2372
rect 15936 2320 15988 2372
rect 14740 2252 14792 2304
rect 19984 2456 20036 2508
rect 20168 2456 20220 2508
rect 22284 2456 22336 2508
rect 24400 2456 24452 2508
rect 26516 2456 26568 2508
rect 37740 2499 37792 2508
rect 37740 2465 37749 2499
rect 37749 2465 37783 2499
rect 37783 2465 37792 2499
rect 37740 2456 37792 2465
rect 41328 2456 41380 2508
rect 49148 2499 49200 2508
rect 49148 2465 49157 2499
rect 49157 2465 49191 2499
rect 49191 2465 49200 2499
rect 49148 2456 49200 2465
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 22100 2388 22152 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 29000 2388 29052 2440
rect 30748 2388 30800 2440
rect 33140 2431 33192 2440
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 34980 2388 35032 2440
rect 38292 2388 38344 2440
rect 45652 2388 45704 2440
rect 47124 2388 47176 2440
rect 48504 2320 48556 2372
rect 37096 2295 37148 2304
rect 37096 2261 37105 2295
rect 37105 2261 37139 2295
rect 37139 2261 37148 2295
rect 37096 2252 37148 2261
rect 43444 2252 43496 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26330 2926 27000
rect 2870 26302 3372 26330
rect 2870 26200 2926 26302
rect 1596 22778 1624 26200
rect 1768 23044 1820 23050
rect 1768 22986 1820 22992
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1032 21956 1084 21962
rect 1032 21898 1084 21904
rect 1044 20777 1072 21898
rect 1780 21593 1808 22986
rect 2240 22234 2268 26200
rect 3146 25664 3202 25673
rect 3146 25599 3202 25608
rect 3160 25498 3188 25599
rect 3148 25492 3200 25498
rect 3148 25434 3200 25440
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2778 24440 2834 24449
rect 2950 24443 3258 24452
rect 2778 24375 2834 24384
rect 2792 23526 2820 24375
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2962 23216 3018 23225
rect 2962 23151 3018 23160
rect 2780 22500 2832 22506
rect 2780 22442 2832 22448
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 1766 21584 1822 21593
rect 1766 21519 1822 21528
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1030 20768 1086 20777
rect 1030 20703 1086 20712
rect 1308 20528 1360 20534
rect 1308 20470 1360 20476
rect 1320 20369 1348 20470
rect 1306 20360 1362 20369
rect 1306 20295 1362 20304
rect 1780 19961 1808 21422
rect 2792 21185 2820 22442
rect 2976 22438 3004 23151
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3238 21992 3294 22001
rect 3238 21927 3240 21936
rect 3292 21927 3294 21936
rect 3240 21898 3292 21904
rect 3344 21622 3372 26302
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26200 4858 27000
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26330 8078 27000
rect 7852 26302 8078 26330
rect 3528 24274 3556 26200
rect 3790 25256 3846 25265
rect 3790 25191 3846 25200
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3514 24032 3570 24041
rect 3514 23967 3570 23976
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2778 21176 2834 21185
rect 2950 21179 3258 21188
rect 2778 21111 2834 21120
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 1766 19952 1822 19961
rect 1766 19887 1822 19896
rect 1492 19780 1544 19786
rect 1492 19722 1544 19728
rect 1504 18737 1532 19722
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1490 18728 1546 18737
rect 1400 18692 1452 18698
rect 1490 18663 1546 18672
rect 1400 18634 1452 18640
rect 1412 17921 1440 18634
rect 1780 18329 1808 19314
rect 2792 19145 2820 20266
rect 2884 19553 2912 20946
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19854 3372 20266
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 2870 19544 2926 19553
rect 2870 19479 2926 19488
rect 3436 19446 3464 22714
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3528 18834 3556 23967
rect 3608 23044 3660 23050
rect 3608 22986 3660 22992
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3620 18426 3648 22986
rect 3804 21350 3832 25191
rect 3882 24848 3938 24857
rect 3882 24783 3884 24792
rect 3936 24783 3938 24792
rect 3884 24754 3936 24760
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3896 19310 3924 24142
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 3974 23624 4030 23633
rect 3974 23559 3976 23568
rect 4028 23559 4030 23568
rect 3976 23530 4028 23536
rect 3974 22808 4030 22817
rect 3974 22743 4030 22752
rect 3988 22166 4016 22743
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 1766 18320 1822 18329
rect 4080 18290 4108 23666
rect 4172 23662 4200 26200
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4632 23866 4660 24142
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4724 23322 4752 23666
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4252 22228 4304 22234
rect 4252 22170 4304 22176
rect 4158 22128 4214 22137
rect 4158 22063 4214 22072
rect 4172 21010 4200 22063
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 18358 4200 20198
rect 4264 19922 4292 22170
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 1766 18255 1822 18264
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 1032 17604 1084 17610
rect 1032 17546 1084 17552
rect 940 17128 992 17134
rect 1044 17105 1072 17546
rect 1780 17513 1808 18158
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 1766 17504 1822 17513
rect 1766 17439 1822 17448
rect 3332 17264 3384 17270
rect 3332 17206 3384 17212
rect 940 17070 992 17076
rect 1030 17096 1086 17105
rect 952 16697 980 17070
rect 1030 17031 1086 17040
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 938 16688 994 16697
rect 938 16623 994 16632
rect 3344 16590 3372 17206
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 1032 16516 1084 16522
rect 1032 16458 1084 16464
rect 1044 16289 1072 16458
rect 1030 16280 1086 16289
rect 1030 16215 1086 16224
rect 4264 16114 4292 18158
rect 4356 17202 4384 18634
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4448 16658 4476 23054
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4632 21554 4660 22918
rect 4816 22710 4844 26200
rect 5460 23662 5488 26200
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5816 23588 5868 23594
rect 5816 23530 5868 23536
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 4816 20058 4844 20402
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 5276 19990 5304 20402
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5368 19854 5396 22918
rect 5644 21962 5672 23258
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5354 18864 5410 18873
rect 5354 18799 5410 18808
rect 5368 18766 5396 18799
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5644 18358 5672 21422
rect 5736 19922 5764 23462
rect 5828 21486 5856 23530
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 5920 20398 5948 24754
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 6012 22642 6040 23462
rect 6104 23186 6132 26200
rect 6748 24274 6776 26200
rect 6736 24268 6788 24274
rect 6736 24210 6788 24216
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6656 23118 6684 24006
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 7116 22710 7144 24142
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 6368 22500 6420 22506
rect 6368 22442 6420 22448
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6012 21010 6040 22374
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 6380 20466 6408 22442
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 21690 6776 21830
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6550 21584 6606 21593
rect 6550 21519 6552 21528
rect 6604 21519 6606 21528
rect 6644 21548 6696 21554
rect 6552 21490 6604 21496
rect 6644 21490 6696 21496
rect 6656 20602 6684 21490
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6840 20534 6868 21966
rect 7208 21622 7236 22578
rect 7392 22574 7420 26200
rect 7470 24304 7526 24313
rect 7470 24239 7526 24248
rect 7484 24206 7512 24239
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 22642 7512 24006
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26200 10654 27000
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26330 12586 27000
rect 13174 26330 13230 27000
rect 12530 26302 12848 26330
rect 12530 26200 12586 26302
rect 8680 24274 8708 26200
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7196 21616 7248 21622
rect 7196 21558 7248 21564
rect 7208 21146 7236 21558
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 7300 19514 7328 22510
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8312 21298 8340 23666
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8404 21894 8432 23598
rect 9140 23118 9168 24006
rect 9220 23656 9272 23662
rect 9324 23610 9352 26200
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 9272 23604 9352 23610
rect 9220 23598 9352 23604
rect 9232 23582 9352 23598
rect 9220 23248 9272 23254
rect 9220 23190 9272 23196
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 22030 9168 22442
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8312 21270 8432 21298
rect 8404 20942 8432 21270
rect 8392 20936 8444 20942
rect 8390 20904 8392 20913
rect 8444 20904 8446 20913
rect 8496 20874 8524 21898
rect 9232 21146 9260 23190
rect 9508 21690 9536 24074
rect 9784 22098 9812 25434
rect 9968 22710 9996 26200
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9586 21584 9642 21593
rect 9586 21519 9588 21528
rect 9640 21519 9642 21528
rect 9588 21490 9640 21496
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 8390 20839 8446 20848
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5828 19174 5856 19314
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5632 18352 5684 18358
rect 5632 18294 5684 18300
rect 5828 17134 5856 19110
rect 6840 18970 6868 19246
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 1032 16040 1084 16046
rect 1032 15982 1084 15988
rect 1044 15881 1072 15982
rect 1030 15872 1086 15881
rect 1030 15807 1086 15816
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 938 15464 994 15473
rect 938 15399 940 15408
rect 992 15399 994 15408
rect 940 15370 992 15376
rect 938 15056 994 15065
rect 938 14991 940 15000
rect 992 14991 994 15000
rect 940 14962 992 14968
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 938 14648 994 14657
rect 2950 14651 3258 14660
rect 938 14583 994 14592
rect 952 14482 980 14583
rect 940 14476 992 14482
rect 940 14418 992 14424
rect 1030 14240 1086 14249
rect 1030 14175 1086 14184
rect 1044 14006 1072 14175
rect 1032 14000 1084 14006
rect 1032 13942 1084 13948
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 1766 13832 1822 13841
rect 1766 13767 1822 13776
rect 1780 13394 1808 13767
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3528 13433 3556 13874
rect 3514 13424 3570 13433
rect 1768 13388 1820 13394
rect 3514 13359 3570 13368
rect 1768 13330 1820 13336
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 12918 1348 12951
rect 1308 12912 1360 12918
rect 1308 12854 1360 12860
rect 1216 12844 1268 12850
rect 1216 12786 1268 12792
rect 1228 12617 1256 12786
rect 1214 12608 1270 12617
rect 1214 12543 1270 12552
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 1308 12300 1360 12306
rect 1308 12242 1360 12248
rect 1214 12200 1270 12209
rect 1214 12135 1270 12144
rect 1228 11762 1256 12135
rect 1320 11801 1348 12242
rect 4264 11898 4292 16050
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4724 15026 4752 15370
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 5460 12986 5488 16594
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5828 12238 5856 17070
rect 6840 15910 6868 18090
rect 7760 16590 7788 19450
rect 8312 19174 8340 19926
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 17338 7880 18566
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16250 8340 19110
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9048 16454 9076 16594
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 9048 16046 9076 16390
rect 9232 16250 9260 19382
rect 9600 19378 9628 20946
rect 9692 20602 9720 22034
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9862 20496 9918 20505
rect 9772 20460 9824 20466
rect 9862 20431 9864 20440
rect 9772 20402 9824 20408
rect 9916 20431 9918 20440
rect 9864 20402 9916 20408
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9784 18086 9812 20402
rect 9968 19990 9996 21490
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9968 19417 9996 19790
rect 9954 19408 10010 19417
rect 9954 19343 10010 19352
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9876 18426 9904 19246
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 10060 18358 10088 24346
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10336 20602 10364 23802
rect 10612 23662 10640 26200
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 11164 22642 11192 24006
rect 11256 23186 11284 26200
rect 11900 25242 11928 26200
rect 11808 25214 11928 25242
rect 11808 24274 11836 25214
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23798 11836 24006
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11888 23112 11940 23118
rect 11334 23080 11390 23089
rect 11888 23054 11940 23060
rect 11334 23015 11390 23024
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11244 22500 11296 22506
rect 11244 22442 11296 22448
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10782 20360 10838 20369
rect 10782 20295 10784 20304
rect 10836 20295 10838 20304
rect 10784 20266 10836 20272
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 10244 17882 10272 18634
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10612 17882 10640 18158
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9508 16998 9536 17138
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 9048 15366 9076 15982
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 9048 13258 9076 15302
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 9508 12782 9536 16934
rect 10428 16794 10456 17614
rect 10506 17232 10562 17241
rect 10506 17167 10508 17176
rect 10560 17167 10562 17176
rect 10508 17138 10560 17144
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9692 15162 9720 16458
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15162 9812 15914
rect 10336 15910 10364 16662
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9784 13734 9812 14894
rect 10244 14550 10272 15438
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 14074 9996 14350
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10336 13870 10364 15846
rect 10520 15337 10548 16458
rect 10704 15706 10732 18634
rect 10796 17202 10824 19926
rect 10888 19718 10916 20742
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10888 16697 10916 19654
rect 10980 19122 11008 21490
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20602 11100 20878
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11072 19281 11100 20334
rect 11058 19272 11114 19281
rect 11058 19207 11114 19216
rect 10980 19094 11100 19122
rect 11072 18970 11100 19094
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10874 16688 10930 16697
rect 10980 16658 11008 18906
rect 11164 18902 11192 20742
rect 11152 18896 11204 18902
rect 11256 18873 11284 22442
rect 11348 20942 11376 23015
rect 11900 22234 11928 23054
rect 11980 22500 12032 22506
rect 11980 22442 12032 22448
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11992 22098 12020 22442
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 11702 21992 11758 22001
rect 11702 21927 11758 21936
rect 11716 21622 11744 21927
rect 11428 21616 11480 21622
rect 11428 21558 11480 21564
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11440 19786 11468 21558
rect 12360 21554 12388 22374
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11716 20448 11744 21286
rect 11808 20942 11836 21354
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 21146 12296 21286
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 12072 20936 12124 20942
rect 12360 20890 12388 21490
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12452 21146 12480 21422
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12072 20878 12124 20884
rect 11888 20460 11940 20466
rect 11716 20420 11888 20448
rect 11888 20402 11940 20408
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11152 18838 11204 18844
rect 11242 18864 11298 18873
rect 11242 18799 11298 18808
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 10874 16623 10930 16632
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10796 15609 10824 15982
rect 10782 15600 10838 15609
rect 10782 15535 10838 15544
rect 10506 15328 10562 15337
rect 10506 15263 10562 15272
rect 10888 15094 10916 16118
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15706 11008 15982
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 15094 11008 15370
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10612 14822 10640 14962
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10414 14376 10470 14385
rect 10414 14311 10416 14320
rect 10468 14311 10470 14320
rect 10416 14282 10468 14288
rect 10428 14074 10456 14282
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10520 14006 10548 14214
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 9784 12170 9812 13670
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 2136 11824 2188 11830
rect 1306 11792 1362 11801
rect 1216 11756 1268 11762
rect 2136 11766 2188 11772
rect 1306 11727 1362 11736
rect 1216 11698 1268 11704
rect 1228 11354 1256 11698
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1320 11393 1348 11630
rect 1306 11384 1362 11393
rect 1216 11348 1268 11354
rect 1306 11319 1362 11328
rect 1216 11290 1268 11296
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10985 1624 11086
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1216 10736 1268 10742
rect 1216 10678 1268 10684
rect 1228 10169 1256 10678
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10577 1348 10610
rect 1306 10568 1362 10577
rect 1306 10503 1362 10512
rect 1214 10160 1270 10169
rect 2148 10130 2176 11766
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 1214 10095 1270 10104
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 1306 9752 1362 9761
rect 2424 9722 2452 9998
rect 1306 9687 1308 9696
rect 1360 9687 1362 9696
rect 2412 9716 2464 9722
rect 1308 9658 1360 9664
rect 2412 9658 2464 9664
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 9353 1348 9522
rect 1766 9480 1822 9489
rect 1766 9415 1768 9424
rect 1820 9415 1822 9424
rect 1768 9386 1820 9392
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1306 8936 1362 8945
rect 1228 8537 1256 8910
rect 1306 8871 1308 8880
rect 1360 8871 1362 8880
rect 1308 8842 1360 8848
rect 1214 8528 1270 8537
rect 2148 8498 2176 9046
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3160 8838 3188 8978
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 1214 8463 1270 8472
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 1306 8120 1362 8129
rect 2424 8090 2452 8366
rect 1306 8055 1308 8064
rect 1360 8055 1362 8064
rect 2412 8084 2464 8090
rect 1308 8026 1360 8032
rect 2412 8026 2464 8032
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 7721 1348 7822
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 7313 1348 7346
rect 1306 7304 1362 7313
rect 1306 7239 1362 7248
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6730 1256 6831
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1216 6724 1268 6730
rect 1216 6666 1268 6672
rect 1228 6458 1256 6666
rect 1320 6497 1348 6734
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1306 6488 1362 6497
rect 1216 6452 1268 6458
rect 1306 6423 1362 6432
rect 1216 6394 1268 6400
rect 1780 6322 1808 6598
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1320 6089 1348 6258
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 2608 5914 2636 8774
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 1360 5672 1362 5681
rect 1306 5607 1362 5616
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4865 1348 5102
rect 1306 4856 1362 4865
rect 1306 4791 1308 4800
rect 1360 4791 1362 4800
rect 1308 4762 1360 4768
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1320 4457 1348 4558
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1400 4208 1452 4214
rect 1400 4150 1452 4156
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1320 3641 1348 4082
rect 1412 4049 1440 4150
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1306 3632 1362 3641
rect 1306 3567 1362 3576
rect 1122 3496 1178 3505
rect 1122 3431 1178 3440
rect 1308 3460 1360 3466
rect 1136 800 1164 3431
rect 1308 3402 1360 3408
rect 1320 3233 1348 3402
rect 1306 3224 1362 3233
rect 1306 3159 1308 3168
rect 1360 3159 1362 3168
rect 1308 3130 1360 3136
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1320 2825 1348 2994
rect 1780 2922 1808 4218
rect 2700 3602 2728 7822
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 5273 2820 5646
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 4080 4758 4108 6122
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4448 4010 4476 4966
rect 4816 4282 4844 10134
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 10612 6730 10640 14758
rect 11256 14618 11284 18294
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 17270 11468 17682
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11624 16561 11652 19314
rect 11716 18222 11744 19722
rect 11808 18426 11836 20198
rect 11900 19689 11928 20402
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11992 19922 12020 19994
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11886 19680 11942 19689
rect 11886 19615 11942 19624
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18970 11928 19110
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 17542 11744 18022
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11610 16552 11666 16561
rect 11610 16487 11666 16496
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11348 16250 11376 16390
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11440 15910 11468 16118
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11256 14006 11284 14282
rect 11244 14000 11296 14006
rect 11242 13968 11244 13977
rect 11296 13968 11298 13977
rect 11242 13903 11298 13912
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10796 12306 10824 13330
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11150 13152 11206 13161
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10888 12238 10916 13126
rect 10980 12986 11008 13126
rect 11150 13087 11206 13096
rect 11164 12986 11192 13087
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11150 12880 11206 12889
rect 11150 12815 11206 12824
rect 11164 12646 11192 12815
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11898 10916 12174
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11072 11218 11100 12106
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 9518 11100 11154
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 11164 6254 11192 12582
rect 11440 11626 11468 15846
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11624 10713 11652 15030
rect 11716 12866 11744 16050
rect 11808 15162 11836 18226
rect 11992 17610 12020 18566
rect 12084 17728 12112 20878
rect 12268 20862 12388 20890
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12176 18873 12204 19314
rect 12268 19242 12296 20862
rect 12452 20058 12480 21082
rect 12544 20534 12572 21626
rect 12636 21622 12664 24074
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12728 21078 12756 23666
rect 12820 22710 12848 26302
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 23186 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26200 16450 27000
rect 17038 26200 17094 27000
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26330 25466 27000
rect 25240 26302 25466 26330
rect 13832 24274 13860 26200
rect 14476 24290 14504 26200
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 14384 24262 14504 24290
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 14200 23322 14228 23734
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13280 21962 13308 22034
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12716 21072 12768 21078
rect 12820 21049 12848 21286
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 21146 13400 21830
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 12716 21014 12768 21020
rect 12806 21040 12862 21049
rect 12806 20975 12862 20984
rect 13452 21004 13504 21010
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12544 19530 12572 20334
rect 12360 19502 12572 19530
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12162 18864 12218 18873
rect 12162 18799 12218 18808
rect 12360 18630 12388 19502
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12452 18358 12480 19314
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12544 18222 12572 18838
rect 12636 18442 12664 20810
rect 12820 20534 12848 20975
rect 13452 20946 13504 20952
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 13188 20262 13216 20810
rect 13464 20534 13492 20946
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 12820 19768 12848 20198
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12900 19780 12952 19786
rect 12820 19740 12900 19768
rect 12900 19722 12952 19728
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18902 12756 19110
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12820 18698 12848 19382
rect 12912 19378 12940 19722
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12636 18414 12756 18442
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12532 17740 12584 17746
rect 12084 17700 12388 17728
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11900 17105 11928 17206
rect 11886 17096 11942 17105
rect 11886 17031 11942 17040
rect 11992 15434 12020 17546
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11888 15360 11940 15366
rect 11940 15308 12020 15314
rect 11888 15302 12020 15308
rect 11900 15286 12020 15302
rect 11992 15162 12020 15286
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12084 14890 12112 17546
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12176 16998 12204 17206
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 11992 12986 12020 14826
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 12084 13394 12112 13738
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12176 12986 12204 15642
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 11716 12838 12020 12866
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 12442 11836 12718
rect 11992 12442 12020 12838
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11808 11762 11836 12378
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11808 11218 11836 11698
rect 12268 11626 12296 16526
rect 12360 15162 12388 17700
rect 12532 17682 12584 17688
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16658 12480 16934
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12360 14074 12388 15098
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12360 13394 12388 13670
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12360 12306 12388 13194
rect 12452 12782 12480 16390
rect 12544 15570 12572 17682
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12636 15502 12664 17002
rect 12728 16454 12756 18414
rect 13188 18358 13216 18770
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13280 18358 13308 18566
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17338 13400 18838
rect 13464 18766 13492 19450
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13464 18290 13492 18702
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13464 17746 13492 18226
rect 13556 17882 13584 21966
rect 13648 19961 13676 22578
rect 13740 21690 13768 23054
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22438 14136 22918
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 21894 14136 22374
rect 14292 22098 14320 24142
rect 14384 23798 14412 24262
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13924 20806 13952 21830
rect 14108 21690 14136 21830
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13634 19952 13690 19961
rect 13634 19887 13690 19896
rect 13648 18902 13676 19887
rect 13832 19825 13860 20742
rect 13818 19816 13874 19825
rect 13818 19751 13874 19760
rect 13726 19408 13782 19417
rect 13726 19343 13782 19352
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13544 17536 13596 17542
rect 13648 17524 13676 18022
rect 13596 17496 13676 17524
rect 13544 17478 13596 17484
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12820 16640 12848 17070
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12820 16612 12940 16640
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 14822 12572 15370
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12728 14362 12756 15846
rect 12820 14618 12848 16458
rect 12912 15910 12940 16612
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 16114 13308 16390
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13188 16017 13216 16050
rect 13360 16040 13412 16046
rect 13174 16008 13230 16017
rect 13360 15982 13412 15988
rect 13174 15943 13230 15952
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12900 15632 12952 15638
rect 12900 15574 12952 15580
rect 12912 15162 12940 15574
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13372 14482 13400 15982
rect 13464 15502 13492 16934
rect 13556 16130 13584 17478
rect 13556 16102 13676 16130
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13464 14550 13492 15030
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 12544 14334 12756 14362
rect 12808 14340 12860 14346
rect 12544 12986 12572 14334
rect 12808 14282 12860 14288
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13172 12664 14214
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13240 12756 13670
rect 12820 13394 12848 14282
rect 13280 14006 13308 14418
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13280 13716 13308 13942
rect 13280 13688 13400 13716
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12728 13212 12940 13240
rect 12636 13144 12848 13172
rect 12532 12980 12584 12986
rect 12584 12940 12664 12968
rect 12532 12922 12584 12928
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12636 12646 12664 12940
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12544 12434 12572 12582
rect 12544 12406 12664 12434
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12360 11898 12388 12242
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11610 10704 11666 10713
rect 11610 10639 11666 10648
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10470 12296 10610
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5354 4040 5410 4049
rect 4436 4004 4488 4010
rect 5354 3975 5410 3984
rect 4436 3946 4488 3952
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 2320 2848 2372 2854
rect 1306 2816 1362 2825
rect 2320 2790 2372 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1306 2751 1362 2760
rect 1308 2440 1360 2446
rect 1306 2408 1308 2417
rect 1360 2408 1362 2417
rect 1216 2372 1268 2378
rect 2332 2378 2360 2790
rect 2792 2446 2820 2790
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 1306 2343 1362 2352
rect 2320 2372 2372 2378
rect 1216 2314 1268 2320
rect 2320 2314 2372 2320
rect 1228 2009 1256 2314
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1601 1348 2246
rect 3344 1850 3372 3538
rect 3252 1822 3372 1850
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 3252 800 3280 1822
rect 5368 800 5396 3975
rect 6840 3942 6868 4762
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7484 800 7512 3606
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 10336 3194 10364 3470
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9600 800 9628 2994
rect 9784 2582 9812 2994
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 10704 2446 10732 3334
rect 12268 2514 12296 10406
rect 12360 9586 12388 11494
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10810 12572 10950
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 10198 12572 10406
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12452 7886 12480 9862
rect 12636 9654 12664 12406
rect 12728 11898 12756 12650
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12728 11286 12756 11562
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12728 8634 12756 11086
rect 12820 10810 12848 13144
rect 12912 12714 12940 13212
rect 13268 12980 13320 12986
rect 13372 12968 13400 13688
rect 13320 12940 13400 12968
rect 13268 12922 13320 12928
rect 13556 12866 13584 15302
rect 13648 14482 13676 16102
rect 13740 16028 13768 19343
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18329 13952 18566
rect 13910 18320 13966 18329
rect 13820 18284 13872 18290
rect 13910 18255 13966 18264
rect 13820 18226 13872 18232
rect 13832 16590 13860 18226
rect 13924 17270 13952 18255
rect 14016 17338 14044 21490
rect 14108 20874 14136 21626
rect 14188 21616 14240 21622
rect 14188 21558 14240 21564
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 14200 18290 14228 21558
rect 14292 21146 14320 21558
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14384 21146 14412 21490
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14292 20398 14320 21082
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14476 20058 14504 24142
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22642 14688 22918
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14568 21486 14596 22374
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19553 14320 19790
rect 14278 19544 14334 19553
rect 14278 19479 14334 19488
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16658 14136 16934
rect 14476 16833 14504 19110
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14568 18222 14596 18634
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14568 17882 14596 18158
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14660 17134 14688 21898
rect 14936 20602 14964 24074
rect 15120 22710 15148 26200
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 14922 20360 14978 20369
rect 14922 20295 14978 20304
rect 14936 19990 14964 20295
rect 14924 19984 14976 19990
rect 14924 19926 14976 19932
rect 15028 19514 15056 22646
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15488 22234 15516 22510
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15304 21622 15332 21898
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 15474 21584 15530 21593
rect 15474 21519 15530 21528
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 15120 18306 15148 20402
rect 15290 20360 15346 20369
rect 15290 20295 15346 20304
rect 15198 19408 15254 19417
rect 15198 19343 15200 19352
rect 15252 19343 15254 19352
rect 15200 19314 15252 19320
rect 15304 19310 15332 20295
rect 15488 20262 15516 21519
rect 15580 20602 15608 24278
rect 15660 23248 15712 23254
rect 15660 23190 15712 23196
rect 15672 20602 15700 23190
rect 15764 23186 15792 26200
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19854 15516 20198
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15292 19304 15344 19310
rect 15568 19304 15620 19310
rect 15292 19246 15344 19252
rect 15566 19272 15568 19281
rect 15620 19272 15622 19281
rect 15304 19174 15332 19246
rect 15566 19207 15622 19216
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15028 18278 15148 18306
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14462 16824 14518 16833
rect 14462 16759 14518 16768
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 13820 16040 13872 16046
rect 13740 16000 13820 16028
rect 13740 15502 13768 16000
rect 13820 15982 13872 15988
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13924 15162 13952 15914
rect 14016 15910 14044 16118
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14016 14521 14044 14554
rect 14002 14512 14058 14521
rect 13636 14476 13688 14482
rect 14002 14447 14058 14456
rect 13636 14418 13688 14424
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13648 12986 13676 13806
rect 13728 13524 13780 13530
rect 13832 13512 13860 14350
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13780 13484 13860 13512
rect 13728 13466 13780 13472
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13556 12838 13676 12866
rect 13544 12776 13596 12782
rect 13450 12744 13506 12753
rect 12900 12708 12952 12714
rect 13544 12718 13596 12724
rect 13450 12679 13506 12688
rect 12900 12650 12952 12656
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13464 12434 13492 12679
rect 13280 12406 13492 12434
rect 13280 11694 13308 12406
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13358 11928 13414 11937
rect 13358 11863 13360 11872
rect 13412 11863 13414 11872
rect 13360 11834 13412 11840
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12912 10690 12940 11018
rect 12820 10662 12940 10690
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12820 5234 12848 10662
rect 13268 10600 13320 10606
rect 13266 10568 13268 10577
rect 13320 10568 13322 10577
rect 13266 10503 13322 10512
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13096 9926 13124 9998
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13372 9042 13400 11834
rect 13464 10538 13492 12106
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13556 8974 13584 12718
rect 13648 11898 13676 12838
rect 13740 12753 13768 13466
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13832 13190 13860 13330
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13726 12744 13782 12753
rect 13726 12679 13782 12688
rect 13832 12434 13860 13126
rect 13740 12406 13860 12434
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13648 9466 13676 11630
rect 13740 9654 13768 12406
rect 13818 12200 13874 12209
rect 13818 12135 13874 12144
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13648 9438 13768 9466
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13740 8906 13768 9438
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13740 7818 13768 8842
rect 13832 8838 13860 12135
rect 13924 11354 13952 14214
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14016 13394 14044 13466
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14108 13274 14136 16594
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14200 14618 14228 16390
rect 14292 16153 14320 16662
rect 14752 16590 14780 17206
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14278 16144 14334 16153
rect 14334 16102 14412 16130
rect 14278 16079 14334 16088
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14292 15094 14320 15914
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14292 14822 14320 15030
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14292 14074 14320 14758
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14384 13920 14412 16102
rect 14844 16046 14872 16730
rect 15028 16114 15056 18278
rect 15108 18080 15160 18086
rect 15160 18040 15240 18068
rect 15108 18022 15160 18028
rect 15212 17202 15240 18040
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15120 16810 15148 17138
rect 15120 16782 15240 16810
rect 15106 16688 15162 16697
rect 15106 16623 15162 16632
rect 15120 16250 15148 16623
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14832 16040 14884 16046
rect 14554 16008 14610 16017
rect 14832 15982 14884 15988
rect 14554 15943 14610 15952
rect 14568 15162 14596 15943
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14464 14952 14516 14958
rect 14516 14900 14596 14906
rect 14464 14894 14596 14900
rect 14476 14878 14596 14894
rect 14568 14090 14596 14878
rect 14660 14618 14688 15302
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14752 14822 14780 15030
rect 14844 14958 14872 15982
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14844 14278 14872 14418
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14568 14062 14872 14090
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14384 13892 14596 13920
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14370 13696 14426 13705
rect 14370 13631 14426 13640
rect 14016 13246 14136 13274
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14016 11830 14044 13246
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14016 10538 14044 11630
rect 14108 10742 14136 13126
rect 14292 12434 14320 13262
rect 14200 12406 14320 12434
rect 14200 12102 14228 12406
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 14016 10146 14044 10474
rect 13924 10118 14044 10146
rect 13924 9926 13952 10118
rect 14200 9994 14228 12038
rect 14384 11744 14412 13631
rect 14476 13326 14504 13738
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14476 13161 14504 13262
rect 14462 13152 14518 13161
rect 14462 13087 14518 13096
rect 14568 13002 14596 13892
rect 14752 13462 14780 13942
rect 14740 13456 14792 13462
rect 14738 13424 14740 13433
rect 14792 13424 14794 13433
rect 14738 13359 14794 13368
rect 14292 11716 14412 11744
rect 14476 12974 14596 13002
rect 14292 10062 14320 11716
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14384 10810 14412 11562
rect 14476 11218 14504 12974
rect 14648 12912 14700 12918
rect 14752 12900 14780 13359
rect 14700 12872 14780 12900
rect 14648 12854 14700 12860
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 11354 14596 12718
rect 14752 12238 14780 12872
rect 14844 12306 14872 14062
rect 14936 13258 14964 15506
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15028 13530 15056 14350
rect 15120 13870 15148 15574
rect 15212 14226 15240 16782
rect 15304 15978 15332 17546
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15396 15638 15424 17682
rect 15580 17338 15608 18566
rect 15672 17610 15700 18702
rect 15764 18154 15792 21082
rect 16040 20602 16068 24754
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 16224 23866 16252 24618
rect 16212 23860 16264 23866
rect 16212 23802 16264 23808
rect 16408 23662 16436 26200
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16592 22234 16620 22578
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16592 21350 16620 21898
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15842 19680 15898 19689
rect 15842 19615 15898 19624
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15856 17524 15884 19615
rect 15948 19514 15976 20334
rect 16132 19854 16160 20810
rect 16316 19922 16344 21082
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15936 19236 15988 19242
rect 15936 19178 15988 19184
rect 15948 18970 15976 19178
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 16040 17746 16068 19382
rect 16132 19310 16160 19790
rect 16210 19408 16266 19417
rect 16210 19343 16212 19352
rect 16264 19343 16266 19352
rect 16212 19314 16264 19320
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15936 17536 15988 17542
rect 15856 17496 15936 17524
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15396 14482 15424 14826
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15212 14198 15332 14226
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11762 14780 12174
rect 14844 11830 14872 12242
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14740 11756 14792 11762
rect 14660 11716 14740 11744
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14568 10606 14596 11290
rect 14660 11014 14688 11716
rect 14740 11698 14792 11704
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11218 14872 11494
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14660 10062 14688 10950
rect 14752 10198 14780 10950
rect 14936 10606 14964 13194
rect 15028 12986 15056 13466
rect 15120 13394 15148 13806
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15212 11898 15240 14010
rect 15304 12714 15332 14198
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15396 12594 15424 14418
rect 15488 13394 15516 16390
rect 15580 16046 15608 16662
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15580 15570 15608 15982
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15580 13326 15608 15302
rect 15672 14958 15700 16390
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15764 14770 15792 17206
rect 15856 16590 15884 17496
rect 15936 17478 15988 17484
rect 16040 17270 16068 17682
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15842 16144 15898 16153
rect 15842 16079 15898 16088
rect 15856 16046 15884 16079
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15672 14742 15792 14770
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15488 12782 15516 12854
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15304 12566 15424 12594
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15304 11218 15332 12566
rect 15488 12306 15516 12718
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15580 12170 15608 12582
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15568 11688 15620 11694
rect 15672 11676 15700 14742
rect 15856 13938 15884 15574
rect 16040 15094 16068 17206
rect 16132 17134 16160 18906
rect 16592 18902 16620 21286
rect 16684 21078 16712 21626
rect 16868 21418 16896 22578
rect 17052 22166 17080 26200
rect 17696 24274 17724 26200
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17040 22160 17092 22166
rect 17040 22102 17092 22108
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16684 18970 16712 21014
rect 16868 20942 16896 21354
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16776 18970 16804 20742
rect 16868 20466 16896 20878
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16316 18154 16344 18838
rect 16684 18766 16712 18906
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16684 18222 16712 18702
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16316 17542 16344 17682
rect 16500 17678 16528 18158
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16500 17066 16528 17478
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16394 16552 16450 16561
rect 16394 16487 16450 16496
rect 16408 16250 16436 16487
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16210 15600 16266 15609
rect 16120 15564 16172 15570
rect 16210 15535 16266 15544
rect 16120 15506 16172 15512
rect 16028 15088 16080 15094
rect 16028 15030 16080 15036
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14074 15976 14758
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 16132 13462 16160 15506
rect 16120 13456 16172 13462
rect 16120 13398 16172 13404
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15764 12306 15792 13330
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15856 12889 15884 12922
rect 15842 12880 15898 12889
rect 15842 12815 15898 12824
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15856 12050 15884 12650
rect 15620 11648 15700 11676
rect 15764 12022 15884 12050
rect 15568 11630 15620 11636
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 10266 15056 10542
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14280 10056 14332 10062
rect 14648 10056 14700 10062
rect 14280 9998 14332 10004
rect 14646 10024 14648 10033
rect 14700 10024 14702 10033
rect 14188 9988 14240 9994
rect 14646 9959 14702 9968
rect 14188 9930 14240 9936
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13924 8566 13952 9862
rect 14752 9722 14780 10134
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15120 9738 15148 9959
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 15120 9710 15332 9738
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 14476 6254 14504 8774
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13740 3602 13768 4218
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 14108 2446 14136 3402
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 11716 800 11744 2314
rect 13832 800 13860 2314
rect 14752 2310 14780 9658
rect 15120 9654 15148 9710
rect 15108 9648 15160 9654
rect 15108 9590 15160 9596
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14936 7886 14964 9318
rect 15120 9042 15148 9454
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15120 8430 15148 8978
rect 15212 8634 15240 9590
rect 15304 8838 15332 9710
rect 15396 9110 15424 11494
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15488 9042 15516 11562
rect 15580 11082 15608 11630
rect 15764 11370 15792 12022
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15672 11342 15792 11370
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15672 10470 15700 11342
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15580 8974 15608 10406
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15212 8498 15240 8570
rect 15304 8566 15332 8774
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15212 3194 15240 8434
rect 15672 6866 15700 9318
rect 15764 9178 15792 11154
rect 15856 9586 15884 11834
rect 15948 11218 15976 13126
rect 16132 12782 16160 13398
rect 16224 12918 16252 15535
rect 16316 15366 16344 16118
rect 16592 15706 16620 18022
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16408 15366 16436 15506
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16316 14890 16344 15302
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16316 13734 16344 14826
rect 16578 14512 16634 14521
rect 16578 14447 16634 14456
rect 16592 14278 16620 14447
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16486 13832 16542 13841
rect 16486 13767 16542 13776
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16316 12918 16344 13330
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16210 12744 16266 12753
rect 16210 12679 16266 12688
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 11354 16160 11630
rect 16224 11558 16252 12679
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16132 10266 16160 11154
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16224 10062 16252 10610
rect 16316 10130 16344 12582
rect 16500 11914 16528 13767
rect 16408 11898 16528 11914
rect 16396 11892 16528 11898
rect 16448 11886 16528 11892
rect 16396 11834 16448 11840
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16040 9654 16068 9998
rect 16224 9654 16252 9998
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 5030 15700 6802
rect 15948 6798 15976 8774
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16316 5642 16344 9318
rect 16408 7818 16436 11290
rect 16592 11082 16620 14010
rect 16684 12442 16712 17818
rect 16776 17626 16804 18566
rect 16868 17746 16896 20266
rect 16960 19446 16988 21966
rect 17144 21962 17172 22918
rect 17512 22692 17540 23054
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17592 22704 17644 22710
rect 17512 22664 17592 22692
rect 17512 22574 17540 22664
rect 17592 22646 17644 22652
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17144 20602 17172 21898
rect 17236 21622 17264 22170
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17420 20505 17448 21626
rect 17512 21078 17540 22510
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17512 20942 17540 21014
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17512 20602 17540 20878
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17406 20496 17462 20505
rect 17406 20431 17462 20440
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 17052 19378 17080 20198
rect 17144 19718 17172 20198
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16776 17598 16896 17626
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16776 15434 16804 16934
rect 16868 16658 16896 17598
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16960 16522 16988 17138
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16856 16176 16908 16182
rect 16856 16118 16908 16124
rect 16868 15473 16896 16118
rect 16948 15904 17000 15910
rect 17052 15892 17080 19314
rect 17236 17882 17264 19654
rect 17328 19514 17356 19654
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17512 19446 17540 20538
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 17604 19378 17632 19858
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17406 18728 17462 18737
rect 17406 18663 17408 18672
rect 17460 18663 17462 18672
rect 17408 18634 17460 18640
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 16998 17448 17478
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16794 17448 16934
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17512 16590 17540 18158
rect 17788 18057 17816 22918
rect 17880 21690 17908 24550
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23662 18368 26200
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18892 24206 18920 24686
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18696 24132 18748 24138
rect 18696 24074 18748 24080
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17866 20496 17922 20505
rect 17866 20431 17922 20440
rect 17774 18048 17830 18057
rect 17774 17983 17830 17992
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17144 16182 17172 16390
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17000 15864 17080 15892
rect 16948 15846 17000 15852
rect 16854 15464 16910 15473
rect 16764 15428 16816 15434
rect 16854 15399 16910 15408
rect 16764 15370 16816 15376
rect 16868 14278 16896 15399
rect 16960 14958 16988 15846
rect 17144 15434 17172 15982
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16776 12186 16804 13874
rect 16684 12158 16804 12186
rect 16684 12102 16712 12158
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16776 10742 16804 12038
rect 16960 11626 16988 14894
rect 17144 13705 17172 15370
rect 17328 15337 17356 15846
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 14278 17264 14826
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17130 13696 17186 13705
rect 17130 13631 17186 13640
rect 17130 13424 17186 13433
rect 17130 13359 17186 13368
rect 17144 13258 17172 13359
rect 17132 13252 17184 13258
rect 17052 13212 17132 13240
rect 17052 12850 17080 13212
rect 17132 13194 17184 13200
rect 17236 13138 17264 14214
rect 17328 13841 17356 15263
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17314 13832 17370 13841
rect 17314 13767 17370 13776
rect 17314 13696 17370 13705
rect 17314 13631 17370 13640
rect 17144 13110 17264 13138
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 11898 17080 12786
rect 17144 12714 17172 13110
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 17144 11354 17172 12650
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 11937 17264 12174
rect 17222 11928 17278 11937
rect 17222 11863 17278 11872
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 16764 10736 16816 10742
rect 16486 10704 16542 10713
rect 16764 10678 16816 10684
rect 16486 10639 16542 10648
rect 16500 10266 16528 10639
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9722 16620 9862
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16684 9654 16712 10542
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16776 9110 16804 9930
rect 16868 9654 16896 11290
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17052 10742 17080 11086
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 17328 10674 17356 13631
rect 17420 12306 17448 14350
rect 17512 14074 17540 14826
rect 17604 14074 17632 15914
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17696 13938 17724 14350
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17788 12714 17816 16050
rect 17880 15706 17908 20431
rect 18340 20058 18368 21490
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18340 18970 18368 19722
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18524 18850 18552 20742
rect 18616 19854 18644 24006
rect 18708 23050 18736 24074
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 18708 22778 18736 22986
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18800 22234 18828 23462
rect 18892 22982 18920 23734
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22574 18920 22918
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18694 21992 18750 22001
rect 18694 21927 18750 21936
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18708 19360 18736 21927
rect 18800 21622 18828 22170
rect 18984 21962 19012 26200
rect 19524 24268 19576 24274
rect 19628 24256 19656 26200
rect 19576 24228 19656 24256
rect 19524 24210 19576 24216
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 19076 22574 19104 23122
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19352 22778 19380 23054
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18892 21842 18920 21898
rect 18892 21814 19012 21842
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18984 21486 19012 21814
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18892 20602 18920 21422
rect 19064 21072 19116 21078
rect 19064 21014 19116 21020
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18892 19990 18920 20538
rect 19076 20534 19104 21014
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 19076 19718 19104 20470
rect 19260 19990 19288 22510
rect 19352 21350 19380 22714
rect 19444 22030 19472 24006
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19628 23254 19656 23802
rect 20272 23322 20300 26200
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19812 22681 19840 22986
rect 20364 22982 20392 23734
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 19798 22672 19854 22681
rect 19798 22607 19854 22616
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20942 19380 21286
rect 19720 21146 19748 22510
rect 19892 22160 19944 22166
rect 19892 22102 19944 22108
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19812 21146 19840 21626
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19432 20868 19484 20874
rect 19432 20810 19484 20816
rect 19444 20602 19472 20810
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 18708 19332 18828 19360
rect 18604 19304 18656 19310
rect 18656 19264 18736 19292
rect 18604 19246 18656 19252
rect 18432 18822 18552 18850
rect 18602 18864 18658 18873
rect 18432 18630 18460 18822
rect 18602 18799 18658 18808
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18524 18358 18552 18702
rect 18616 18630 18644 18799
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 17524 18276 18226
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18340 17746 18368 18090
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18604 17536 18656 17542
rect 18248 17496 18552 17524
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16658 18000 17206
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17880 15434 17908 15642
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 14074 18368 16186
rect 18420 15632 18472 15638
rect 18418 15600 18420 15609
rect 18472 15600 18474 15609
rect 18418 15535 18474 15544
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18432 14618 18460 15438
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18432 13938 18460 14214
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17972 13530 18000 13738
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17972 11082 18000 11494
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17604 10606 17632 10746
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16500 8498 16528 8978
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16776 7954 16804 8502
rect 16960 7954 16988 9862
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 17052 7886 17080 10406
rect 17696 10198 17724 10542
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17328 9450 17356 9862
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17144 8566 17172 9114
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17420 8634 17448 8842
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17788 8430 17816 11018
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10266 18368 11086
rect 18432 10674 18460 13466
rect 18524 13462 18552 17496
rect 18604 17478 18656 17484
rect 18616 16522 18644 17478
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18616 13870 18644 16458
rect 18708 15366 18736 19264
rect 18800 15706 18828 19332
rect 19444 18834 19472 20538
rect 19628 20262 19656 20742
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19628 19174 19656 20198
rect 19708 19440 19760 19446
rect 19708 19382 19760 19388
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19338 18728 19394 18737
rect 19338 18663 19340 18672
rect 19392 18663 19394 18672
rect 19340 18634 19392 18640
rect 19628 18630 19656 19110
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18892 17202 18920 17614
rect 19168 17338 19196 18294
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19338 18048 19394 18057
rect 19338 17983 19394 17992
rect 19352 17882 19380 17983
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18892 15910 18920 17138
rect 18970 16824 19026 16833
rect 18970 16759 19026 16768
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18800 15042 18828 15642
rect 18708 15026 18828 15042
rect 18696 15020 18828 15026
rect 18748 15014 18828 15020
rect 18696 14962 18748 14968
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18616 11694 18644 12106
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18510 11112 18566 11121
rect 18510 11047 18512 11056
rect 18564 11047 18566 11056
rect 18604 11076 18656 11082
rect 18512 11018 18564 11024
rect 18604 11018 18656 11024
rect 18616 10962 18644 11018
rect 18524 10934 18644 10962
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18432 10130 18460 10610
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 17880 9178 17908 10066
rect 18524 10010 18552 10934
rect 18708 10792 18736 13874
rect 18800 13297 18828 14894
rect 18786 13288 18842 13297
rect 18786 13223 18842 13232
rect 18616 10764 18736 10792
rect 18616 10130 18644 10764
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18432 9982 18552 10010
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18340 9194 18368 9590
rect 18432 9382 18460 9982
rect 18616 9602 18644 10066
rect 18524 9574 18644 9602
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 17868 9172 17920 9178
rect 18340 9166 18460 9194
rect 17868 9114 17920 9120
rect 18432 8906 18460 9166
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18432 8566 18460 8842
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18432 7546 18460 8502
rect 18524 8090 18552 9574
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 8634 18644 9454
rect 18708 8974 18736 10610
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18616 7954 18644 8570
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16592 3534 16620 3946
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 17880 3126 17908 7482
rect 18800 7274 18828 13223
rect 18892 12850 18920 15846
rect 18984 15706 19012 16759
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 18984 14278 19012 15642
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 19076 14074 19104 16390
rect 19168 16114 19196 16594
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19352 14414 19380 16186
rect 19444 15162 19472 18090
rect 19536 17785 19564 18566
rect 19628 18222 19656 18566
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19628 17882 19656 18158
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19522 17776 19578 17785
rect 19522 17711 19578 17720
rect 19536 15706 19564 17711
rect 19720 17338 19748 19382
rect 19812 19310 19840 20878
rect 19904 20602 19932 22102
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 20180 19666 20208 20334
rect 20364 20058 20392 22918
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20640 20262 20668 21898
rect 20732 21622 20760 24346
rect 20916 24274 20944 26200
rect 21560 24954 21588 26200
rect 21548 24948 21600 24954
rect 21548 24890 21600 24896
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 21744 24614 21772 24754
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21732 24608 21784 24614
rect 21732 24550 21784 24556
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20996 24268 21048 24274
rect 20996 24210 21048 24216
rect 20812 22500 20864 22506
rect 20812 22442 20864 22448
rect 20824 22234 20852 22442
rect 21008 22438 21036 24210
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21468 23526 21496 24142
rect 21652 23866 21680 24550
rect 22204 24274 22232 26200
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 21560 23730 21588 23802
rect 21548 23724 21600 23730
rect 21548 23666 21600 23672
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21100 23050 21128 23462
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21088 23044 21140 23050
rect 21088 22986 21140 22992
rect 21100 22710 21128 22986
rect 21192 22778 21220 23122
rect 22112 23118 22140 23598
rect 22480 23322 22508 24210
rect 22572 23662 22600 24346
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 21086 22128 21142 22137
rect 21086 22063 21142 22072
rect 21100 21894 21128 22063
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20916 21350 20944 21490
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 20534 20944 21286
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20916 19854 20944 20470
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20260 19712 20312 19718
rect 20180 19660 20260 19666
rect 20180 19654 20312 19660
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19904 18970 19932 19450
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19996 18358 20024 19654
rect 20180 19638 20300 19654
rect 20180 18834 20208 19638
rect 20364 19446 20392 19790
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 20364 18222 20392 18566
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19996 17134 20024 17750
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20272 17542 20300 17682
rect 20352 17604 20404 17610
rect 20456 17592 20484 19110
rect 20404 17564 20484 17592
rect 20352 17546 20404 17552
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19904 15706 19932 17070
rect 20640 16046 20668 19178
rect 20732 18873 20760 19722
rect 20916 19310 20944 19790
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20812 18896 20864 18902
rect 20718 18864 20774 18873
rect 20812 18838 20864 18844
rect 20718 18799 20774 18808
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19536 15026 19564 15642
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19614 14648 19670 14657
rect 19614 14583 19670 14592
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19444 13938 19472 14282
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 14006 19564 14214
rect 19524 14000 19576 14006
rect 19628 13977 19656 14583
rect 19890 14512 19946 14521
rect 19890 14447 19946 14456
rect 19904 14414 19932 14447
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 14074 19932 14350
rect 19996 14346 20024 15302
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19524 13942 19576 13948
rect 19614 13968 19670 13977
rect 19432 13932 19484 13938
rect 19614 13903 19670 13912
rect 19432 13874 19484 13880
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18984 12918 19012 13806
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18892 12170 18920 12786
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 9518 18920 11630
rect 19168 11286 19196 13466
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19260 11898 19288 12106
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19260 11354 19288 11834
rect 19352 11762 19380 12582
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19444 11354 19472 13874
rect 19892 13184 19944 13190
rect 19996 13172 20024 14282
rect 20088 13530 20116 14418
rect 20272 13530 20300 15302
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 19944 13144 20024 13172
rect 20260 13184 20312 13190
rect 19892 13126 19944 13132
rect 20260 13126 20312 13132
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19536 12238 19564 12718
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19444 10810 19472 10950
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 18970 10704 19026 10713
rect 18970 10639 18972 10648
rect 19024 10639 19026 10648
rect 18972 10610 19024 10616
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18892 9042 18920 9454
rect 19444 9042 19472 10066
rect 19536 9654 19564 11086
rect 19628 10130 19656 12786
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 19720 10810 19748 12718
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19536 9178 19564 9590
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19444 8090 19472 8978
rect 19904 8634 19932 12242
rect 19982 12064 20038 12073
rect 19982 11999 20038 12008
rect 19996 11218 20024 11999
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 20088 11354 20116 11698
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 20180 10656 20208 12718
rect 20272 11626 20300 13126
rect 20364 11830 20392 15302
rect 20732 15042 20760 16730
rect 20824 15706 20852 18838
rect 20916 17592 20944 19246
rect 21008 18970 21036 19858
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21192 18834 21220 22714
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 21652 22234 21680 22578
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21376 21457 21404 21490
rect 21362 21448 21418 21457
rect 21362 21383 21418 21392
rect 21456 21412 21508 21418
rect 21456 21354 21508 21360
rect 21270 21040 21326 21049
rect 21270 20975 21326 20984
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 20996 17604 21048 17610
rect 20916 17564 20996 17592
rect 20916 17338 20944 17564
rect 20996 17546 21048 17552
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20916 16998 20944 17274
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16590 20944 16934
rect 21008 16794 21036 17206
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20916 16454 20944 16526
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20916 16182 20944 16390
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20916 15366 20944 15914
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20548 15014 20760 15042
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20548 14958 20576 15014
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20536 14272 20588 14278
rect 20640 14260 20668 14894
rect 20588 14232 20668 14260
rect 20720 14272 20772 14278
rect 20536 14214 20588 14220
rect 20720 14214 20772 14220
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20456 11558 20484 12718
rect 20548 11937 20576 14214
rect 20628 14000 20680 14006
rect 20732 13988 20760 14214
rect 20680 13960 20760 13988
rect 20628 13942 20680 13948
rect 20640 12764 20668 13942
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20732 13394 20760 13806
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20732 12889 20760 12922
rect 20718 12880 20774 12889
rect 20718 12815 20774 12824
rect 20640 12736 20760 12764
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20534 11928 20590 11937
rect 20534 11863 20590 11872
rect 20534 11792 20590 11801
rect 20534 11727 20536 11736
rect 20588 11727 20590 11736
rect 20536 11698 20588 11704
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20456 11354 20484 11494
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20260 10668 20312 10674
rect 20180 10628 20260 10656
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19996 9722 20024 10542
rect 20180 10266 20208 10628
rect 20260 10610 20312 10616
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 20352 9648 20404 9654
rect 20456 9602 20484 10066
rect 20404 9596 20484 9602
rect 20352 9590 20484 9596
rect 20364 9574 20484 9590
rect 20456 8906 20484 9574
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 4010 18368 6190
rect 18892 5234 18920 7958
rect 19904 7954 19932 8570
rect 20456 8566 20484 8842
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 20456 7818 20484 8502
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 19628 6798 19656 7754
rect 20456 7546 20484 7754
rect 20640 7546 20668 12038
rect 20732 11132 20760 12736
rect 20824 11626 20852 15030
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20916 13530 20944 14962
rect 21100 14890 21128 17818
rect 21192 17746 21220 17818
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21284 15552 21312 20975
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 21376 20602 21404 20810
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 18086 21404 20198
rect 21468 19922 21496 21354
rect 21652 21350 21680 22170
rect 21928 22098 21956 22986
rect 22008 22636 22060 22642
rect 22112 22624 22140 23054
rect 22204 22778 22232 23122
rect 22664 23066 22692 24074
rect 22744 23588 22796 23594
rect 22744 23530 22796 23536
rect 22756 23254 22784 23530
rect 22744 23248 22796 23254
rect 22744 23190 22796 23196
rect 22664 23038 22784 23066
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22060 22596 22232 22624
rect 22008 22578 22060 22584
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 22204 21486 22232 22596
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21546 20632 21602 20641
rect 21546 20567 21602 20576
rect 21560 20534 21588 20567
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21560 20398 21588 20470
rect 22204 20466 22232 21422
rect 22388 20890 22416 21966
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22480 21690 22508 21830
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22572 21010 22600 21830
rect 22664 21010 22692 22034
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22388 20862 22600 20890
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21560 19242 21588 20198
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21468 18358 21496 18566
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21376 17116 21404 18022
rect 21468 17270 21496 18022
rect 21652 17746 21680 19858
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22112 18834 22140 19722
rect 22204 19310 22232 20402
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22192 19304 22244 19310
rect 22192 19246 22244 19252
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21744 17610 21772 18294
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21456 17264 21508 17270
rect 21456 17206 21508 17212
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 21376 17088 21496 17116
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21376 15706 21404 15914
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21468 15570 21496 17088
rect 21560 16998 21588 17206
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21744 16794 21772 17546
rect 21824 17128 21876 17134
rect 21928 17116 21956 18566
rect 22020 17660 22048 18702
rect 22100 17808 22152 17814
rect 22100 17750 22152 17756
rect 22112 17660 22140 17750
rect 22204 17746 22232 19246
rect 22296 17882 22324 20266
rect 22480 20058 22508 20334
rect 22376 20052 22428 20058
rect 22376 19994 22428 20000
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22388 19786 22416 19994
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22572 19666 22600 20862
rect 22756 20330 22784 23038
rect 22848 22982 22876 26200
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23492 23526 23520 26200
rect 24032 24676 24084 24682
rect 24032 24618 24084 24624
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23294 23080 23350 23089
rect 23294 23015 23350 23024
rect 23308 22982 23336 23015
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22848 21894 22876 21966
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 23032 21622 23060 22170
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23216 21332 23244 21558
rect 23216 21304 23336 21332
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 21010 23336 21304
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22940 20602 22968 20878
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22940 20244 22968 20538
rect 23400 20466 23428 23258
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23584 22234 23612 22578
rect 23768 22273 23796 23054
rect 24044 22710 24072 24618
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23754 22264 23810 22273
rect 23572 22228 23624 22234
rect 23754 22199 23810 22208
rect 23572 22170 23624 22176
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23768 20913 23796 21830
rect 23952 21706 23980 21966
rect 24044 21894 24072 22374
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 23952 21678 24072 21706
rect 24044 21622 24072 21678
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 24136 21146 24164 26200
rect 24780 24614 24808 26200
rect 24492 24608 24544 24614
rect 24492 24550 24544 24556
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24504 24138 24532 24550
rect 25240 24206 25268 26302
rect 25410 26200 25466 26302
rect 26054 26330 26110 27000
rect 26698 26330 26754 27000
rect 26054 26302 26188 26330
rect 26054 26200 26110 26302
rect 25964 24948 26016 24954
rect 25964 24890 26016 24896
rect 26056 24948 26108 24954
rect 26056 24890 26108 24896
rect 25872 24880 25924 24886
rect 25872 24822 25924 24828
rect 25780 24336 25832 24342
rect 25778 24304 25780 24313
rect 25832 24304 25834 24313
rect 25778 24239 25834 24248
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 24492 24132 24544 24138
rect 24492 24074 24544 24080
rect 24400 24064 24452 24070
rect 24452 24012 24716 24018
rect 24400 24006 24716 24012
rect 24412 23990 24716 24006
rect 24308 23792 24360 23798
rect 24308 23734 24360 23740
rect 24216 23656 24268 23662
rect 24216 23598 24268 23604
rect 24228 23322 24256 23598
rect 24216 23316 24268 23322
rect 24216 23258 24268 23264
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 24228 22137 24256 22442
rect 24320 22166 24348 23734
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24412 22642 24440 23462
rect 24584 22704 24636 22710
rect 24584 22646 24636 22652
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24596 22438 24624 22646
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24308 22160 24360 22166
rect 24214 22128 24270 22137
rect 24308 22102 24360 22108
rect 24214 22063 24270 22072
rect 24228 21486 24256 22063
rect 24688 21978 24716 23990
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 23322 24900 23462
rect 25056 23322 25084 23666
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 24872 23186 24900 23258
rect 25240 23254 25268 24142
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 25228 23248 25280 23254
rect 25228 23190 25280 23196
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 22545 24808 23054
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24780 22098 24808 22374
rect 24872 22166 24900 22374
rect 25056 22216 25084 22714
rect 25148 22409 25176 22986
rect 25332 22982 25360 24074
rect 25780 23792 25832 23798
rect 25780 23734 25832 23740
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25320 22976 25372 22982
rect 25318 22944 25320 22953
rect 25372 22944 25374 22953
rect 25318 22879 25374 22888
rect 25134 22400 25190 22409
rect 25134 22335 25190 22344
rect 25136 22228 25188 22234
rect 25056 22188 25136 22216
rect 25136 22170 25188 22176
rect 24860 22160 24912 22166
rect 24858 22128 24860 22137
rect 24912 22128 24914 22137
rect 24768 22092 24820 22098
rect 25148 22098 25176 22170
rect 24858 22063 24914 22072
rect 25136 22092 25188 22098
rect 24768 22034 24820 22040
rect 25136 22034 25188 22040
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 24952 22024 25004 22030
rect 24858 21992 24914 22001
rect 24688 21962 24808 21978
rect 24584 21956 24636 21962
rect 24688 21956 24820 21962
rect 24688 21950 24768 21956
rect 24584 21898 24636 21904
rect 24952 21966 25004 21972
rect 24858 21927 24914 21936
rect 24768 21898 24820 21904
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 23940 21072 23992 21078
rect 23940 21014 23992 21020
rect 23754 20904 23810 20913
rect 23572 20868 23624 20874
rect 23754 20839 23810 20848
rect 23572 20810 23624 20816
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 22848 20216 22968 20244
rect 22848 19922 22876 20216
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23018 19952 23074 19961
rect 22836 19916 22888 19922
rect 23018 19887 23074 19896
rect 23480 19916 23532 19922
rect 22836 19858 22888 19864
rect 23032 19854 23060 19887
rect 23480 19858 23532 19864
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22388 19638 22600 19666
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22020 17632 22140 17660
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22008 17128 22060 17134
rect 21928 17088 22008 17116
rect 21824 17070 21876 17076
rect 22008 17070 22060 17076
rect 21836 16794 21864 17070
rect 21732 16788 21784 16794
rect 21732 16730 21784 16736
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21560 15910 21588 16118
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21192 15524 21312 15552
rect 21364 15564 21416 15570
rect 21192 15094 21220 15524
rect 21364 15506 21416 15512
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21284 14958 21312 15370
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 21100 14482 21128 14826
rect 21376 14482 21404 15506
rect 21454 15464 21510 15473
rect 21454 15399 21510 15408
rect 21468 15366 21496 15399
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21468 14890 21496 15098
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21178 14376 21234 14385
rect 21178 14311 21234 14320
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21192 13258 21220 14311
rect 21376 14074 21404 14418
rect 21468 14346 21496 14418
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21560 14278 21588 15846
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21272 13184 21324 13190
rect 21192 13132 21272 13138
rect 21192 13126 21324 13132
rect 21192 13110 21312 13126
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21008 11830 21036 12174
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 21192 11234 21220 13110
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21284 11830 21312 12582
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21376 11694 21404 13330
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21560 12442 21588 12650
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21652 11558 21680 13194
rect 21744 13190 21772 16730
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21836 15473 21864 15846
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 21822 15464 21878 15473
rect 21928 15434 21956 15574
rect 21822 15399 21878 15408
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21836 14006 21864 14282
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21928 13870 21956 14894
rect 22020 14657 22048 17070
rect 22006 14648 22062 14657
rect 22006 14583 22062 14592
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 22112 13530 22140 17478
rect 22204 17202 22232 17682
rect 22388 17377 22416 19638
rect 22664 19378 22692 19654
rect 23492 19446 23520 19858
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22480 18222 22508 18906
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22572 17882 22600 19314
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22374 17368 22430 17377
rect 22374 17303 22430 17312
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22388 15450 22416 17303
rect 22664 16810 22692 19178
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 22756 17354 22784 18634
rect 23308 18426 23336 19314
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23308 18290 23336 18362
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22848 17785 22876 18022
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22834 17776 22890 17785
rect 22834 17711 22890 17720
rect 22756 17326 22876 17354
rect 22848 17270 22876 17326
rect 22836 17264 22888 17270
rect 22836 17206 22888 17212
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22572 16782 22692 16810
rect 22572 16674 22600 16782
rect 22480 16658 22600 16674
rect 22468 16652 22600 16658
rect 22520 16646 22600 16652
rect 22468 16594 22520 16600
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22480 15638 22508 15846
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22388 15422 22508 15450
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21730 12880 21786 12889
rect 22204 12850 22232 15302
rect 22374 15192 22430 15201
rect 22374 15127 22430 15136
rect 22388 14822 22416 15127
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22480 14362 22508 15422
rect 22572 14521 22600 16458
rect 22664 14906 22692 16782
rect 22756 16658 22784 17138
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16794 23336 18226
rect 23492 17678 23520 18634
rect 23584 17882 23612 20810
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23768 18154 23796 20470
rect 23846 19952 23902 19961
rect 23846 19887 23848 19896
rect 23900 19887 23902 19896
rect 23848 19858 23900 19864
rect 23952 19514 23980 21014
rect 24136 20942 24164 21082
rect 24216 21004 24268 21010
rect 24216 20946 24268 20952
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 24228 20534 24256 20946
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24228 19446 24256 20470
rect 24596 19922 24624 21898
rect 24872 21894 24900 21927
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24688 20398 24716 21830
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 24308 19916 24360 19922
rect 24308 19858 24360 19864
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24320 19514 24348 19858
rect 24308 19508 24360 19514
rect 24308 19450 24360 19456
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23860 18698 23888 19110
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 24136 18358 24164 18702
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23662 18048 23718 18057
rect 23662 17983 23718 17992
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23492 17338 23520 17614
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23676 17241 23704 17983
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23662 17232 23718 17241
rect 23662 17167 23718 17176
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 22664 14878 22784 14906
rect 22848 14890 22876 16390
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23308 15570 23336 16390
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22558 14512 22614 14521
rect 22558 14447 22614 14456
rect 22480 14334 22600 14362
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 21730 12815 21786 12824
rect 21916 12844 21968 12850
rect 21744 12238 21772 12815
rect 21916 12786 21968 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21192 11206 21864 11234
rect 20812 11144 20864 11150
rect 20732 11104 20812 11132
rect 20732 10130 20760 11104
rect 20812 11086 20864 11092
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 20996 10736 21048 10742
rect 21652 10724 21680 11018
rect 21048 10696 21680 10724
rect 20996 10678 21048 10684
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 21100 10130 21128 10542
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21100 9722 21128 10066
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21284 9654 21312 10474
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21836 9382 21864 11206
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21468 8430 21496 8910
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21468 7886 21496 8366
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4554 19104 5102
rect 19260 4690 19288 6598
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 19076 3058 19104 4490
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19352 3194 19380 3402
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17420 2446 17448 2790
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 15948 800 15976 2314
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 2926
rect 19444 2446 19472 6054
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 2514 20024 4558
rect 20640 3058 20668 4966
rect 20732 4826 20760 7210
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 21008 3534 21036 7754
rect 21456 7744 21508 7750
rect 21560 7698 21588 9318
rect 21508 7692 21588 7698
rect 21456 7686 21588 7692
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21468 7670 21588 7686
rect 21468 7206 21496 7670
rect 21652 7274 21680 7686
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21744 4690 21772 6598
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21836 4486 21864 9318
rect 21928 8090 21956 12786
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22020 11762 22048 12718
rect 22112 12306 22140 12718
rect 22480 12442 22508 13398
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22374 12200 22430 12209
rect 22374 12135 22376 12144
rect 22428 12135 22430 12144
rect 22468 12164 22520 12170
rect 22376 12106 22428 12112
rect 22468 12106 22520 12112
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22388 11694 22416 12106
rect 22480 12073 22508 12106
rect 22466 12064 22522 12073
rect 22466 11999 22522 12008
rect 22572 11880 22600 14334
rect 22664 12986 22692 14758
rect 22756 14550 22784 14878
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22756 13530 22784 14486
rect 23124 13734 23152 14554
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22480 11852 22600 11880
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11014 22048 11494
rect 22480 11121 22508 11852
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22466 11112 22522 11121
rect 22466 11047 22522 11056
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22020 10690 22048 10950
rect 22284 10736 22336 10742
rect 22020 10662 22232 10690
rect 22284 10678 22336 10684
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10062 22048 10542
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22020 8974 22048 9998
rect 22112 9178 22140 10406
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22020 7206 22048 8434
rect 22112 8430 22140 9114
rect 22204 8922 22232 10662
rect 22296 9722 22324 10678
rect 22572 9994 22600 11698
rect 22664 11626 22692 12786
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22664 10810 22692 10950
rect 22848 10826 22876 13194
rect 22926 13016 22982 13025
rect 23032 12986 23060 13330
rect 22926 12951 22928 12960
rect 22980 12951 22982 12960
rect 23020 12980 23072 12986
rect 22928 12922 22980 12928
rect 23020 12922 23072 12928
rect 22940 12714 22968 12922
rect 22928 12708 22980 12714
rect 22928 12650 22980 12656
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11354 23336 14962
rect 23400 12714 23428 15982
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23492 12374 23520 16050
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23584 12782 23612 14894
rect 23676 13530 23704 16390
rect 23768 15162 23796 17478
rect 24136 17270 24164 18294
rect 24124 17264 24176 17270
rect 24124 17206 24176 17212
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 24596 16046 24624 17002
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 23848 15632 23900 15638
rect 23848 15574 23900 15580
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23860 14929 23888 15574
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 23952 15026 23980 15506
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23846 14920 23902 14929
rect 23846 14855 23902 14864
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23860 13410 23888 14214
rect 24044 14006 24072 15506
rect 24688 14958 24716 20334
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24872 19310 24900 20198
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24780 17610 24808 18566
rect 24872 17746 24900 19246
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24780 16182 24808 17546
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24872 15978 24900 17478
rect 24964 17338 24992 21966
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25148 21049 25176 21490
rect 25134 21040 25190 21049
rect 25134 20975 25190 20984
rect 25240 20874 25268 22034
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25412 21480 25464 21486
rect 25412 21422 25464 21428
rect 25228 20868 25280 20874
rect 25228 20810 25280 20816
rect 25332 20312 25360 21422
rect 25424 20641 25452 21422
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25410 20632 25466 20641
rect 25410 20567 25466 20576
rect 25332 20284 25452 20312
rect 25318 20224 25374 20233
rect 25318 20159 25374 20168
rect 25332 19938 25360 20159
rect 25148 19910 25360 19938
rect 25148 19825 25176 19910
rect 25228 19848 25280 19854
rect 25134 19816 25190 19825
rect 25228 19790 25280 19796
rect 25134 19751 25190 19760
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 25056 19145 25084 19654
rect 25042 19136 25098 19145
rect 25042 19071 25098 19080
rect 25148 18850 25176 19751
rect 25240 19514 25268 19790
rect 25332 19718 25360 19910
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25056 18834 25176 18850
rect 25044 18828 25176 18834
rect 25096 18822 25176 18828
rect 25044 18770 25096 18776
rect 25134 18320 25190 18329
rect 25044 18284 25096 18290
rect 25134 18255 25136 18264
rect 25044 18226 25096 18232
rect 25188 18255 25190 18264
rect 25136 18226 25188 18232
rect 25056 18193 25084 18226
rect 25240 18222 25268 19450
rect 25228 18216 25280 18222
rect 25042 18184 25098 18193
rect 25228 18158 25280 18164
rect 25042 18119 25098 18128
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17746 25084 18022
rect 25228 17808 25280 17814
rect 25228 17750 25280 17756
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 25240 16590 25268 17750
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24964 16425 24992 16458
rect 24950 16416 25006 16425
rect 24950 16351 25006 16360
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 25240 15366 25268 16526
rect 25332 16454 25360 19654
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24596 14618 24624 14894
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23676 13382 23888 13410
rect 23676 13258 23704 13382
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 22848 10810 22968 10826
rect 22652 10804 22704 10810
rect 22848 10804 22980 10810
rect 22848 10798 22928 10804
rect 22652 10746 22704 10752
rect 22928 10746 22980 10752
rect 23584 10742 23612 10950
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23400 9994 23428 10610
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 22572 9722 22600 9930
rect 23584 9926 23612 10474
rect 23676 10266 23704 12922
rect 23860 12918 23888 13126
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23860 12170 23888 12718
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 23756 11280 23808 11286
rect 23756 11222 23808 11228
rect 23768 10470 23796 11222
rect 23848 11212 23900 11218
rect 23848 11154 23900 11160
rect 23860 11121 23888 11154
rect 23846 11112 23902 11121
rect 23952 11082 23980 13806
rect 24412 13394 24440 14214
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24400 13388 24452 13394
rect 24400 13330 24452 13336
rect 24044 12646 24072 13330
rect 24596 12986 24624 13738
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24688 13326 24716 13670
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 24044 12434 24072 12582
rect 24044 12406 24164 12434
rect 23846 11047 23902 11056
rect 23940 11076 23992 11082
rect 23860 11014 23888 11047
rect 23940 11018 23992 11024
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22204 8894 22324 8922
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22204 7886 22232 8774
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22296 7546 22324 8894
rect 22468 8356 22520 8362
rect 22520 8316 22600 8344
rect 22468 8298 22520 8304
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22388 7410 22416 7686
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 21008 2990 21036 3470
rect 21284 3058 21312 4422
rect 21376 4282 21404 4422
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 22020 3738 22048 7142
rect 22388 6866 22416 7346
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22112 4214 22140 4558
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22020 3466 22048 3674
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21376 2854 21404 3402
rect 22112 3126 22140 4150
rect 22100 3120 22152 3126
rect 22152 3068 22232 3074
rect 22100 3062 22232 3068
rect 22112 3046 22232 3062
rect 22204 2922 22232 3046
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20180 800 20208 2450
rect 22112 2446 22140 2858
rect 22480 2582 22508 7686
rect 22572 7342 22600 8316
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22664 7274 22692 9522
rect 23768 9466 23796 10406
rect 23860 10130 23888 10950
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23952 9926 23980 10542
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23676 9438 23796 9466
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23676 7954 23704 9438
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 9042 23796 9318
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 22652 7268 22704 7274
rect 22652 7210 22704 7216
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23952 6186 23980 9862
rect 24044 9042 24072 9998
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24044 8498 24072 8978
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 22940 4146 22968 4626
rect 23216 4146 23244 4626
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22848 3602 22876 3878
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22756 2922 22784 3334
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 23308 2854 23336 4014
rect 23584 3738 23612 4558
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 24136 3534 24164 12406
rect 24596 12238 24624 12922
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11830 24256 12038
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 24596 11558 24624 12174
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11150 24624 11494
rect 24584 11144 24636 11150
rect 24636 11092 24716 11098
rect 24584 11086 24716 11092
rect 24596 11070 24716 11086
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24504 10606 24532 10950
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24400 9988 24452 9994
rect 24400 9930 24452 9936
rect 24412 9654 24440 9930
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24412 9042 24440 9590
rect 24504 9518 24532 10202
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24596 9178 24624 9658
rect 24688 9654 24716 11070
rect 24780 10470 24808 15098
rect 25240 15026 25268 15302
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24872 14618 24900 14894
rect 24964 14822 24992 14962
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 24872 12918 24900 13398
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24872 11694 24900 12242
rect 24964 11801 24992 14758
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25148 13326 25176 14214
rect 25332 14074 25360 15506
rect 25424 14822 25452 20284
rect 25608 20262 25636 20946
rect 25700 20602 25728 23054
rect 25792 22710 25820 23734
rect 25780 22704 25832 22710
rect 25780 22646 25832 22652
rect 25792 22574 25820 22646
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25792 22438 25820 22510
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25884 22094 25912 24822
rect 25976 22522 26004 24890
rect 26068 23474 26096 24890
rect 26160 24188 26188 26302
rect 26698 26302 27016 26330
rect 26698 26200 26754 26302
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 26436 24410 26464 24618
rect 26332 24404 26384 24410
rect 26332 24346 26384 24352
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26240 24200 26292 24206
rect 26160 24160 26240 24188
rect 26240 24142 26292 24148
rect 26068 23446 26188 23474
rect 25976 22494 26096 22522
rect 25792 22066 25912 22094
rect 25792 22001 25820 22066
rect 25872 22024 25924 22030
rect 25778 21992 25834 22001
rect 25872 21966 25924 21972
rect 25778 21927 25834 21936
rect 25792 21690 25820 21927
rect 25780 21684 25832 21690
rect 25780 21626 25832 21632
rect 25778 21040 25834 21049
rect 25778 20975 25834 20984
rect 25792 20806 25820 20975
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25700 19378 25728 20538
rect 25792 19990 25820 20538
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25700 18834 25728 19314
rect 25884 19242 25912 21966
rect 26068 21146 26096 22494
rect 26160 21554 26188 23446
rect 26344 23168 26372 24346
rect 26436 24274 26464 24346
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 26606 24168 26662 24177
rect 26606 24103 26608 24112
rect 26660 24103 26662 24112
rect 26608 24074 26660 24080
rect 26988 24070 27016 26302
rect 27342 26200 27398 27000
rect 27986 26330 28042 27000
rect 27986 26302 28396 26330
rect 27986 26200 28042 26302
rect 27252 24744 27304 24750
rect 27252 24686 27304 24692
rect 27264 24410 27292 24686
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 27356 24274 27384 26200
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27252 24132 27304 24138
rect 27252 24074 27304 24080
rect 27344 24132 27396 24138
rect 27344 24074 27396 24080
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 26344 23140 26556 23168
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26252 22778 26280 22986
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26344 22710 26372 22918
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26528 22094 26556 23140
rect 26620 22778 26648 23598
rect 26700 23180 26752 23186
rect 26700 23122 26752 23128
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26620 22642 26648 22714
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26712 22234 26740 23122
rect 27264 23050 27292 24074
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 27264 22438 27292 22986
rect 27356 22506 27384 24074
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27632 22574 27660 23734
rect 27816 23730 27844 24006
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27816 23254 27844 23666
rect 28368 23662 28396 26302
rect 28630 26200 28686 27000
rect 29274 26330 29330 27000
rect 29274 26302 29592 26330
rect 29274 26200 29330 26302
rect 28644 24342 28672 26200
rect 29564 24750 29592 26302
rect 29918 26200 29974 27000
rect 30562 26330 30618 27000
rect 30562 26302 30880 26330
rect 30562 26200 30618 26302
rect 29932 24818 29960 26200
rect 29920 24812 29972 24818
rect 29920 24754 29972 24760
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30668 24614 30696 24686
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 28632 24336 28684 24342
rect 28632 24278 28684 24284
rect 30392 24206 30420 24550
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28632 24064 28684 24070
rect 28632 24006 28684 24012
rect 28356 23656 28408 23662
rect 28356 23598 28408 23604
rect 28356 23520 28408 23526
rect 28356 23462 28408 23468
rect 27804 23248 27856 23254
rect 27804 23190 27856 23196
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27344 22500 27396 22506
rect 27344 22442 27396 22448
rect 27436 22500 27488 22506
rect 27436 22442 27488 22448
rect 27252 22432 27304 22438
rect 27252 22374 27304 22380
rect 26700 22228 26752 22234
rect 26700 22170 26752 22176
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 26252 22066 26556 22094
rect 26606 22128 26662 22137
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 26252 21350 26280 22066
rect 26606 22063 26608 22072
rect 26660 22063 26662 22072
rect 26608 22034 26660 22040
rect 26422 21448 26478 21457
rect 26422 21383 26424 21392
rect 26476 21383 26478 21392
rect 26884 21412 26936 21418
rect 26424 21354 26476 21360
rect 26884 21354 26936 21360
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26056 21140 26108 21146
rect 26056 21082 26108 21088
rect 26068 20466 26096 21082
rect 26160 20992 26188 21286
rect 26516 21072 26568 21078
rect 26516 21014 26568 21020
rect 26332 21004 26384 21010
rect 26160 20964 26332 20992
rect 26332 20946 26384 20952
rect 26528 20806 26556 21014
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 26148 20392 26200 20398
rect 26054 20360 26110 20369
rect 26148 20334 26200 20340
rect 26054 20295 26056 20304
rect 26108 20295 26110 20304
rect 26056 20266 26108 20272
rect 26068 19514 26096 20266
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25792 18426 25820 19110
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25962 18320 26018 18329
rect 25962 18255 26018 18264
rect 25976 17270 26004 18255
rect 26056 18148 26108 18154
rect 26056 18090 26108 18096
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25516 14618 25544 17070
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25516 14074 25544 14554
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25332 12918 25360 14010
rect 25608 13530 25636 17138
rect 25976 16697 26004 17206
rect 26068 16726 26096 18090
rect 26056 16720 26108 16726
rect 25962 16688 26018 16697
rect 25688 16652 25740 16658
rect 26056 16662 26108 16668
rect 25962 16623 26018 16632
rect 25688 16594 25740 16600
rect 25700 13734 25728 16594
rect 25962 16552 26018 16561
rect 25962 16487 26018 16496
rect 25780 16176 25832 16182
rect 25780 16118 25832 16124
rect 25792 14346 25820 16118
rect 25976 15434 26004 16487
rect 26160 16454 26188 20334
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 26528 19446 26556 20198
rect 26804 20058 26832 20810
rect 26896 20534 26924 21354
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 20806 27016 21286
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 27068 20800 27120 20806
rect 27068 20742 27120 20748
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26896 19922 26924 20470
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26712 19446 26740 19654
rect 26516 19440 26568 19446
rect 26516 19382 26568 19388
rect 26700 19440 26752 19446
rect 26700 19382 26752 19388
rect 26424 18216 26476 18222
rect 26238 18184 26294 18193
rect 26424 18158 26476 18164
rect 26238 18119 26294 18128
rect 26252 17882 26280 18119
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26252 16998 26280 17818
rect 26436 17202 26464 18158
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 26148 16448 26200 16454
rect 26240 16448 26292 16454
rect 26148 16390 26200 16396
rect 26238 16416 26240 16425
rect 26292 16416 26294 16425
rect 26238 16351 26294 16360
rect 26148 16176 26200 16182
rect 26252 16164 26280 16351
rect 26200 16136 26280 16164
rect 26148 16118 26200 16124
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 26068 15706 26096 15982
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25884 15094 25912 15302
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25976 15026 26004 15370
rect 26238 15056 26294 15065
rect 25964 15020 26016 15026
rect 26238 14991 26240 15000
rect 25964 14962 26016 14968
rect 26292 14991 26294 15000
rect 26240 14962 26292 14968
rect 25780 14340 25832 14346
rect 25780 14282 25832 14288
rect 25792 14006 25820 14282
rect 25780 14000 25832 14006
rect 25780 13942 25832 13948
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25792 13530 25820 13942
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 25792 12986 25820 13466
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25332 12434 25360 12854
rect 25240 12406 25360 12434
rect 24950 11792 25006 11801
rect 24950 11727 25006 11736
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24872 11218 24900 11630
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24964 11098 24992 11727
rect 25240 11354 25268 12406
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25884 11830 25912 12174
rect 25872 11824 25924 11830
rect 25872 11766 25924 11772
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 24872 11070 24992 11098
rect 25884 11082 25912 11766
rect 25872 11076 25924 11082
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24412 8906 24440 8978
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24412 8634 24440 8842
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24872 4078 24900 11070
rect 25872 11018 25924 11024
rect 25884 10810 25912 11018
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25780 9988 25832 9994
rect 25884 9976 25912 10746
rect 25832 9948 25912 9976
rect 25780 9930 25832 9936
rect 25608 9042 25636 9930
rect 25976 9602 26004 14962
rect 26344 14618 26372 15370
rect 26424 15360 26476 15366
rect 26424 15302 26476 15308
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 26068 12889 26096 13194
rect 26436 13025 26464 15302
rect 26528 14618 26556 19382
rect 26988 19378 27016 20742
rect 27080 20602 27108 20742
rect 27068 20596 27120 20602
rect 27068 20538 27120 20544
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 27080 19718 27108 19994
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 26792 18624 26844 18630
rect 26792 18566 26844 18572
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26712 16114 26740 16390
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26516 14612 26568 14618
rect 26516 14554 26568 14560
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26422 13016 26478 13025
rect 26528 12986 26556 13126
rect 26422 12951 26424 12960
rect 26476 12951 26478 12960
rect 26516 12980 26568 12986
rect 26424 12922 26476 12928
rect 26516 12922 26568 12928
rect 26054 12880 26110 12889
rect 26054 12815 26110 12824
rect 26056 12776 26108 12782
rect 26056 12718 26108 12724
rect 25884 9574 26004 9602
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25700 8838 25728 9386
rect 25884 9382 25912 9574
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25976 9178 26004 9454
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25700 7750 25728 8774
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25700 6186 25728 7686
rect 26068 6644 26096 12718
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26344 12102 26372 12310
rect 26332 12096 26384 12102
rect 26332 12038 26384 12044
rect 26148 11824 26200 11830
rect 26148 11766 26200 11772
rect 26160 10742 26188 11766
rect 26620 11354 26648 15506
rect 26712 12442 26740 15846
rect 26804 15706 26832 18566
rect 26884 17060 26936 17066
rect 26884 17002 26936 17008
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26804 12782 26832 15642
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26896 12306 26924 17002
rect 26988 16522 27016 19314
rect 27080 18086 27108 19654
rect 27172 18970 27200 22170
rect 27448 22030 27476 22442
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27448 20942 27476 21626
rect 27436 20936 27488 20942
rect 27434 20904 27436 20913
rect 27488 20904 27490 20913
rect 27434 20839 27490 20848
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27264 19378 27292 19654
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27160 18964 27212 18970
rect 27160 18906 27212 18912
rect 27264 18426 27292 19110
rect 27540 18834 27568 22034
rect 27620 22024 27672 22030
rect 27618 21992 27620 22001
rect 27672 21992 27674 22001
rect 27618 21927 27674 21936
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27632 20754 27660 21830
rect 27724 20874 27752 22578
rect 27816 21690 27844 22646
rect 28080 22568 28132 22574
rect 28080 22510 28132 22516
rect 27896 22432 27948 22438
rect 27896 22374 27948 22380
rect 27908 22234 27936 22374
rect 27896 22228 27948 22234
rect 27896 22170 27948 22176
rect 28092 22098 28120 22510
rect 28262 22264 28318 22273
rect 28262 22199 28318 22208
rect 28276 22166 28304 22199
rect 28264 22160 28316 22166
rect 28264 22102 28316 22108
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 28368 21962 28396 23462
rect 28356 21956 28408 21962
rect 28356 21898 28408 21904
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27908 21010 27936 21490
rect 27896 21004 27948 21010
rect 27896 20946 27948 20952
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 27632 20726 27752 20754
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27528 18828 27580 18834
rect 27528 18770 27580 18776
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27528 18692 27580 18698
rect 27528 18634 27580 18640
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27068 17196 27120 17202
rect 27068 17138 27120 17144
rect 26976 16516 27028 16522
rect 26976 16458 27028 16464
rect 26974 15464 27030 15473
rect 26974 15399 27030 15408
rect 26988 15366 27016 15399
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 27080 14346 27108 17138
rect 27172 15502 27200 18022
rect 27448 17678 27476 18634
rect 27540 18426 27568 18634
rect 27528 18420 27580 18426
rect 27528 18362 27580 18368
rect 27632 18306 27660 19654
rect 27724 19009 27752 20726
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28446 19952 28502 19961
rect 28356 19916 28408 19922
rect 28446 19887 28502 19896
rect 28356 19858 28408 19864
rect 27804 19780 27856 19786
rect 27804 19722 27856 19728
rect 27710 19000 27766 19009
rect 27710 18935 27766 18944
rect 27712 18828 27764 18834
rect 27712 18770 27764 18776
rect 27724 18426 27752 18770
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27540 18290 27660 18306
rect 27528 18284 27660 18290
rect 27580 18278 27660 18284
rect 27528 18226 27580 18232
rect 27712 18216 27764 18222
rect 27540 18164 27712 18170
rect 27540 18158 27764 18164
rect 27540 18142 27752 18158
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27252 17604 27304 17610
rect 27252 17546 27304 17552
rect 27264 16708 27292 17546
rect 27344 16720 27396 16726
rect 27264 16680 27344 16708
rect 27264 16232 27292 16680
rect 27344 16662 27396 16668
rect 27448 16454 27476 17614
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27264 16204 27384 16232
rect 27250 16144 27306 16153
rect 27356 16114 27384 16204
rect 27250 16079 27306 16088
rect 27344 16108 27396 16114
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27264 15434 27292 16079
rect 27344 16050 27396 16056
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27264 15162 27292 15370
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27250 15056 27306 15065
rect 27250 14991 27252 15000
rect 27304 14991 27306 15000
rect 27252 14962 27304 14968
rect 27160 14952 27212 14958
rect 27160 14894 27212 14900
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27080 13870 27108 14282
rect 27068 13864 27120 13870
rect 27068 13806 27120 13812
rect 27080 13394 27108 13806
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 27068 12980 27120 12986
rect 27068 12922 27120 12928
rect 27080 12434 27108 12922
rect 26988 12406 27108 12434
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26988 12102 27016 12406
rect 27068 12300 27120 12306
rect 27068 12242 27120 12248
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26976 11824 27028 11830
rect 26976 11766 27028 11772
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 26148 10736 26200 10742
rect 26148 10678 26200 10684
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26344 10266 26372 10610
rect 26620 10606 26648 11290
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26620 10198 26648 10542
rect 26712 10198 26740 10746
rect 26608 10192 26660 10198
rect 26608 10134 26660 10140
rect 26700 10192 26752 10198
rect 26700 10134 26752 10140
rect 26712 9926 26740 10134
rect 26896 10130 26924 11086
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 25792 6616 26096 6644
rect 25688 6180 25740 6186
rect 25688 6122 25740 6128
rect 25792 4078 25820 6616
rect 26988 6254 27016 11766
rect 27080 11064 27108 12242
rect 27172 11694 27200 14894
rect 27356 12374 27384 15914
rect 27540 15638 27568 18142
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27632 17542 27660 18022
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27632 16658 27660 17478
rect 27710 17368 27766 17377
rect 27816 17338 27844 19722
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28368 19514 28396 19858
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28460 19378 28488 19887
rect 28172 19372 28224 19378
rect 28172 19314 28224 19320
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 28000 18902 28028 19246
rect 27988 18896 28040 18902
rect 27988 18838 28040 18844
rect 28000 18630 28028 18838
rect 28184 18630 28212 19314
rect 28356 19304 28408 19310
rect 28408 19252 28488 19258
rect 28356 19246 28488 19252
rect 28368 19230 28488 19246
rect 28552 19242 28580 24006
rect 28644 19854 28672 24006
rect 29932 23905 29960 24142
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 29918 23896 29974 23905
rect 29918 23831 29974 23840
rect 30010 23760 30066 23769
rect 30010 23695 30066 23704
rect 30380 23724 30432 23730
rect 29184 23656 29236 23662
rect 29104 23616 29184 23644
rect 29104 22250 29132 23616
rect 29184 23598 29236 23604
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29368 23520 29420 23526
rect 29368 23462 29420 23468
rect 29276 23180 29328 23186
rect 29276 23122 29328 23128
rect 29288 22710 29316 23122
rect 29276 22704 29328 22710
rect 29276 22646 29328 22652
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 29196 22386 29224 22510
rect 29196 22358 29316 22386
rect 29000 22228 29052 22234
rect 29104 22222 29224 22250
rect 29000 22170 29052 22176
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 28828 21593 28856 21626
rect 28814 21584 28870 21593
rect 28814 21519 28870 21528
rect 28920 21486 28948 22034
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 29012 21298 29040 22170
rect 29196 22098 29224 22222
rect 29184 22092 29236 22098
rect 29184 22034 29236 22040
rect 29184 21888 29236 21894
rect 29184 21830 29236 21836
rect 28920 21270 29040 21298
rect 28724 20800 28776 20806
rect 28724 20742 28776 20748
rect 28632 19848 28684 19854
rect 28632 19790 28684 19796
rect 28736 19514 28764 20742
rect 28920 20534 28948 21270
rect 29196 20534 29224 21830
rect 28908 20528 28960 20534
rect 28908 20470 28960 20476
rect 29184 20528 29236 20534
rect 29184 20470 29236 20476
rect 29288 20398 29316 22358
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 28908 20324 28960 20330
rect 28908 20266 28960 20272
rect 28920 19990 28948 20266
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28816 19508 28868 19514
rect 28816 19450 28868 19456
rect 28354 18728 28410 18737
rect 28354 18663 28410 18672
rect 27988 18624 28040 18630
rect 27988 18566 28040 18572
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27710 17303 27712 17312
rect 27764 17303 27766 17312
rect 27804 17332 27856 17338
rect 27712 17274 27764 17280
rect 27804 17274 27856 17280
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 27804 17128 27856 17134
rect 27804 17070 27856 17076
rect 27986 17096 28042 17105
rect 27816 16726 27844 17070
rect 27986 17031 28042 17040
rect 28000 16998 28028 17031
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 27804 16720 27856 16726
rect 27804 16662 27856 16668
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 28000 16436 28028 16934
rect 28078 16688 28134 16697
rect 28276 16658 28304 17138
rect 28078 16623 28080 16632
rect 28132 16623 28134 16632
rect 28264 16652 28316 16658
rect 28080 16594 28132 16600
rect 28264 16594 28316 16600
rect 28276 16454 28304 16594
rect 27724 16408 28028 16436
rect 28264 16448 28316 16454
rect 27528 15632 27580 15638
rect 27528 15574 27580 15580
rect 27724 15502 27752 16408
rect 28264 16390 28316 16396
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27448 13326 27476 15302
rect 27526 15192 27582 15201
rect 27526 15127 27528 15136
rect 27580 15127 27582 15136
rect 27528 15098 27580 15104
rect 27540 14278 27568 15098
rect 27816 15026 27844 16118
rect 28368 15609 28396 18663
rect 28460 18630 28488 19230
rect 28540 19236 28592 19242
rect 28540 19178 28592 19184
rect 28538 19136 28594 19145
rect 28828 19122 28856 19450
rect 28920 19258 28948 19926
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 29000 19304 29052 19310
rect 28920 19252 29000 19258
rect 28920 19246 29052 19252
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 28920 19230 29040 19246
rect 29104 19122 29132 19246
rect 28594 19094 28856 19122
rect 28920 19094 29132 19122
rect 28538 19071 28594 19080
rect 28448 18624 28500 18630
rect 28448 18566 28500 18572
rect 28460 18193 28488 18566
rect 28446 18184 28502 18193
rect 28446 18119 28502 18128
rect 28448 17740 28500 17746
rect 28448 17682 28500 17688
rect 28354 15600 28410 15609
rect 28354 15535 28410 15544
rect 28368 15434 28396 15535
rect 28356 15428 28408 15434
rect 28356 15370 28408 15376
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 28460 15162 28488 17682
rect 28552 16658 28580 19071
rect 28630 19000 28686 19009
rect 28630 18935 28686 18944
rect 28644 16998 28672 18935
rect 28920 18902 28948 19094
rect 29092 18964 29144 18970
rect 29092 18906 29144 18912
rect 28908 18896 28960 18902
rect 29000 18896 29052 18902
rect 28908 18838 28960 18844
rect 28998 18864 29000 18873
rect 29052 18864 29054 18873
rect 28998 18799 29054 18808
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28828 17882 28856 18702
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 28828 17762 28856 17818
rect 28828 17734 29040 17762
rect 29104 17746 29132 18906
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28630 16824 28686 16833
rect 28828 16794 28856 17478
rect 28630 16759 28686 16768
rect 28816 16788 28868 16794
rect 28644 16658 28672 16759
rect 28816 16730 28868 16736
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28552 15892 28580 16594
rect 28632 16448 28684 16454
rect 28632 16390 28684 16396
rect 28644 16046 28672 16390
rect 28632 16040 28684 16046
rect 28684 16000 28764 16028
rect 28632 15982 28684 15988
rect 28632 15904 28684 15910
rect 28552 15864 28632 15892
rect 28632 15846 28684 15852
rect 28448 15156 28500 15162
rect 28448 15098 28500 15104
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 27988 14816 28040 14822
rect 27986 14784 27988 14793
rect 28040 14784 28042 14793
rect 27986 14719 28042 14728
rect 28736 14482 28764 16000
rect 27896 14476 27948 14482
rect 27896 14418 27948 14424
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 27620 14408 27672 14414
rect 27908 14362 27936 14418
rect 27620 14350 27672 14356
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27632 14090 27660 14350
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27816 14334 27936 14362
rect 27540 14074 27660 14090
rect 27528 14068 27660 14074
rect 27580 14062 27660 14068
rect 27528 14010 27580 14016
rect 27724 13530 27752 14282
rect 27816 13530 27844 14334
rect 28448 14272 28500 14278
rect 28500 14232 28580 14260
rect 28448 14214 28500 14220
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27540 12918 27568 13466
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27344 12368 27396 12374
rect 27344 12310 27396 12316
rect 27540 12238 27568 12854
rect 27528 12232 27580 12238
rect 27580 12192 27660 12220
rect 27528 12174 27580 12180
rect 27252 12096 27304 12102
rect 27252 12038 27304 12044
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27160 11688 27212 11694
rect 27160 11630 27212 11636
rect 27160 11076 27212 11082
rect 27080 11036 27160 11064
rect 27160 11018 27212 11024
rect 27068 10804 27120 10810
rect 27068 10746 27120 10752
rect 27080 10606 27108 10746
rect 27068 10600 27120 10606
rect 27068 10542 27120 10548
rect 27172 9518 27200 11018
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 27264 7750 27292 12038
rect 27356 11898 27384 12038
rect 27434 11928 27490 11937
rect 27344 11892 27396 11898
rect 27434 11863 27490 11872
rect 27344 11834 27396 11840
rect 27448 11694 27476 11863
rect 27632 11830 27660 12192
rect 27620 11824 27672 11830
rect 27620 11766 27672 11772
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27344 11620 27396 11626
rect 27344 11562 27396 11568
rect 27356 9994 27384 11562
rect 27448 10742 27476 11630
rect 27632 11082 27660 11766
rect 27724 11121 27752 13466
rect 27816 12646 27844 13466
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27804 12640 27856 12646
rect 27804 12582 27856 12588
rect 27908 12442 27936 12922
rect 27896 12436 27948 12442
rect 27896 12378 27948 12384
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27710 11112 27766 11121
rect 27620 11076 27672 11082
rect 27710 11047 27766 11056
rect 27620 11018 27672 11024
rect 27436 10736 27488 10742
rect 27436 10678 27488 10684
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27540 10282 27568 10610
rect 27724 10418 27752 11047
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27448 10266 27568 10282
rect 27436 10260 27568 10266
rect 27488 10254 27568 10260
rect 27436 10202 27488 10208
rect 27344 9988 27396 9994
rect 27344 9930 27396 9936
rect 27356 9654 27384 9930
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 27540 6390 27568 10254
rect 27632 10390 27752 10418
rect 27632 7410 27660 10390
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 27528 6384 27580 6390
rect 27528 6326 27580 6332
rect 27816 6322 27844 8774
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 28368 5234 28396 13466
rect 28552 12753 28580 14232
rect 28828 14074 28856 16730
rect 28920 16590 28948 17614
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 28920 16182 28948 16526
rect 28908 16176 28960 16182
rect 28908 16118 28960 16124
rect 29012 16046 29040 17734
rect 29092 17740 29144 17746
rect 29092 17682 29144 17688
rect 29196 17202 29224 19654
rect 29276 19168 29328 19174
rect 29276 19110 29328 19116
rect 29288 17338 29316 19110
rect 29380 18630 29408 23462
rect 29748 23322 29776 23530
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29460 23112 29512 23118
rect 29460 23054 29512 23060
rect 29472 22710 29500 23054
rect 29920 23044 29972 23050
rect 29920 22986 29972 22992
rect 29460 22704 29512 22710
rect 29460 22646 29512 22652
rect 29642 22672 29698 22681
rect 29472 22234 29500 22646
rect 29642 22607 29698 22616
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 29460 22092 29512 22098
rect 29460 22034 29512 22040
rect 29472 21622 29500 22034
rect 29460 21616 29512 21622
rect 29460 21558 29512 21564
rect 29472 18766 29500 21558
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29564 21078 29592 21286
rect 29656 21146 29684 22607
rect 29932 22574 29960 22986
rect 30024 22982 30052 23695
rect 30380 23666 30432 23672
rect 30196 23588 30248 23594
rect 30196 23530 30248 23536
rect 30208 23186 30236 23530
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23186 30328 23462
rect 30196 23180 30248 23186
rect 30196 23122 30248 23128
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30392 22982 30420 23666
rect 30012 22976 30064 22982
rect 30012 22918 30064 22924
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30380 22976 30432 22982
rect 30380 22918 30432 22924
rect 29920 22568 29972 22574
rect 29920 22510 29972 22516
rect 29734 22400 29790 22409
rect 29734 22335 29790 22344
rect 29748 21894 29776 22335
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29932 21729 29960 21966
rect 29918 21720 29974 21729
rect 30024 21690 30052 22170
rect 29918 21655 29974 21664
rect 30012 21684 30064 21690
rect 30012 21626 30064 21632
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29932 21418 29960 21490
rect 29920 21412 29972 21418
rect 29920 21354 29972 21360
rect 30024 21146 30052 21626
rect 29644 21140 29696 21146
rect 29644 21082 29696 21088
rect 30012 21140 30064 21146
rect 30012 21082 30064 21088
rect 29552 21072 29604 21078
rect 29828 21072 29880 21078
rect 29552 21014 29604 21020
rect 29748 21020 29828 21026
rect 29748 21014 29880 21020
rect 30010 21040 30066 21049
rect 29748 20998 29868 21014
rect 29552 20936 29604 20942
rect 29748 20924 29776 20998
rect 30010 20975 30066 20984
rect 29604 20896 29776 20924
rect 29920 20936 29972 20942
rect 29826 20904 29882 20913
rect 29552 20878 29604 20884
rect 29564 20398 29592 20878
rect 29920 20878 29972 20884
rect 29826 20839 29882 20848
rect 29552 20392 29604 20398
rect 29552 20334 29604 20340
rect 29564 19718 29592 20334
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29642 19544 29698 19553
rect 29642 19479 29698 19488
rect 29656 19446 29684 19479
rect 29644 19440 29696 19446
rect 29644 19382 29696 19388
rect 29552 18828 29604 18834
rect 29552 18770 29604 18776
rect 29460 18760 29512 18766
rect 29460 18702 29512 18708
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29276 17332 29328 17338
rect 29276 17274 29328 17280
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29288 16658 29316 17274
rect 29276 16652 29328 16658
rect 29276 16594 29328 16600
rect 29380 16522 29408 18566
rect 29460 16652 29512 16658
rect 29460 16594 29512 16600
rect 29368 16516 29420 16522
rect 29368 16458 29420 16464
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29380 15366 29408 15982
rect 29368 15360 29420 15366
rect 29368 15302 29420 15308
rect 29380 15026 29408 15302
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29276 14544 29328 14550
rect 29276 14486 29328 14492
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28538 12744 28594 12753
rect 28538 12679 28594 12688
rect 28736 11898 28764 13126
rect 28828 12170 28856 14010
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 28920 13530 28948 13874
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 29012 13326 29040 14214
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28908 12776 28960 12782
rect 28908 12718 28960 12724
rect 28816 12164 28868 12170
rect 28816 12106 28868 12112
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28828 11354 28856 12106
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 28828 10742 28856 11290
rect 28920 11286 28948 12718
rect 29288 11558 29316 14486
rect 29276 11552 29328 11558
rect 29276 11494 29328 11500
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28816 10736 28868 10742
rect 28816 10678 28868 10684
rect 28828 9722 28856 10678
rect 28920 9926 28948 11086
rect 29288 11082 29316 11494
rect 29276 11076 29328 11082
rect 29276 11018 29328 11024
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 28908 9920 28960 9926
rect 28908 9862 28960 9868
rect 28920 9722 28948 9862
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 29104 8566 29132 10202
rect 29288 10198 29316 11018
rect 29276 10192 29328 10198
rect 29276 10134 29328 10140
rect 29276 9512 29328 9518
rect 29196 9460 29276 9466
rect 29196 9454 29328 9460
rect 29196 9438 29316 9454
rect 29472 9450 29500 16594
rect 29564 15026 29592 18770
rect 29656 17882 29684 19382
rect 29748 18426 29776 19654
rect 29840 19122 29868 20839
rect 29932 19281 29960 20878
rect 30024 19922 30052 20975
rect 30116 20806 30144 22918
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30196 22228 30248 22234
rect 30196 22170 30248 22176
rect 30208 22001 30236 22170
rect 30194 21992 30250 22001
rect 30484 21962 30512 22714
rect 30576 22098 30604 24006
rect 30852 23322 30880 26302
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26200 33838 27000
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26330 37058 27000
rect 37646 26330 37702 27000
rect 38290 26330 38346 27000
rect 37002 26302 37136 26330
rect 37002 26200 37058 26302
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 30840 23316 30892 23322
rect 30840 23258 30892 23264
rect 31036 23186 31064 24550
rect 31114 23760 31170 23769
rect 31114 23695 31170 23704
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 30654 22672 30710 22681
rect 30654 22607 30656 22616
rect 30708 22607 30710 22616
rect 30656 22578 30708 22584
rect 31024 22500 31076 22506
rect 31024 22442 31076 22448
rect 31036 22216 31064 22442
rect 30760 22188 31064 22216
rect 30564 22092 30616 22098
rect 30760 22094 30788 22188
rect 31128 22148 31156 23695
rect 31220 22982 31248 26200
rect 31576 24336 31628 24342
rect 31864 24313 31892 26200
rect 32508 24857 32536 26200
rect 32494 24848 32550 24857
rect 32494 24783 32550 24792
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32496 24608 32548 24614
rect 32496 24550 32548 24556
rect 31576 24278 31628 24284
rect 31850 24304 31906 24313
rect 31300 23248 31352 23254
rect 31300 23190 31352 23196
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 30564 22034 30616 22040
rect 30668 22066 30788 22094
rect 30194 21927 30250 21936
rect 30472 21956 30524 21962
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30208 20466 30236 21927
rect 30472 21898 30524 21904
rect 30576 21894 30604 22034
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30392 21593 30420 21830
rect 30668 21706 30696 22066
rect 30760 21962 30788 22066
rect 31036 22120 31156 22148
rect 30840 22024 30892 22030
rect 30840 21966 30892 21972
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30576 21678 30696 21706
rect 30378 21584 30434 21593
rect 30378 21519 30434 21528
rect 30472 21480 30524 21486
rect 30472 21422 30524 21428
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30012 19916 30064 19922
rect 30012 19858 30064 19864
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30288 19916 30340 19922
rect 30288 19858 30340 19864
rect 30104 19848 30156 19854
rect 30024 19796 30104 19802
rect 30024 19790 30156 19796
rect 30024 19774 30144 19790
rect 29918 19272 29974 19281
rect 29918 19207 29974 19216
rect 30024 19156 30052 19774
rect 30104 19712 30156 19718
rect 30104 19654 30156 19660
rect 30116 19417 30144 19654
rect 30102 19408 30158 19417
rect 30102 19343 30158 19352
rect 30104 19168 30156 19174
rect 30024 19136 30104 19156
rect 30156 19136 30158 19145
rect 30024 19128 30102 19136
rect 29840 19094 29960 19122
rect 29932 18834 29960 19094
rect 30102 19071 30158 19080
rect 30104 18896 30156 18902
rect 30010 18864 30066 18873
rect 29920 18828 29972 18834
rect 30104 18838 30156 18844
rect 30010 18799 30066 18808
rect 29920 18770 29972 18776
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29828 18420 29880 18426
rect 29828 18362 29880 18368
rect 29840 18170 29868 18362
rect 29748 18142 29868 18170
rect 29748 18086 29776 18142
rect 29736 18080 29788 18086
rect 29736 18022 29788 18028
rect 29644 17876 29696 17882
rect 29644 17818 29696 17824
rect 29656 17270 29684 17818
rect 29644 17264 29696 17270
rect 29644 17206 29696 17212
rect 29642 16008 29698 16017
rect 29642 15943 29698 15952
rect 29552 15020 29604 15026
rect 29552 14962 29604 14968
rect 29564 11694 29592 14962
rect 29656 14278 29684 15943
rect 29748 14550 29776 18022
rect 30024 17814 30052 18799
rect 30116 18193 30144 18838
rect 30102 18184 30158 18193
rect 30102 18119 30158 18128
rect 30012 17808 30064 17814
rect 30012 17750 30064 17756
rect 29920 17740 29972 17746
rect 29920 17682 29972 17688
rect 29932 17134 29960 17682
rect 30012 17604 30064 17610
rect 30012 17546 30064 17552
rect 30024 17513 30052 17546
rect 30010 17504 30066 17513
rect 30010 17439 30066 17448
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 30116 16794 30144 18119
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30116 16658 30144 16730
rect 30104 16652 30156 16658
rect 30104 16594 30156 16600
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 29828 16040 29880 16046
rect 30116 16017 30144 16050
rect 29828 15982 29880 15988
rect 30102 16008 30158 16017
rect 29840 15162 29868 15982
rect 30102 15943 30158 15952
rect 30208 15706 30236 19858
rect 30300 18970 30328 19858
rect 30392 19689 30420 19994
rect 30378 19680 30434 19689
rect 30378 19615 30434 19624
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30392 19174 30420 19314
rect 30484 19310 30512 21422
rect 30576 20398 30604 21678
rect 30656 21616 30708 21622
rect 30656 21558 30708 21564
rect 30564 20392 30616 20398
rect 30564 20334 30616 20340
rect 30564 20256 30616 20262
rect 30564 20198 30616 20204
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 30104 15428 30156 15434
rect 30104 15370 30156 15376
rect 29828 15156 29880 15162
rect 29880 15116 29960 15144
rect 29828 15098 29880 15104
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29656 12918 29684 14214
rect 29932 13462 29960 15116
rect 30116 14414 30144 15370
rect 30300 14958 30328 17682
rect 30392 17513 30420 19110
rect 30472 18624 30524 18630
rect 30472 18566 30524 18572
rect 30378 17504 30434 17513
rect 30378 17439 30434 17448
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30012 14408 30064 14414
rect 30012 14350 30064 14356
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30024 14074 30052 14350
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 29920 13456 29972 13462
rect 29920 13398 29972 13404
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29644 12912 29696 12918
rect 29644 12854 29696 12860
rect 29656 11801 29684 12854
rect 29642 11792 29698 11801
rect 29642 11727 29698 11736
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29656 11150 29684 11630
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29552 10600 29604 10606
rect 29656 10588 29684 11086
rect 29840 10606 29868 13330
rect 29932 12170 29960 13398
rect 30024 12850 30052 14010
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 30024 12306 30052 12786
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 30116 12209 30144 14350
rect 30208 13326 30236 14758
rect 30300 13818 30328 14894
rect 30392 14822 30420 14894
rect 30380 14816 30432 14822
rect 30378 14784 30380 14793
rect 30432 14784 30434 14793
rect 30378 14719 30434 14728
rect 30380 14612 30432 14618
rect 30380 14554 30432 14560
rect 30392 14278 30420 14554
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30300 13790 30420 13818
rect 30392 13462 30420 13790
rect 30380 13456 30432 13462
rect 30380 13398 30432 13404
rect 30484 13394 30512 18566
rect 30576 18222 30604 20198
rect 30668 18970 30696 21558
rect 30748 21344 30800 21350
rect 30748 21286 30800 21292
rect 30656 18964 30708 18970
rect 30656 18906 30708 18912
rect 30656 18828 30708 18834
rect 30656 18770 30708 18776
rect 30668 18630 30696 18770
rect 30656 18624 30708 18630
rect 30656 18566 30708 18572
rect 30564 18216 30616 18222
rect 30564 18158 30616 18164
rect 30760 18086 30788 21286
rect 30852 20602 30880 21966
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 30944 20874 30972 21490
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 31036 20534 31064 22120
rect 31208 21616 31260 21622
rect 31206 21584 31208 21593
rect 31260 21584 31262 21593
rect 31206 21519 31262 21528
rect 31116 21412 31168 21418
rect 31116 21354 31168 21360
rect 31128 21049 31156 21354
rect 31114 21040 31170 21049
rect 31114 20975 31170 20984
rect 31312 20806 31340 23190
rect 31392 23112 31444 23118
rect 31392 23054 31444 23060
rect 31404 22710 31432 23054
rect 31392 22704 31444 22710
rect 31392 22646 31444 22652
rect 31404 22094 31432 22646
rect 31482 22536 31538 22545
rect 31482 22471 31538 22480
rect 31496 22438 31524 22471
rect 31484 22432 31536 22438
rect 31484 22374 31536 22380
rect 31484 22094 31536 22098
rect 31404 22092 31536 22094
rect 31404 22066 31484 22092
rect 31484 22034 31536 22040
rect 31496 22003 31524 22034
rect 31392 21956 31444 21962
rect 31392 21898 31444 21904
rect 31404 21690 31432 21898
rect 31392 21684 31444 21690
rect 31392 21626 31444 21632
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31024 20528 31076 20534
rect 31024 20470 31076 20476
rect 31116 20392 31168 20398
rect 31116 20334 31168 20340
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30748 17604 30800 17610
rect 30748 17546 30800 17552
rect 30760 17270 30788 17546
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 30562 16416 30618 16425
rect 30562 16351 30618 16360
rect 30576 14482 30604 16351
rect 30668 16250 30696 17206
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 30656 16244 30708 16250
rect 30656 16186 30708 16192
rect 30760 15910 30788 17070
rect 30852 16114 30880 20198
rect 30930 19408 30986 19417
rect 30930 19343 30986 19352
rect 30944 18902 30972 19343
rect 31024 19236 31076 19242
rect 31024 19178 31076 19184
rect 30932 18896 30984 18902
rect 30932 18838 30984 18844
rect 30944 18737 30972 18838
rect 30930 18728 30986 18737
rect 30930 18663 30986 18672
rect 30932 18624 30984 18630
rect 30930 18592 30932 18601
rect 30984 18592 30986 18601
rect 30930 18527 30986 18536
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 30944 17338 30972 18158
rect 31036 18154 31064 19178
rect 31024 18148 31076 18154
rect 31024 18090 31076 18096
rect 31128 17746 31156 20334
rect 31220 18426 31248 20742
rect 31312 20534 31340 20742
rect 31484 20596 31536 20602
rect 31484 20538 31536 20544
rect 31300 20528 31352 20534
rect 31300 20470 31352 20476
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31300 19712 31352 19718
rect 31300 19654 31352 19660
rect 31312 18850 31340 19654
rect 31404 19514 31432 20198
rect 31392 19508 31444 19514
rect 31392 19450 31444 19456
rect 31496 19446 31524 20538
rect 31588 19854 31616 24278
rect 31850 24239 31906 24248
rect 32508 24206 32536 24550
rect 32876 24206 32904 24754
rect 33152 24614 33180 26200
rect 33796 24721 33824 26200
rect 33968 24744 34020 24750
rect 33782 24712 33838 24721
rect 33968 24686 34020 24692
rect 33782 24647 33838 24656
rect 33140 24608 33192 24614
rect 33140 24550 33192 24556
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 33048 24404 33100 24410
rect 33048 24346 33100 24352
rect 32496 24200 32548 24206
rect 32496 24142 32548 24148
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 31852 24064 31904 24070
rect 31852 24006 31904 24012
rect 32036 24064 32088 24070
rect 32036 24006 32088 24012
rect 32956 24064 33008 24070
rect 32956 24006 33008 24012
rect 31864 23662 31892 24006
rect 31760 23656 31812 23662
rect 31666 23624 31722 23633
rect 31760 23598 31812 23604
rect 31852 23656 31904 23662
rect 31852 23598 31904 23604
rect 31666 23559 31722 23568
rect 31680 22642 31708 23559
rect 31772 23186 31800 23598
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 31760 23044 31812 23050
rect 31864 23032 31892 23598
rect 32048 23594 32076 24006
rect 32588 23792 32640 23798
rect 32968 23769 32996 24006
rect 33060 23798 33088 24346
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33600 24064 33652 24070
rect 33600 24006 33652 24012
rect 33612 23905 33640 24006
rect 33598 23896 33654 23905
rect 33598 23831 33654 23840
rect 33048 23792 33100 23798
rect 32588 23734 32640 23740
rect 32954 23760 33010 23769
rect 32036 23588 32088 23594
rect 32036 23530 32088 23536
rect 31812 23004 31892 23032
rect 31760 22986 31812 22992
rect 31668 22636 31720 22642
rect 31668 22578 31720 22584
rect 31772 21690 31800 22986
rect 32128 22228 32180 22234
rect 32128 22170 32180 22176
rect 32140 22137 32168 22170
rect 32126 22128 32182 22137
rect 32126 22063 32182 22072
rect 31944 21888 31996 21894
rect 31944 21830 31996 21836
rect 32036 21888 32088 21894
rect 32036 21830 32088 21836
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31956 21554 31984 21830
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 31666 21040 31722 21049
rect 31666 20975 31722 20984
rect 31576 19848 31628 19854
rect 31576 19790 31628 19796
rect 31484 19440 31536 19446
rect 31484 19382 31536 19388
rect 31482 19136 31538 19145
rect 31482 19071 31538 19080
rect 31312 18822 31432 18850
rect 31404 18630 31432 18822
rect 31392 18624 31444 18630
rect 31392 18566 31444 18572
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31116 17740 31168 17746
rect 31116 17682 31168 17688
rect 31022 17368 31078 17377
rect 30932 17332 30984 17338
rect 31022 17303 31078 17312
rect 30932 17274 30984 17280
rect 31036 16726 31064 17303
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 31312 16726 31340 16934
rect 31024 16720 31076 16726
rect 31024 16662 31076 16668
rect 31300 16720 31352 16726
rect 31300 16662 31352 16668
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 31036 16114 31064 16526
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 31024 16108 31076 16114
rect 31024 16050 31076 16056
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30760 15434 30788 15846
rect 31116 15564 31168 15570
rect 31116 15506 31168 15512
rect 30656 15428 30708 15434
rect 30656 15370 30708 15376
rect 30748 15428 30800 15434
rect 30748 15370 30800 15376
rect 30668 15201 30696 15370
rect 30654 15192 30710 15201
rect 30654 15127 30656 15136
rect 30708 15127 30710 15136
rect 30656 15098 30708 15104
rect 30760 14482 30788 15370
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30852 14414 30880 15302
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 31128 14074 31156 15506
rect 31312 15162 31340 16390
rect 31404 16046 31432 18566
rect 31496 17882 31524 19071
rect 31588 18714 31616 19790
rect 31680 19514 31708 20975
rect 32048 20942 32076 21830
rect 32036 20936 32088 20942
rect 31758 20904 31814 20913
rect 32036 20878 32088 20884
rect 31758 20839 31760 20848
rect 31812 20839 31814 20848
rect 31760 20810 31812 20816
rect 32140 20534 32168 22063
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32416 21690 32444 21966
rect 32600 21894 32628 23734
rect 32680 23724 32732 23730
rect 33048 23734 33100 23740
rect 32954 23695 33010 23704
rect 32680 23666 32732 23672
rect 32692 21894 32720 23666
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33888 23322 33916 24142
rect 33232 23316 33284 23322
rect 33232 23258 33284 23264
rect 33876 23316 33928 23322
rect 33876 23258 33928 23264
rect 33244 23225 33272 23258
rect 33980 23254 34008 24686
rect 34244 24268 34296 24274
rect 34244 24210 34296 24216
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 34072 23254 34100 23666
rect 34256 23322 34284 24210
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 33968 23248 34020 23254
rect 33230 23216 33286 23225
rect 33968 23190 34020 23196
rect 34060 23248 34112 23254
rect 34060 23190 34112 23196
rect 33230 23151 33286 23160
rect 33784 22976 33836 22982
rect 33784 22918 33836 22924
rect 33600 22704 33652 22710
rect 33600 22646 33652 22652
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33428 22409 33456 22578
rect 33414 22400 33470 22409
rect 32950 22332 33258 22341
rect 33414 22335 33470 22344
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33612 22234 33640 22646
rect 33692 22500 33744 22506
rect 33692 22442 33744 22448
rect 33600 22228 33652 22234
rect 33600 22170 33652 22176
rect 33704 22094 33732 22442
rect 33612 22066 33732 22094
rect 32772 21956 32824 21962
rect 32772 21898 32824 21904
rect 32588 21888 32640 21894
rect 32588 21830 32640 21836
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 32128 20528 32180 20534
rect 32128 20470 32180 20476
rect 32324 20398 32352 20946
rect 32416 20874 32444 21626
rect 32496 20936 32548 20942
rect 32496 20878 32548 20884
rect 32586 20904 32642 20913
rect 32404 20868 32456 20874
rect 32404 20810 32456 20816
rect 32416 20534 32444 20810
rect 32508 20602 32536 20878
rect 32586 20839 32642 20848
rect 32496 20596 32548 20602
rect 32496 20538 32548 20544
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32312 20392 32364 20398
rect 31942 20360 31998 20369
rect 32312 20334 32364 20340
rect 31942 20295 31944 20304
rect 31996 20295 31998 20304
rect 31944 20266 31996 20272
rect 31956 19786 31984 20266
rect 31944 19780 31996 19786
rect 31944 19722 31996 19728
rect 32128 19712 32180 19718
rect 32128 19654 32180 19660
rect 31668 19508 31720 19514
rect 31668 19450 31720 19456
rect 31588 18686 31800 18714
rect 31668 18624 31720 18630
rect 31668 18566 31720 18572
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31484 17740 31536 17746
rect 31484 17682 31536 17688
rect 31392 16040 31444 16046
rect 31392 15982 31444 15988
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31116 14068 31168 14074
rect 31116 14010 31168 14016
rect 31128 13938 31156 14010
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 30840 13728 30892 13734
rect 30840 13670 30892 13676
rect 30472 13388 30524 13394
rect 30472 13330 30524 13336
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30562 13288 30618 13297
rect 30562 13223 30618 13232
rect 30196 12912 30248 12918
rect 30196 12854 30248 12860
rect 30102 12200 30158 12209
rect 29920 12164 29972 12170
rect 30102 12135 30158 12144
rect 29920 12106 29972 12112
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 29604 10560 29684 10588
rect 29828 10600 29880 10606
rect 29552 10542 29604 10548
rect 29828 10542 29880 10548
rect 29564 10130 29592 10542
rect 29840 10266 29868 10542
rect 29828 10260 29880 10266
rect 29828 10202 29880 10208
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 29564 9518 29592 10066
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29460 9444 29512 9450
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29196 8430 29224 9438
rect 29460 9386 29512 9392
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 26148 4752 26200 4758
rect 26148 4694 26200 4700
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25884 4214 25912 4422
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 24860 4072 24912 4078
rect 24858 4040 24860 4049
rect 25780 4072 25832 4078
rect 24912 4040 24914 4049
rect 25780 4014 25832 4020
rect 24858 3975 24914 3984
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24124 3528 24176 3534
rect 25792 3505 25820 4014
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 24124 3470 24176 3476
rect 25778 3496 25834 3505
rect 24044 3126 24072 3470
rect 25778 3431 25834 3440
rect 24584 3188 24636 3194
rect 24584 3130 24636 3136
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 24044 2650 24072 3062
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 22468 2576 22520 2582
rect 22468 2518 22520 2524
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22296 800 22324 2450
rect 24412 800 24440 2450
rect 24596 2446 24624 3130
rect 25976 2990 26004 3674
rect 26160 3058 26188 4694
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26344 3126 26372 3334
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26344 2650 26372 3062
rect 27540 2922 27568 3878
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 26528 800 26556 2450
rect 27172 2446 27200 2790
rect 27632 2650 27660 4082
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28828 3058 28856 8366
rect 29932 7954 29960 10610
rect 30116 9926 30144 12135
rect 30208 10810 30236 12854
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 30484 11286 30512 11494
rect 30472 11280 30524 11286
rect 30472 11222 30524 11228
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 30116 9518 30144 9590
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 30104 9512 30156 9518
rect 30104 9454 30156 9460
rect 30024 9110 30052 9454
rect 30484 9382 30512 10542
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30012 9104 30064 9110
rect 30012 9046 30064 9052
rect 30576 8090 30604 13223
rect 30852 11694 30880 13670
rect 31404 13172 31432 15846
rect 31496 15570 31524 17682
rect 31576 17332 31628 17338
rect 31576 17274 31628 17280
rect 31484 15564 31536 15570
rect 31484 15506 31536 15512
rect 31484 14884 31536 14890
rect 31484 14826 31536 14832
rect 31496 14346 31524 14826
rect 31484 14340 31536 14346
rect 31484 14282 31536 14288
rect 31588 13394 31616 17274
rect 31680 16454 31708 18566
rect 31772 17678 31800 18686
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 32036 18624 32088 18630
rect 32036 18566 32088 18572
rect 31956 18465 31984 18566
rect 31942 18456 31998 18465
rect 31942 18391 31998 18400
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31944 17536 31996 17542
rect 31944 17478 31996 17484
rect 31850 17368 31906 17377
rect 31850 17303 31906 17312
rect 31864 16998 31892 17303
rect 31760 16992 31812 16998
rect 31760 16934 31812 16940
rect 31852 16992 31904 16998
rect 31852 16934 31904 16940
rect 31668 16448 31720 16454
rect 31668 16390 31720 16396
rect 31772 16250 31800 16934
rect 31852 16584 31904 16590
rect 31852 16526 31904 16532
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 31668 16176 31720 16182
rect 31668 16118 31720 16124
rect 31680 13433 31708 16118
rect 31864 15910 31892 16526
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31852 15904 31904 15910
rect 31852 15846 31904 15852
rect 31772 15484 31800 15846
rect 31852 15496 31904 15502
rect 31772 15456 31852 15484
rect 31852 15438 31904 15444
rect 31760 15020 31812 15026
rect 31760 14962 31812 14968
rect 31666 13424 31722 13433
rect 31576 13388 31628 13394
rect 31666 13359 31722 13368
rect 31576 13330 31628 13336
rect 31668 13184 31720 13190
rect 31404 13144 31524 13172
rect 31496 12434 31524 13144
rect 31668 13126 31720 13132
rect 31496 12406 31616 12434
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31404 11830 31432 12038
rect 31588 11830 31616 12406
rect 31392 11824 31444 11830
rect 31392 11766 31444 11772
rect 31576 11824 31628 11830
rect 31576 11766 31628 11772
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 30840 11688 30892 11694
rect 30840 11630 30892 11636
rect 30748 11008 30800 11014
rect 30748 10950 30800 10956
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 30668 10130 30696 10610
rect 30656 10124 30708 10130
rect 30656 10066 30708 10072
rect 30656 9716 30708 9722
rect 30656 9658 30708 9664
rect 30668 8974 30696 9658
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30668 8838 30696 8910
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 30668 8566 30696 8774
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 30576 7886 30604 8026
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30484 7342 30512 7754
rect 30668 7750 30696 8502
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30472 7336 30524 7342
rect 30472 7278 30524 7284
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 29012 2650 29040 3470
rect 29644 3392 29696 3398
rect 29644 3334 29696 3340
rect 29656 3126 29684 3334
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 29656 2990 29684 3062
rect 30668 2990 30696 7686
rect 30760 6322 30788 10950
rect 31128 10810 31156 11698
rect 31576 11620 31628 11626
rect 31576 11562 31628 11568
rect 31392 11552 31444 11558
rect 31588 11506 31616 11562
rect 31444 11500 31616 11506
rect 31392 11494 31616 11500
rect 31404 11478 31616 11494
rect 31484 11212 31536 11218
rect 31484 11154 31536 11160
rect 31390 11112 31446 11121
rect 31496 11082 31524 11154
rect 31390 11047 31392 11056
rect 31444 11047 31446 11056
rect 31484 11076 31536 11082
rect 31392 11018 31444 11024
rect 31484 11018 31536 11024
rect 30840 10804 30892 10810
rect 30840 10746 30892 10752
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 30852 10606 30880 10746
rect 30840 10600 30892 10606
rect 30840 10542 30892 10548
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30852 10130 30880 10406
rect 31404 10266 31432 11018
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30840 9988 30892 9994
rect 30840 9930 30892 9936
rect 30852 9722 30880 9930
rect 31496 9722 31524 11018
rect 30840 9716 30892 9722
rect 30840 9658 30892 9664
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 31680 9654 31708 13126
rect 31772 11898 31800 14962
rect 31864 14006 31892 15438
rect 31852 14000 31904 14006
rect 31852 13942 31904 13948
rect 31864 13190 31892 13942
rect 31852 13184 31904 13190
rect 31852 13126 31904 13132
rect 31864 12850 31892 13126
rect 31852 12844 31904 12850
rect 31852 12786 31904 12792
rect 31864 12442 31892 12786
rect 31852 12436 31904 12442
rect 31852 12378 31904 12384
rect 31864 12170 31892 12378
rect 31852 12164 31904 12170
rect 31852 12106 31904 12112
rect 31864 11898 31892 12106
rect 31956 11898 31984 17478
rect 32048 16182 32076 18566
rect 32140 18358 32168 19654
rect 32508 19446 32536 20402
rect 32496 19440 32548 19446
rect 32496 19382 32548 19388
rect 32600 19378 32628 20839
rect 32784 20058 32812 21898
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33428 21690 33456 21830
rect 33416 21684 33468 21690
rect 33416 21626 33468 21632
rect 33506 21584 33562 21593
rect 33416 21548 33468 21554
rect 33506 21519 33508 21528
rect 33416 21490 33468 21496
rect 33560 21519 33562 21528
rect 33508 21490 33560 21496
rect 33324 21480 33376 21486
rect 33324 21422 33376 21428
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32864 21004 32916 21010
rect 32864 20946 32916 20952
rect 32772 20052 32824 20058
rect 32772 19994 32824 20000
rect 32876 19938 32904 20946
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32784 19910 32904 19938
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 32496 19304 32548 19310
rect 32496 19246 32548 19252
rect 32312 18420 32364 18426
rect 32312 18362 32364 18368
rect 32128 18352 32180 18358
rect 32128 18294 32180 18300
rect 32324 17542 32352 18362
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32312 17536 32364 17542
rect 32312 17478 32364 17484
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 32128 17060 32180 17066
rect 32128 17002 32180 17008
rect 32036 16176 32088 16182
rect 32036 16118 32088 16124
rect 32036 15156 32088 15162
rect 32036 15098 32088 15104
rect 32048 14346 32076 15098
rect 32036 14340 32088 14346
rect 32036 14282 32088 14288
rect 32140 12850 32168 17002
rect 32232 16658 32260 17138
rect 32324 17066 32352 17478
rect 32416 17377 32444 18158
rect 32402 17368 32458 17377
rect 32402 17303 32458 17312
rect 32312 17060 32364 17066
rect 32312 17002 32364 17008
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 32220 16516 32272 16522
rect 32220 16458 32272 16464
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 31760 11892 31812 11898
rect 31760 11834 31812 11840
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 31944 11892 31996 11898
rect 31944 11834 31996 11840
rect 31944 11688 31996 11694
rect 31944 11630 31996 11636
rect 31956 10470 31984 11630
rect 32140 11218 32168 12174
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 31760 10464 31812 10470
rect 31760 10406 31812 10412
rect 31944 10464 31996 10470
rect 31944 10406 31996 10412
rect 31668 9648 31720 9654
rect 31668 9590 31720 9596
rect 31772 9586 31800 10406
rect 31956 10146 31984 10406
rect 31956 10118 32076 10146
rect 32140 10130 32168 11154
rect 32232 10198 32260 16458
rect 32324 15366 32352 17002
rect 32416 16522 32444 17303
rect 32404 16516 32456 16522
rect 32404 16458 32456 16464
rect 32416 16425 32444 16458
rect 32402 16416 32458 16425
rect 32402 16351 32458 16360
rect 32508 16046 32536 19246
rect 32784 18834 32812 19910
rect 32864 19508 32916 19514
rect 32864 19450 32916 19456
rect 32772 18828 32824 18834
rect 32772 18770 32824 18776
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 32496 16040 32548 16046
rect 32496 15982 32548 15988
rect 32600 16028 32628 17070
rect 32772 16040 32824 16046
rect 32600 16000 32772 16028
rect 32404 15564 32456 15570
rect 32404 15506 32456 15512
rect 32312 15360 32364 15366
rect 32312 15302 32364 15308
rect 32312 15088 32364 15094
rect 32312 15030 32364 15036
rect 32324 13870 32352 15030
rect 32416 14482 32444 15506
rect 32404 14476 32456 14482
rect 32404 14418 32456 14424
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32416 13172 32444 14418
rect 32324 13144 32444 13172
rect 32324 11121 32352 13144
rect 32404 12980 32456 12986
rect 32404 12922 32456 12928
rect 32416 12306 32444 12922
rect 32404 12300 32456 12306
rect 32404 12242 32456 12248
rect 32310 11112 32366 11121
rect 32310 11047 32366 11056
rect 32312 10804 32364 10810
rect 32312 10746 32364 10752
rect 32324 10606 32352 10746
rect 32416 10606 32444 12242
rect 32508 10810 32536 15982
rect 32600 15638 32628 16000
rect 32772 15982 32824 15988
rect 32680 15904 32732 15910
rect 32680 15846 32732 15852
rect 32588 15632 32640 15638
rect 32588 15574 32640 15580
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 32600 12986 32628 14418
rect 32588 12980 32640 12986
rect 32588 12922 32640 12928
rect 32692 12434 32720 15846
rect 32876 14414 32904 19450
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32954 18864 33010 18873
rect 32954 18799 32956 18808
rect 33008 18799 33010 18808
rect 33048 18828 33100 18834
rect 32956 18770 33008 18776
rect 33048 18770 33100 18776
rect 33060 18578 33088 18770
rect 32968 18550 33088 18578
rect 32968 18426 32996 18550
rect 32956 18420 33008 18426
rect 32956 18362 33008 18368
rect 33336 18290 33364 21422
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 33232 17740 33284 17746
rect 33428 17728 33456 21490
rect 33612 19718 33640 22066
rect 33692 20528 33744 20534
rect 33692 20470 33744 20476
rect 33600 19712 33652 19718
rect 33600 19654 33652 19660
rect 33600 18896 33652 18902
rect 33598 18864 33600 18873
rect 33652 18864 33654 18873
rect 33598 18799 33654 18808
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33284 17700 33456 17728
rect 33232 17682 33284 17688
rect 33416 17536 33468 17542
rect 33416 17478 33468 17484
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 33336 14550 33364 16050
rect 33428 15978 33456 17478
rect 33612 17338 33640 18158
rect 33704 18086 33732 20470
rect 33796 19854 33824 22918
rect 33980 22574 34008 23190
rect 34072 22982 34100 23190
rect 34336 23180 34388 23186
rect 34336 23122 34388 23128
rect 34060 22976 34112 22982
rect 34060 22918 34112 22924
rect 34244 22704 34296 22710
rect 34348 22658 34376 23122
rect 34296 22652 34376 22658
rect 34244 22646 34376 22652
rect 34256 22630 34376 22646
rect 33968 22568 34020 22574
rect 33968 22510 34020 22516
rect 34244 22024 34296 22030
rect 34244 21966 34296 21972
rect 33876 21956 33928 21962
rect 33876 21898 33928 21904
rect 33784 19848 33836 19854
rect 33784 19790 33836 19796
rect 33888 19666 33916 21898
rect 33968 21344 34020 21350
rect 33968 21286 34020 21292
rect 33796 19638 33916 19666
rect 33692 18080 33744 18086
rect 33692 18022 33744 18028
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 33416 15972 33468 15978
rect 33416 15914 33468 15920
rect 33692 15904 33744 15910
rect 33692 15846 33744 15852
rect 33508 15360 33560 15366
rect 33508 15302 33560 15308
rect 33520 14550 33548 15302
rect 33324 14544 33376 14550
rect 33324 14486 33376 14492
rect 33508 14544 33560 14550
rect 33508 14486 33560 14492
rect 32864 14408 32916 14414
rect 33520 14396 33548 14486
rect 33704 14414 33732 15846
rect 33796 15162 33824 19638
rect 33980 19446 34008 21286
rect 34256 21078 34284 21966
rect 34348 21894 34376 22630
rect 34440 22001 34468 26200
rect 34888 24812 34940 24818
rect 34888 24754 34940 24760
rect 34612 24404 34664 24410
rect 34612 24346 34664 24352
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 34532 23050 34560 23598
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34520 22704 34572 22710
rect 34520 22646 34572 22652
rect 34532 22098 34560 22646
rect 34520 22092 34572 22098
rect 34520 22034 34572 22040
rect 34426 21992 34482 22001
rect 34426 21927 34482 21936
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 34244 21072 34296 21078
rect 34244 21014 34296 21020
rect 34348 21010 34376 21830
rect 34428 21412 34480 21418
rect 34428 21354 34480 21360
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 34440 20806 34468 21354
rect 34532 20942 34560 22034
rect 34624 21690 34652 24346
rect 34794 23760 34850 23769
rect 34794 23695 34850 23704
rect 34808 22681 34836 23695
rect 34794 22672 34850 22681
rect 34794 22607 34850 22616
rect 34704 22228 34756 22234
rect 34704 22170 34756 22176
rect 34716 21690 34744 22170
rect 34808 21690 34836 22607
rect 34900 22137 34928 24754
rect 34980 24676 35032 24682
rect 34980 24618 35032 24624
rect 34992 24070 35020 24618
rect 34980 24064 35032 24070
rect 34980 24006 35032 24012
rect 35084 23497 35112 26200
rect 35164 24744 35216 24750
rect 35164 24686 35216 24692
rect 35176 24274 35204 24686
rect 35164 24268 35216 24274
rect 35164 24210 35216 24216
rect 35532 24132 35584 24138
rect 35532 24074 35584 24080
rect 35440 24064 35492 24070
rect 35438 24032 35440 24041
rect 35492 24032 35494 24041
rect 35438 23967 35494 23976
rect 35452 23730 35480 23967
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 35348 23656 35400 23662
rect 35348 23598 35400 23604
rect 35070 23488 35126 23497
rect 35070 23423 35126 23432
rect 35360 23186 35388 23598
rect 35440 23588 35492 23594
rect 35440 23530 35492 23536
rect 35348 23180 35400 23186
rect 35348 23122 35400 23128
rect 35162 23080 35218 23089
rect 35162 23015 35218 23024
rect 35176 22794 35204 23015
rect 35176 22778 35296 22794
rect 35452 22778 35480 23530
rect 35544 22778 35572 24074
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35636 23798 35664 24006
rect 35624 23792 35676 23798
rect 35624 23734 35676 23740
rect 35624 23656 35676 23662
rect 35624 23598 35676 23604
rect 35176 22772 35308 22778
rect 35176 22766 35256 22772
rect 35072 22432 35124 22438
rect 35072 22374 35124 22380
rect 34886 22128 34942 22137
rect 35084 22098 35112 22374
rect 34886 22063 34942 22072
rect 35072 22092 35124 22098
rect 35072 22034 35124 22040
rect 34612 21684 34664 21690
rect 34612 21626 34664 21632
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 34796 21684 34848 21690
rect 34796 21626 34848 21632
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 35072 20936 35124 20942
rect 35072 20878 35124 20884
rect 34428 20800 34480 20806
rect 34428 20742 34480 20748
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34072 20398 34100 20538
rect 34440 20534 34468 20742
rect 35084 20641 35112 20878
rect 35070 20632 35126 20641
rect 35070 20567 35126 20576
rect 34428 20528 34480 20534
rect 34428 20470 34480 20476
rect 34888 20460 34940 20466
rect 34888 20402 34940 20408
rect 35072 20460 35124 20466
rect 35072 20402 35124 20408
rect 34060 20392 34112 20398
rect 34060 20334 34112 20340
rect 33968 19440 34020 19446
rect 33968 19382 34020 19388
rect 33968 19168 34020 19174
rect 33968 19110 34020 19116
rect 33980 17814 34008 19110
rect 34072 18834 34100 20334
rect 34518 20224 34574 20233
rect 34518 20159 34574 20168
rect 34336 20052 34388 20058
rect 34336 19994 34388 20000
rect 34244 19780 34296 19786
rect 34244 19722 34296 19728
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 34060 18828 34112 18834
rect 34060 18770 34112 18776
rect 34164 18630 34192 19314
rect 34256 19242 34284 19722
rect 34348 19718 34376 19994
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 34244 19236 34296 19242
rect 34244 19178 34296 19184
rect 34244 18896 34296 18902
rect 34242 18864 34244 18873
rect 34296 18864 34298 18873
rect 34242 18799 34298 18808
rect 34152 18624 34204 18630
rect 34152 18566 34204 18572
rect 33968 17808 34020 17814
rect 33968 17750 34020 17756
rect 34058 17368 34114 17377
rect 34058 17303 34060 17312
rect 34112 17303 34114 17312
rect 34060 17274 34112 17280
rect 33876 17264 33928 17270
rect 33876 17206 33928 17212
rect 33888 16522 33916 17206
rect 33876 16516 33928 16522
rect 33876 16458 33928 16464
rect 33968 16448 34020 16454
rect 33968 16390 34020 16396
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33888 15162 33916 15302
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 33876 15156 33928 15162
rect 33876 15098 33928 15104
rect 33980 15026 34008 16390
rect 34072 15502 34100 16390
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 33968 15020 34020 15026
rect 33968 14962 34020 14968
rect 33784 14952 33836 14958
rect 33784 14894 33836 14900
rect 33796 14618 33824 14894
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 32864 14350 32916 14356
rect 33428 14368 33548 14396
rect 33692 14408 33744 14414
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 32600 12406 32720 12434
rect 32496 10804 32548 10810
rect 32496 10746 32548 10752
rect 32312 10600 32364 10606
rect 32312 10542 32364 10548
rect 32404 10600 32456 10606
rect 32404 10542 32456 10548
rect 32600 10266 32628 12406
rect 32784 11898 32812 14214
rect 33324 14000 33376 14006
rect 33324 13942 33376 13948
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 33336 13190 33364 13942
rect 33324 13184 33376 13190
rect 33324 13126 33376 13132
rect 33336 12646 33364 13126
rect 33324 12640 33376 12646
rect 33324 12582 33376 12588
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32772 11892 32824 11898
rect 32772 11834 32824 11840
rect 32680 11688 32732 11694
rect 32680 11630 32732 11636
rect 32692 11286 32720 11630
rect 32864 11552 32916 11558
rect 32864 11494 32916 11500
rect 32680 11280 32732 11286
rect 32680 11222 32732 11228
rect 32876 11234 32904 11494
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 32956 11280 33008 11286
rect 32876 11228 32956 11234
rect 32876 11222 33008 11228
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 32220 10192 32272 10198
rect 32220 10134 32272 10140
rect 31852 9988 31904 9994
rect 31852 9930 31904 9936
rect 31944 9988 31996 9994
rect 31944 9930 31996 9936
rect 31116 9580 31168 9586
rect 31116 9522 31168 9528
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 31128 9382 31156 9522
rect 31864 9518 31892 9930
rect 31852 9512 31904 9518
rect 31852 9454 31904 9460
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 31128 8974 31156 9318
rect 31760 9036 31812 9042
rect 31760 8978 31812 8984
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31128 7546 31156 8570
rect 31772 8498 31800 8978
rect 31760 8492 31812 8498
rect 31760 8434 31812 8440
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31312 7342 31340 8366
rect 31864 8362 31892 9454
rect 31956 8838 31984 9930
rect 31944 8832 31996 8838
rect 31944 8774 31996 8780
rect 31944 8560 31996 8566
rect 31944 8502 31996 8508
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31404 7546 31432 7686
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31956 7478 31984 8502
rect 32048 8498 32076 10118
rect 32128 10124 32180 10130
rect 32128 10066 32180 10072
rect 32588 10124 32640 10130
rect 32588 10066 32640 10072
rect 32140 9654 32168 10066
rect 32128 9648 32180 9654
rect 32128 9590 32180 9596
rect 32140 9042 32168 9590
rect 32600 9450 32628 10066
rect 32588 9444 32640 9450
rect 32588 9386 32640 9392
rect 32128 9036 32180 9042
rect 32128 8978 32180 8984
rect 32140 8498 32168 8978
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32600 8566 32628 8910
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32036 8492 32088 8498
rect 32036 8434 32088 8440
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 32692 8430 32720 11222
rect 32876 11206 32996 11222
rect 33336 11150 33364 11290
rect 33232 11144 33284 11150
rect 33232 11086 33284 11092
rect 33324 11144 33376 11150
rect 33324 11086 33376 11092
rect 33244 10742 33272 11086
rect 33232 10736 33284 10742
rect 33232 10678 33284 10684
rect 32864 10464 32916 10470
rect 32864 10406 32916 10412
rect 32772 10056 32824 10062
rect 32772 9998 32824 10004
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32680 8424 32732 8430
rect 32680 8366 32732 8372
rect 32232 7954 32260 8366
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32784 7886 32812 9998
rect 32876 9160 32904 10406
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33232 9920 33284 9926
rect 33284 9868 33364 9874
rect 33232 9862 33364 9868
rect 33244 9846 33364 9862
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32876 9132 32996 9160
rect 32968 8430 32996 9132
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32772 7880 32824 7886
rect 32772 7822 32824 7828
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 31944 7472 31996 7478
rect 31944 7414 31996 7420
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 32600 7274 32628 7686
rect 33336 7410 33364 9846
rect 33324 7404 33376 7410
rect 33324 7346 33376 7352
rect 32588 7268 32640 7274
rect 32588 7210 32640 7216
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32772 4616 32824 4622
rect 32772 4558 32824 4564
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 32784 2582 32812 4558
rect 32864 4072 32916 4078
rect 32864 4014 32916 4020
rect 32876 2650 32904 4014
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 33336 3534 33364 5170
rect 33428 3670 33456 14368
rect 33692 14350 33744 14356
rect 33692 14272 33744 14278
rect 33692 14214 33744 14220
rect 33704 13462 33732 14214
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 33784 13524 33836 13530
rect 33784 13466 33836 13472
rect 33692 13456 33744 13462
rect 33692 13398 33744 13404
rect 33704 13190 33732 13398
rect 33692 13184 33744 13190
rect 33692 13126 33744 13132
rect 33704 12986 33732 13126
rect 33692 12980 33744 12986
rect 33692 12922 33744 12928
rect 33704 12434 33732 12922
rect 33612 12406 33732 12434
rect 33508 12232 33560 12238
rect 33508 12174 33560 12180
rect 33520 10742 33548 12174
rect 33508 10736 33560 10742
rect 33508 10678 33560 10684
rect 33520 9722 33548 10678
rect 33508 9716 33560 9722
rect 33508 9658 33560 9664
rect 33520 9178 33548 9658
rect 33508 9172 33560 9178
rect 33508 9114 33560 9120
rect 33612 9042 33640 12406
rect 33796 11744 33824 13466
rect 33876 13388 33928 13394
rect 33876 13330 33928 13336
rect 33888 12782 33916 13330
rect 34072 13326 34100 13806
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 33968 13252 34020 13258
rect 33968 13194 34020 13200
rect 33876 12776 33928 12782
rect 33876 12718 33928 12724
rect 33980 12594 34008 13194
rect 34072 12986 34100 13262
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 33888 12566 34008 12594
rect 33888 12442 33916 12566
rect 33876 12436 33928 12442
rect 34164 12434 34192 18566
rect 34244 17808 34296 17814
rect 34244 17750 34296 17756
rect 34256 15094 34284 17750
rect 34348 16454 34376 19654
rect 34532 19514 34560 20159
rect 34900 20058 34928 20402
rect 34980 20392 35032 20398
rect 34980 20334 35032 20340
rect 34888 20052 34940 20058
rect 34888 19994 34940 20000
rect 34704 19984 34756 19990
rect 34704 19926 34756 19932
rect 34520 19508 34572 19514
rect 34520 19450 34572 19456
rect 34532 18902 34560 19450
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 34520 18216 34572 18222
rect 34520 18158 34572 18164
rect 34532 17746 34560 18158
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34532 16794 34560 17682
rect 34520 16788 34572 16794
rect 34520 16730 34572 16736
rect 34336 16448 34388 16454
rect 34336 16390 34388 16396
rect 34336 15972 34388 15978
rect 34336 15914 34388 15920
rect 34244 15088 34296 15094
rect 34244 15030 34296 15036
rect 34244 14816 34296 14822
rect 34244 14758 34296 14764
rect 34256 14618 34284 14758
rect 34244 14612 34296 14618
rect 34244 14554 34296 14560
rect 34348 13190 34376 15914
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 34428 15632 34480 15638
rect 34428 15574 34480 15580
rect 34440 14074 34468 15574
rect 34624 15473 34652 15846
rect 34610 15464 34666 15473
rect 34610 15399 34666 15408
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 34716 13938 34744 19926
rect 34900 19514 34928 19994
rect 34888 19508 34940 19514
rect 34888 19450 34940 19456
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34808 16250 34836 17070
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 34808 15570 34836 16186
rect 34900 16153 34928 19450
rect 34992 19310 35020 20334
rect 35084 19922 35112 20402
rect 35072 19916 35124 19922
rect 35072 19858 35124 19864
rect 34980 19304 35032 19310
rect 34980 19246 35032 19252
rect 34992 19009 35020 19246
rect 35084 19174 35112 19858
rect 35176 19854 35204 22766
rect 35256 22714 35308 22720
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 35532 22772 35584 22778
rect 35532 22714 35584 22720
rect 35346 22400 35402 22409
rect 35346 22335 35402 22344
rect 35256 21888 35308 21894
rect 35256 21830 35308 21836
rect 35268 21690 35296 21830
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35268 20505 35296 21626
rect 35254 20496 35310 20505
rect 35254 20431 35310 20440
rect 35164 19848 35216 19854
rect 35164 19790 35216 19796
rect 35360 19718 35388 22335
rect 35452 22166 35480 22714
rect 35440 22160 35492 22166
rect 35440 22102 35492 22108
rect 35636 21434 35664 23598
rect 35728 22681 35756 26200
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 35992 23656 36044 23662
rect 36096 23633 36124 24006
rect 35992 23598 36044 23604
rect 36082 23624 36138 23633
rect 35714 22672 35770 22681
rect 35714 22607 35770 22616
rect 36004 21894 36032 23598
rect 36082 23559 36138 23568
rect 36268 23520 36320 23526
rect 36268 23462 36320 23468
rect 36280 22982 36308 23462
rect 36268 22976 36320 22982
rect 36268 22918 36320 22924
rect 36372 22778 36400 26200
rect 36910 24440 36966 24449
rect 36910 24375 36966 24384
rect 36452 24336 36504 24342
rect 36452 24278 36504 24284
rect 36464 23662 36492 24278
rect 36820 24132 36872 24138
rect 36820 24074 36872 24080
rect 36452 23656 36504 23662
rect 36452 23598 36504 23604
rect 36636 22976 36688 22982
rect 36636 22918 36688 22924
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 36360 22636 36412 22642
rect 36360 22578 36412 22584
rect 36268 22568 36320 22574
rect 36268 22510 36320 22516
rect 36280 21978 36308 22510
rect 36096 21950 36308 21978
rect 35992 21888 36044 21894
rect 35992 21830 36044 21836
rect 35990 21720 36046 21729
rect 35990 21655 36046 21664
rect 35452 21406 35664 21434
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 35072 19168 35124 19174
rect 35072 19110 35124 19116
rect 34978 19000 35034 19009
rect 34978 18935 35034 18944
rect 35254 19000 35310 19009
rect 35254 18935 35310 18944
rect 34980 18080 35032 18086
rect 34980 18022 35032 18028
rect 34992 17814 35020 18022
rect 34980 17808 35032 17814
rect 34980 17750 35032 17756
rect 34992 17270 35020 17750
rect 35072 17536 35124 17542
rect 35072 17478 35124 17484
rect 35084 17338 35112 17478
rect 35072 17332 35124 17338
rect 35072 17274 35124 17280
rect 34980 17264 35032 17270
rect 34980 17206 35032 17212
rect 34992 16726 35020 17206
rect 34980 16720 35032 16726
rect 34980 16662 35032 16668
rect 34992 16182 35020 16662
rect 34980 16176 35032 16182
rect 34886 16144 34942 16153
rect 34980 16118 35032 16124
rect 34886 16079 34942 16088
rect 34992 15706 35020 16118
rect 35164 15904 35216 15910
rect 35164 15846 35216 15852
rect 34980 15700 35032 15706
rect 34980 15642 35032 15648
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 34808 14482 34836 15506
rect 34992 15416 35020 15642
rect 35072 15428 35124 15434
rect 34992 15388 35072 15416
rect 35072 15370 35124 15376
rect 34888 15088 34940 15094
rect 34888 15030 34940 15036
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 34704 13932 34756 13938
rect 34704 13874 34756 13880
rect 34704 13796 34756 13802
rect 34704 13738 34756 13744
rect 34336 13184 34388 13190
rect 34336 13126 34388 13132
rect 34244 12640 34296 12646
rect 34244 12582 34296 12588
rect 33876 12378 33928 12384
rect 33980 12406 34192 12434
rect 33876 11756 33928 11762
rect 33796 11716 33876 11744
rect 33876 11698 33928 11704
rect 33980 11014 34008 12406
rect 34256 12374 34284 12582
rect 34244 12368 34296 12374
rect 34244 12310 34296 12316
rect 34348 12102 34376 13126
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34336 12096 34388 12102
rect 34336 12038 34388 12044
rect 33692 11008 33744 11014
rect 33692 10950 33744 10956
rect 33968 11008 34020 11014
rect 33968 10950 34020 10956
rect 33704 9489 33732 10950
rect 34244 9512 34296 9518
rect 33690 9480 33746 9489
rect 34244 9454 34296 9460
rect 33690 9415 33746 9424
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 33612 8362 33640 8978
rect 33704 8838 33732 9415
rect 34060 9036 34112 9042
rect 34060 8978 34112 8984
rect 34072 8906 34100 8978
rect 34256 8974 34284 9454
rect 34244 8968 34296 8974
rect 34244 8910 34296 8916
rect 34060 8900 34112 8906
rect 34060 8842 34112 8848
rect 34152 8900 34204 8906
rect 34152 8842 34204 8848
rect 33692 8832 33744 8838
rect 33692 8774 33744 8780
rect 34072 8634 34100 8842
rect 33876 8628 33928 8634
rect 33876 8570 33928 8576
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33888 8430 33916 8570
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 34164 8090 34192 8842
rect 34256 8634 34284 8910
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 34152 8084 34204 8090
rect 34152 8026 34204 8032
rect 33416 3664 33468 3670
rect 33416 3606 33468 3612
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 34348 2582 34376 12038
rect 34440 11694 34468 12786
rect 34520 12708 34572 12714
rect 34520 12650 34572 12656
rect 34428 11688 34480 11694
rect 34428 11630 34480 11636
rect 34440 11354 34468 11630
rect 34428 11348 34480 11354
rect 34428 11290 34480 11296
rect 34428 9716 34480 9722
rect 34428 9658 34480 9664
rect 34440 9625 34468 9658
rect 34426 9616 34482 9625
rect 34426 9551 34482 9560
rect 34532 8974 34560 12650
rect 34612 11552 34664 11558
rect 34612 11494 34664 11500
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34624 8838 34652 11494
rect 34716 10130 34744 13738
rect 34900 13410 34928 15030
rect 35176 14346 35204 15846
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 34808 13382 34928 13410
rect 34808 12782 34836 13382
rect 34888 13320 34940 13326
rect 34888 13262 34940 13268
rect 35162 13288 35218 13297
rect 34900 12918 34928 13262
rect 35162 13223 35164 13232
rect 35216 13223 35218 13232
rect 35164 13194 35216 13200
rect 35176 12986 35204 13194
rect 35164 12980 35216 12986
rect 35164 12922 35216 12928
rect 34888 12912 34940 12918
rect 34888 12854 34940 12860
rect 34796 12776 34848 12782
rect 34796 12718 34848 12724
rect 34808 12306 34836 12718
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 34704 10124 34756 10130
rect 34704 10066 34756 10072
rect 34704 9648 34756 9654
rect 34702 9616 34704 9625
rect 34756 9616 34758 9625
rect 34702 9551 34758 9560
rect 34612 8832 34664 8838
rect 34612 8774 34664 8780
rect 34716 8566 34744 9551
rect 34704 8560 34756 8566
rect 34704 8502 34756 8508
rect 34808 7954 34836 12242
rect 34900 12238 34928 12854
rect 35268 12594 35296 18935
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 35360 18426 35388 18702
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35452 17184 35480 21406
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35530 20632 35586 20641
rect 35530 20567 35586 20576
rect 35544 20330 35572 20567
rect 35532 20324 35584 20330
rect 35532 20266 35584 20272
rect 35532 18692 35584 18698
rect 35532 18634 35584 18640
rect 35544 18426 35572 18634
rect 35532 18420 35584 18426
rect 35532 18362 35584 18368
rect 35532 17536 35584 17542
rect 35530 17504 35532 17513
rect 35584 17504 35586 17513
rect 35530 17439 35586 17448
rect 35544 17270 35572 17439
rect 35532 17264 35584 17270
rect 35532 17206 35584 17212
rect 35360 17156 35480 17184
rect 35360 16998 35388 17156
rect 35440 17060 35492 17066
rect 35440 17002 35492 17008
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 35348 15360 35400 15366
rect 35452 15337 35480 17002
rect 35544 16590 35572 17206
rect 35636 17202 35664 21286
rect 35728 21146 35756 21286
rect 35716 21140 35768 21146
rect 35716 21082 35768 21088
rect 36004 20330 36032 21655
rect 35992 20324 36044 20330
rect 35992 20266 36044 20272
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35900 19712 35952 19718
rect 35900 19654 35952 19660
rect 35716 18148 35768 18154
rect 35716 18090 35768 18096
rect 35728 17746 35756 18090
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 35624 17196 35676 17202
rect 35624 17138 35676 17144
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 35714 16008 35770 16017
rect 35532 15972 35584 15978
rect 35714 15943 35770 15952
rect 35532 15914 35584 15920
rect 35348 15302 35400 15308
rect 35438 15328 35494 15337
rect 35360 14362 35388 15302
rect 35438 15263 35494 15272
rect 35360 14346 35480 14362
rect 35360 14340 35492 14346
rect 35360 14334 35440 14340
rect 35440 14282 35492 14288
rect 35348 14272 35400 14278
rect 35452 14249 35480 14282
rect 35348 14214 35400 14220
rect 35438 14240 35494 14249
rect 34992 12566 35296 12594
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 34900 11694 34928 12174
rect 34888 11688 34940 11694
rect 34888 11630 34940 11636
rect 34888 11212 34940 11218
rect 34888 11154 34940 11160
rect 34900 10062 34928 11154
rect 34992 10577 35020 12566
rect 35360 12434 35388 14214
rect 35438 14175 35494 14184
rect 35452 12646 35480 14175
rect 35544 13530 35572 15914
rect 35624 15700 35676 15706
rect 35624 15642 35676 15648
rect 35636 15162 35664 15642
rect 35624 15156 35676 15162
rect 35624 15098 35676 15104
rect 35728 14385 35756 15943
rect 35820 15094 35848 19654
rect 35912 18465 35940 19654
rect 35992 19304 36044 19310
rect 35992 19246 36044 19252
rect 35898 18456 35954 18465
rect 35898 18391 35954 18400
rect 36004 17728 36032 19246
rect 36096 18970 36124 21950
rect 36268 21888 36320 21894
rect 36268 21830 36320 21836
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36188 20602 36216 21422
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36280 19786 36308 21830
rect 36268 19780 36320 19786
rect 36268 19722 36320 19728
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 36084 18964 36136 18970
rect 36280 18952 36308 19314
rect 36084 18906 36136 18912
rect 36188 18924 36308 18952
rect 36188 18358 36216 18924
rect 36372 18850 36400 22578
rect 36648 22506 36676 22918
rect 36636 22500 36688 22506
rect 36636 22442 36688 22448
rect 36832 21894 36860 24074
rect 36924 23032 36952 24375
rect 36924 23004 37044 23032
rect 36912 22500 36964 22506
rect 36912 22442 36964 22448
rect 36820 21888 36872 21894
rect 36820 21830 36872 21836
rect 36820 21548 36872 21554
rect 36820 21490 36872 21496
rect 36452 21480 36504 21486
rect 36452 21422 36504 21428
rect 36464 20874 36492 21422
rect 36636 21140 36688 21146
rect 36636 21082 36688 21088
rect 36452 20868 36504 20874
rect 36452 20810 36504 20816
rect 36464 20602 36492 20810
rect 36648 20806 36676 21082
rect 36728 20868 36780 20874
rect 36728 20810 36780 20816
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36740 20641 36768 20810
rect 36726 20632 36782 20641
rect 36452 20596 36504 20602
rect 36726 20567 36782 20576
rect 36452 20538 36504 20544
rect 36740 20534 36768 20567
rect 36728 20528 36780 20534
rect 36728 20470 36780 20476
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 36280 18822 36400 18850
rect 36280 18630 36308 18822
rect 36268 18624 36320 18630
rect 36268 18566 36320 18572
rect 36176 18352 36228 18358
rect 36176 18294 36228 18300
rect 36268 18284 36320 18290
rect 36268 18226 36320 18232
rect 35912 17700 36032 17728
rect 35912 16522 35940 17700
rect 35992 17604 36044 17610
rect 35992 17546 36044 17552
rect 35900 16516 35952 16522
rect 35900 16458 35952 16464
rect 35912 15570 35940 16458
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 36004 15178 36032 17546
rect 36176 17128 36228 17134
rect 36176 17070 36228 17076
rect 36004 15162 36124 15178
rect 36004 15156 36136 15162
rect 36004 15150 36084 15156
rect 36084 15098 36136 15104
rect 35808 15088 35860 15094
rect 35808 15030 35860 15036
rect 35912 15014 36124 15042
rect 35912 14958 35940 15014
rect 36096 14958 36124 15014
rect 35900 14952 35952 14958
rect 35900 14894 35952 14900
rect 35992 14952 36044 14958
rect 35992 14894 36044 14900
rect 36084 14952 36136 14958
rect 36084 14894 36136 14900
rect 35714 14376 35770 14385
rect 35714 14311 35770 14320
rect 35808 14272 35860 14278
rect 35808 14214 35860 14220
rect 35900 14272 35952 14278
rect 35900 14214 35952 14220
rect 35820 14074 35848 14214
rect 35716 14068 35768 14074
rect 35716 14010 35768 14016
rect 35808 14068 35860 14074
rect 35808 14010 35860 14016
rect 35532 13524 35584 13530
rect 35532 13466 35584 13472
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 35176 12406 35388 12434
rect 35072 11620 35124 11626
rect 35072 11562 35124 11568
rect 35084 11354 35112 11562
rect 35072 11348 35124 11354
rect 35072 11290 35124 11296
rect 35176 11082 35204 12406
rect 35452 12170 35480 12582
rect 35440 12164 35492 12170
rect 35440 12106 35492 12112
rect 35452 11898 35480 12106
rect 35728 11914 35756 14010
rect 35912 13734 35940 14214
rect 36004 13954 36032 14894
rect 36188 14657 36216 17070
rect 36280 16046 36308 18226
rect 36360 17196 36412 17202
rect 36360 17138 36412 17144
rect 36372 16794 36400 17138
rect 36464 17066 36492 20402
rect 36634 20088 36690 20097
rect 36634 20023 36690 20032
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36556 19514 36584 19654
rect 36648 19553 36676 20023
rect 36728 19916 36780 19922
rect 36728 19858 36780 19864
rect 36634 19544 36690 19553
rect 36544 19508 36596 19514
rect 36634 19479 36690 19488
rect 36544 19450 36596 19456
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36544 18080 36596 18086
rect 36544 18022 36596 18028
rect 36556 17610 36584 18022
rect 36544 17604 36596 17610
rect 36544 17546 36596 17552
rect 36648 17542 36676 19110
rect 36740 18154 36768 19858
rect 36832 18426 36860 21490
rect 36924 21486 36952 22442
rect 37016 22094 37044 23004
rect 37108 22273 37136 26302
rect 37646 26302 37872 26330
rect 37646 26200 37702 26302
rect 37556 24676 37608 24682
rect 37556 24618 37608 24624
rect 37648 24676 37700 24682
rect 37648 24618 37700 24624
rect 37188 24268 37240 24274
rect 37188 24210 37240 24216
rect 37372 24268 37424 24274
rect 37372 24210 37424 24216
rect 37094 22264 37150 22273
rect 37094 22199 37150 22208
rect 37016 22066 37136 22094
rect 37004 21956 37056 21962
rect 37004 21898 37056 21904
rect 37016 21554 37044 21898
rect 37004 21548 37056 21554
rect 37004 21490 37056 21496
rect 36912 21480 36964 21486
rect 36912 21422 36964 21428
rect 36912 20800 36964 20806
rect 37108 20788 37136 22066
rect 37200 20806 37228 24210
rect 37280 22772 37332 22778
rect 37280 22714 37332 22720
rect 37292 21962 37320 22714
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37384 21894 37412 24210
rect 37568 24070 37596 24618
rect 37660 24138 37688 24618
rect 37648 24132 37700 24138
rect 37648 24074 37700 24080
rect 37556 24064 37608 24070
rect 37660 24041 37688 24074
rect 37556 24006 37608 24012
rect 37646 24032 37702 24041
rect 37646 23967 37702 23976
rect 37464 23316 37516 23322
rect 37464 23258 37516 23264
rect 37476 22778 37504 23258
rect 37648 23112 37700 23118
rect 37648 23054 37700 23060
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37660 22710 37688 23054
rect 37844 22982 37872 26302
rect 38290 26302 38424 26330
rect 38290 26200 38346 26302
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38292 23180 38344 23186
rect 38292 23122 38344 23128
rect 37832 22976 37884 22982
rect 37832 22918 37884 22924
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 38304 22778 38332 23122
rect 38292 22772 38344 22778
rect 38292 22714 38344 22720
rect 37648 22704 37700 22710
rect 37648 22646 37700 22652
rect 37462 22536 37518 22545
rect 37462 22471 37518 22480
rect 37476 22234 37504 22471
rect 37464 22228 37516 22234
rect 37464 22170 37516 22176
rect 37464 22024 37516 22030
rect 37660 22012 37688 22646
rect 37832 22160 37884 22166
rect 37832 22102 37884 22108
rect 37740 22024 37792 22030
rect 37660 21984 37740 22012
rect 37464 21966 37516 21972
rect 37740 21966 37792 21972
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 37280 21548 37332 21554
rect 37280 21490 37332 21496
rect 37292 21457 37320 21490
rect 37278 21448 37334 21457
rect 37384 21418 37412 21830
rect 37278 21383 37334 21392
rect 37372 21412 37424 21418
rect 37372 21354 37424 21360
rect 37384 21162 37412 21354
rect 37292 21134 37412 21162
rect 36964 20760 37136 20788
rect 37188 20800 37240 20806
rect 36912 20742 36964 20748
rect 37188 20742 37240 20748
rect 36924 20058 36952 20742
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 36912 20052 36964 20058
rect 36912 19994 36964 20000
rect 36924 19514 36952 19994
rect 36912 19508 36964 19514
rect 36912 19450 36964 19456
rect 36912 19168 36964 19174
rect 36912 19110 36964 19116
rect 36924 19009 36952 19110
rect 36910 19000 36966 19009
rect 36910 18935 36966 18944
rect 37200 18902 37228 20402
rect 37292 19310 37320 21134
rect 37476 20602 37504 21966
rect 37740 21684 37792 21690
rect 37740 21626 37792 21632
rect 37556 21480 37608 21486
rect 37556 21422 37608 21428
rect 37568 21350 37596 21422
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37568 21010 37596 21286
rect 37556 21004 37608 21010
rect 37556 20946 37608 20952
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37372 20528 37424 20534
rect 37372 20470 37424 20476
rect 37384 19514 37412 20470
rect 37464 20392 37516 20398
rect 37464 20334 37516 20340
rect 37372 19508 37424 19514
rect 37372 19450 37424 19456
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37372 19236 37424 19242
rect 37372 19178 37424 19184
rect 37384 19122 37412 19178
rect 37292 19094 37412 19122
rect 37188 18896 37240 18902
rect 37188 18838 37240 18844
rect 37096 18828 37148 18834
rect 37096 18770 37148 18776
rect 36820 18420 36872 18426
rect 36820 18362 36872 18368
rect 36728 18148 36780 18154
rect 36728 18090 36780 18096
rect 36636 17536 36688 17542
rect 36636 17478 36688 17484
rect 36452 17060 36504 17066
rect 36452 17002 36504 17008
rect 36728 16992 36780 16998
rect 36728 16934 36780 16940
rect 36360 16788 36412 16794
rect 36360 16730 36412 16736
rect 36544 16448 36596 16454
rect 36544 16390 36596 16396
rect 36268 16040 36320 16046
rect 36268 15982 36320 15988
rect 36452 15360 36504 15366
rect 36452 15302 36504 15308
rect 36360 15088 36412 15094
rect 36360 15030 36412 15036
rect 36372 14822 36400 15030
rect 36360 14816 36412 14822
rect 36360 14758 36412 14764
rect 36174 14648 36230 14657
rect 36174 14583 36230 14592
rect 36358 14648 36414 14657
rect 36358 14583 36360 14592
rect 36004 13926 36124 13954
rect 36188 13938 36216 14583
rect 36412 14583 36414 14592
rect 36360 14554 36412 14560
rect 35992 13864 36044 13870
rect 35992 13806 36044 13812
rect 35900 13728 35952 13734
rect 35900 13670 35952 13676
rect 35806 13424 35862 13433
rect 35806 13359 35862 13368
rect 35820 12918 35848 13359
rect 35808 12912 35860 12918
rect 35808 12854 35860 12860
rect 35728 11898 35848 11914
rect 35440 11892 35492 11898
rect 35728 11892 35860 11898
rect 35728 11886 35808 11892
rect 35440 11834 35492 11840
rect 35808 11834 35860 11840
rect 35532 11824 35584 11830
rect 35900 11824 35952 11830
rect 35584 11784 35756 11812
rect 35532 11766 35584 11772
rect 35624 11552 35676 11558
rect 35728 11540 35756 11784
rect 35900 11766 35952 11772
rect 35808 11552 35860 11558
rect 35728 11512 35808 11540
rect 35624 11494 35676 11500
rect 35808 11494 35860 11500
rect 35164 11076 35216 11082
rect 35164 11018 35216 11024
rect 35256 10736 35308 10742
rect 35256 10678 35308 10684
rect 35268 10606 35296 10678
rect 35636 10674 35664 11494
rect 35912 11150 35940 11766
rect 36004 11558 36032 13806
rect 36096 13682 36124 13926
rect 36176 13932 36228 13938
rect 36176 13874 36228 13880
rect 36360 13932 36412 13938
rect 36360 13874 36412 13880
rect 36268 13864 36320 13870
rect 36268 13806 36320 13812
rect 36096 13654 36216 13682
rect 36084 12912 36136 12918
rect 36084 12854 36136 12860
rect 35992 11552 36044 11558
rect 35992 11494 36044 11500
rect 35900 11144 35952 11150
rect 35900 11086 35952 11092
rect 36096 11082 36124 12854
rect 36188 11694 36216 13654
rect 36280 13530 36308 13806
rect 36268 13524 36320 13530
rect 36268 13466 36320 13472
rect 36372 13394 36400 13874
rect 36360 13388 36412 13394
rect 36360 13330 36412 13336
rect 36464 13274 36492 15302
rect 36372 13258 36492 13274
rect 36360 13252 36492 13258
rect 36412 13246 36492 13252
rect 36360 13194 36412 13200
rect 36556 12918 36584 16390
rect 36636 14340 36688 14346
rect 36636 14282 36688 14288
rect 36648 14249 36676 14282
rect 36634 14240 36690 14249
rect 36634 14175 36690 14184
rect 36648 13870 36676 14175
rect 36740 14006 36768 16934
rect 36832 16658 36860 18362
rect 37108 18154 37136 18770
rect 37188 18284 37240 18290
rect 37188 18226 37240 18232
rect 37096 18148 37148 18154
rect 37096 18090 37148 18096
rect 37004 18080 37056 18086
rect 37004 18022 37056 18028
rect 37016 17610 37044 18022
rect 37004 17604 37056 17610
rect 37004 17546 37056 17552
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 36832 15910 36860 16594
rect 37004 16448 37056 16454
rect 37004 16390 37056 16396
rect 36820 15904 36872 15910
rect 36820 15846 36872 15852
rect 37016 15201 37044 16390
rect 37200 16250 37228 18226
rect 37292 18086 37320 19094
rect 37370 19000 37426 19009
rect 37370 18935 37426 18944
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37384 17921 37412 18935
rect 37476 18358 37504 20334
rect 37568 19718 37596 20946
rect 37648 20800 37700 20806
rect 37648 20742 37700 20748
rect 37660 20398 37688 20742
rect 37648 20392 37700 20398
rect 37648 20334 37700 20340
rect 37752 20346 37780 21626
rect 37844 21350 37872 22102
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 38396 21690 38424 26302
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 42154 26330 42210 27000
rect 42154 26302 42748 26330
rect 42154 26200 42210 26302
rect 38844 24200 38896 24206
rect 38844 24142 38896 24148
rect 38568 24064 38620 24070
rect 38752 24064 38804 24070
rect 38620 24024 38700 24052
rect 38568 24006 38620 24012
rect 38568 23520 38620 23526
rect 38568 23462 38620 23468
rect 38580 23202 38608 23462
rect 38672 23361 38700 24024
rect 38752 24006 38804 24012
rect 38658 23352 38714 23361
rect 38658 23287 38714 23296
rect 38580 23186 38700 23202
rect 38580 23180 38712 23186
rect 38580 23174 38660 23180
rect 38660 23122 38712 23128
rect 38660 23044 38712 23050
rect 38660 22986 38712 22992
rect 38672 22794 38700 22986
rect 38580 22766 38700 22794
rect 38580 22438 38608 22766
rect 38660 22704 38712 22710
rect 38660 22646 38712 22652
rect 38568 22432 38620 22438
rect 38568 22374 38620 22380
rect 38672 22234 38700 22646
rect 38660 22228 38712 22234
rect 38660 22170 38712 22176
rect 38476 22092 38528 22098
rect 38672 22080 38700 22170
rect 38528 22052 38700 22080
rect 38476 22034 38528 22040
rect 38384 21684 38436 21690
rect 38384 21626 38436 21632
rect 38292 21616 38344 21622
rect 38568 21616 38620 21622
rect 38344 21564 38424 21570
rect 38292 21558 38424 21564
rect 38568 21558 38620 21564
rect 38304 21542 38424 21558
rect 38396 21486 38424 21542
rect 38292 21480 38344 21486
rect 38292 21422 38344 21428
rect 38384 21480 38436 21486
rect 38384 21422 38436 21428
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37844 20806 37872 21286
rect 38304 21185 38332 21422
rect 38290 21176 38346 21185
rect 38290 21111 38346 21120
rect 38384 20868 38436 20874
rect 38580 20856 38608 21558
rect 38764 21049 38792 24006
rect 38856 23798 38884 24142
rect 38844 23792 38896 23798
rect 38844 23734 38896 23740
rect 38856 23225 38884 23734
rect 38842 23216 38898 23225
rect 38842 23151 38898 23160
rect 38844 22772 38896 22778
rect 38844 22714 38896 22720
rect 38856 22098 38884 22714
rect 38948 22438 38976 26200
rect 39592 25022 39620 26200
rect 39580 25016 39632 25022
rect 39580 24958 39632 24964
rect 40038 24712 40094 24721
rect 40038 24647 40094 24656
rect 40052 24614 40080 24647
rect 39856 24608 39908 24614
rect 39856 24550 39908 24556
rect 40040 24608 40092 24614
rect 40040 24550 40092 24556
rect 39488 24404 39540 24410
rect 39488 24346 39540 24352
rect 39394 24304 39450 24313
rect 39394 24239 39450 24248
rect 39408 24206 39436 24239
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39304 24064 39356 24070
rect 39304 24006 39356 24012
rect 39212 23588 39264 23594
rect 39212 23530 39264 23536
rect 39120 23520 39172 23526
rect 39120 23462 39172 23468
rect 39028 23316 39080 23322
rect 39028 23258 39080 23264
rect 39040 23225 39068 23258
rect 39026 23216 39082 23225
rect 39026 23151 39082 23160
rect 39132 23050 39160 23462
rect 39120 23044 39172 23050
rect 39120 22986 39172 22992
rect 39132 22953 39160 22986
rect 39118 22944 39174 22953
rect 39118 22879 39174 22888
rect 38936 22432 38988 22438
rect 38936 22374 38988 22380
rect 38844 22092 38896 22098
rect 38844 22034 38896 22040
rect 39224 21434 39252 23530
rect 39316 23089 39344 24006
rect 39408 23526 39436 24142
rect 39500 23594 39528 24346
rect 39672 24336 39724 24342
rect 39672 24278 39724 24284
rect 39580 23724 39632 23730
rect 39580 23666 39632 23672
rect 39488 23588 39540 23594
rect 39488 23530 39540 23536
rect 39396 23520 39448 23526
rect 39396 23462 39448 23468
rect 39488 23180 39540 23186
rect 39488 23122 39540 23128
rect 39302 23080 39358 23089
rect 39302 23015 39358 23024
rect 39500 22778 39528 23122
rect 39592 23089 39620 23666
rect 39578 23080 39634 23089
rect 39578 23015 39634 23024
rect 39488 22772 39540 22778
rect 39488 22714 39540 22720
rect 39500 22166 39528 22714
rect 39488 22160 39540 22166
rect 39488 22102 39540 22108
rect 39224 21418 39344 21434
rect 39224 21412 39356 21418
rect 39224 21406 39304 21412
rect 38750 21040 38806 21049
rect 38750 20975 38806 20984
rect 38436 20828 38608 20856
rect 38384 20810 38436 20816
rect 37832 20800 37884 20806
rect 37832 20742 37884 20748
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37924 20528 37976 20534
rect 38396 20516 38424 20810
rect 37976 20488 38424 20516
rect 37924 20470 37976 20476
rect 37752 20318 37872 20346
rect 37648 20256 37700 20262
rect 37648 20198 37700 20204
rect 37740 20256 37792 20262
rect 37740 20198 37792 20204
rect 37556 19712 37608 19718
rect 37556 19654 37608 19660
rect 37568 18630 37596 19654
rect 37660 19009 37688 20198
rect 37752 19242 37780 20198
rect 37844 20058 37872 20318
rect 39224 20262 39252 21406
rect 39304 21354 39356 21360
rect 39500 21010 39528 22102
rect 39580 21888 39632 21894
rect 39580 21830 39632 21836
rect 39488 21004 39540 21010
rect 39488 20946 39540 20952
rect 39500 20466 39528 20946
rect 39488 20460 39540 20466
rect 39488 20402 39540 20408
rect 39212 20256 39264 20262
rect 39212 20198 39264 20204
rect 37832 20052 37884 20058
rect 37832 19994 37884 20000
rect 37844 19854 37872 19994
rect 38384 19916 38436 19922
rect 38384 19858 38436 19864
rect 39396 19916 39448 19922
rect 39396 19858 39448 19864
rect 37832 19848 37884 19854
rect 38200 19848 38252 19854
rect 37832 19790 37884 19796
rect 38198 19816 38200 19825
rect 38252 19816 38254 19825
rect 38198 19751 38254 19760
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37924 19508 37976 19514
rect 37924 19450 37976 19456
rect 37740 19236 37792 19242
rect 37740 19178 37792 19184
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 37646 19000 37702 19009
rect 37646 18935 37702 18944
rect 37740 18896 37792 18902
rect 37740 18838 37792 18844
rect 37648 18760 37700 18766
rect 37648 18702 37700 18708
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37568 18426 37596 18566
rect 37556 18420 37608 18426
rect 37556 18362 37608 18368
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37370 17912 37426 17921
rect 37370 17847 37426 17856
rect 37280 17740 37332 17746
rect 37280 17682 37332 17688
rect 37188 16244 37240 16250
rect 37188 16186 37240 16192
rect 37292 16046 37320 17682
rect 37372 17604 37424 17610
rect 37372 17546 37424 17552
rect 37384 16232 37412 17546
rect 37476 16454 37504 18022
rect 37568 17678 37596 18362
rect 37556 17672 37608 17678
rect 37556 17614 37608 17620
rect 37568 16726 37596 17614
rect 37556 16720 37608 16726
rect 37556 16662 37608 16668
rect 37464 16448 37516 16454
rect 37464 16390 37516 16396
rect 37384 16204 37596 16232
rect 37372 16108 37424 16114
rect 37372 16050 37424 16056
rect 37280 16040 37332 16046
rect 37280 15982 37332 15988
rect 37292 15706 37320 15982
rect 37280 15700 37332 15706
rect 37280 15642 37332 15648
rect 37384 15570 37412 16050
rect 37464 16040 37516 16046
rect 37464 15982 37516 15988
rect 37476 15638 37504 15982
rect 37464 15632 37516 15638
rect 37464 15574 37516 15580
rect 37372 15564 37424 15570
rect 37372 15506 37424 15512
rect 37002 15192 37058 15201
rect 37002 15127 37058 15136
rect 36820 14816 36872 14822
rect 36820 14758 36872 14764
rect 36832 14618 36860 14758
rect 36820 14612 36872 14618
rect 36820 14554 36872 14560
rect 36728 14000 36780 14006
rect 36728 13942 36780 13948
rect 36636 13864 36688 13870
rect 36636 13806 36688 13812
rect 36648 13258 36676 13806
rect 36820 13388 36872 13394
rect 36820 13330 36872 13336
rect 36636 13252 36688 13258
rect 36636 13194 36688 13200
rect 36544 12912 36596 12918
rect 36544 12854 36596 12860
rect 36832 12850 36860 13330
rect 36912 12912 36964 12918
rect 36912 12854 36964 12860
rect 36820 12844 36872 12850
rect 36820 12786 36872 12792
rect 36924 12646 36952 12854
rect 37016 12782 37044 15127
rect 37384 15026 37412 15506
rect 37372 15020 37424 15026
rect 37372 14962 37424 14968
rect 37096 14952 37148 14958
rect 37096 14894 37148 14900
rect 37004 12776 37056 12782
rect 37004 12718 37056 12724
rect 37016 12646 37044 12718
rect 36912 12640 36964 12646
rect 36912 12582 36964 12588
rect 37004 12640 37056 12646
rect 37004 12582 37056 12588
rect 36728 12096 36780 12102
rect 36728 12038 36780 12044
rect 36176 11688 36228 11694
rect 36176 11630 36228 11636
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 36452 11144 36504 11150
rect 36504 11104 36584 11132
rect 36452 11086 36504 11092
rect 36084 11076 36136 11082
rect 36084 11018 36136 11024
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35716 10668 35768 10674
rect 35716 10610 35768 10616
rect 35256 10600 35308 10606
rect 34978 10568 35034 10577
rect 35728 10554 35756 10610
rect 35256 10542 35308 10548
rect 34978 10503 35034 10512
rect 35636 10526 35756 10554
rect 35636 10130 35664 10526
rect 35716 10260 35768 10266
rect 35716 10202 35768 10208
rect 35728 10130 35756 10202
rect 35624 10124 35676 10130
rect 35624 10066 35676 10072
rect 35716 10124 35768 10130
rect 35716 10066 35768 10072
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 35636 9722 35664 10066
rect 35624 9716 35676 9722
rect 35624 9658 35676 9664
rect 36096 9518 36124 11018
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36084 9512 36136 9518
rect 36084 9454 36136 9460
rect 35164 9376 35216 9382
rect 35164 9318 35216 9324
rect 35176 9042 35204 9318
rect 36372 9178 36400 10542
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 35164 9036 35216 9042
rect 35164 8978 35216 8984
rect 35624 8832 35676 8838
rect 35624 8774 35676 8780
rect 35636 8566 35664 8774
rect 35624 8560 35676 8566
rect 35624 8502 35676 8508
rect 36464 8430 36492 10610
rect 36556 10606 36584 11104
rect 36544 10600 36596 10606
rect 36544 10542 36596 10548
rect 36556 10062 36584 10542
rect 36648 10538 36676 11630
rect 36740 11558 36768 12038
rect 36820 11756 36872 11762
rect 36820 11698 36872 11704
rect 36728 11552 36780 11558
rect 36728 11494 36780 11500
rect 36832 10810 36860 11698
rect 36820 10804 36872 10810
rect 36820 10746 36872 10752
rect 36912 10600 36964 10606
rect 36912 10542 36964 10548
rect 36636 10532 36688 10538
rect 36636 10474 36688 10480
rect 36648 10266 36676 10474
rect 36924 10266 36952 10542
rect 36636 10260 36688 10266
rect 36636 10202 36688 10208
rect 36912 10260 36964 10266
rect 36912 10202 36964 10208
rect 36544 10056 36596 10062
rect 36544 9998 36596 10004
rect 36556 9722 36584 9998
rect 36544 9716 36596 9722
rect 36544 9658 36596 9664
rect 36452 8424 36504 8430
rect 36452 8366 36504 8372
rect 34796 7948 34848 7954
rect 34796 7890 34848 7896
rect 36820 6384 36872 6390
rect 36820 6326 36872 6332
rect 36452 6180 36504 6186
rect 36452 6122 36504 6128
rect 36464 3466 36492 6122
rect 36832 4826 36860 6326
rect 36820 4820 36872 4826
rect 36820 4762 36872 4768
rect 36832 4622 36860 4762
rect 37016 4690 37044 12582
rect 37108 9178 37136 14894
rect 37384 14482 37412 14962
rect 37568 14550 37596 16204
rect 37660 15094 37688 18702
rect 37752 18426 37780 18838
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 37844 18222 37872 19110
rect 37936 18834 37964 19450
rect 38014 19272 38070 19281
rect 38014 19207 38070 19216
rect 38028 18902 38056 19207
rect 38016 18896 38068 18902
rect 38016 18838 38068 18844
rect 37924 18828 37976 18834
rect 37924 18770 37976 18776
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 38396 18442 38424 19858
rect 38476 19712 38528 19718
rect 38476 19654 38528 19660
rect 38304 18414 38424 18442
rect 38016 18352 38068 18358
rect 38016 18294 38068 18300
rect 37924 18284 37976 18290
rect 37924 18226 37976 18232
rect 37740 18216 37792 18222
rect 37740 18158 37792 18164
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 37752 15706 37780 18158
rect 37844 17134 37872 18158
rect 37936 18154 37964 18226
rect 38028 18154 38056 18294
rect 37924 18148 37976 18154
rect 37924 18090 37976 18096
rect 38016 18148 38068 18154
rect 38016 18090 38068 18096
rect 37936 17678 37964 18090
rect 37924 17672 37976 17678
rect 37924 17614 37976 17620
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 37740 15700 37792 15706
rect 37740 15642 37792 15648
rect 37752 15094 37780 15642
rect 37648 15088 37700 15094
rect 37648 15030 37700 15036
rect 37740 15088 37792 15094
rect 37740 15030 37792 15036
rect 37844 14958 37872 16594
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 38304 14958 38332 18414
rect 38384 17876 38436 17882
rect 38384 17818 38436 17824
rect 38396 17134 38424 17818
rect 38384 17128 38436 17134
rect 38384 17070 38436 17076
rect 38488 15314 38516 19654
rect 39408 19310 39436 19858
rect 39500 19446 39528 20402
rect 39592 19718 39620 21830
rect 39684 21010 39712 24278
rect 39868 23798 39896 24550
rect 40132 24132 40184 24138
rect 40132 24074 40184 24080
rect 40040 24064 40092 24070
rect 40040 24006 40092 24012
rect 40052 23866 40080 24006
rect 40040 23860 40092 23866
rect 40040 23802 40092 23808
rect 39764 23792 39816 23798
rect 39764 23734 39816 23740
rect 39856 23792 39908 23798
rect 39856 23734 39908 23740
rect 39776 23662 39804 23734
rect 39764 23656 39816 23662
rect 39764 23598 39816 23604
rect 39762 23352 39818 23361
rect 39762 23287 39818 23296
rect 39948 23316 40000 23322
rect 39776 22778 39804 23287
rect 39948 23258 40000 23264
rect 39960 23118 39988 23258
rect 39948 23112 40000 23118
rect 39948 23054 40000 23060
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 39948 22976 40000 22982
rect 39948 22918 40000 22924
rect 39764 22772 39816 22778
rect 39764 22714 39816 22720
rect 39672 21004 39724 21010
rect 39672 20946 39724 20952
rect 39776 20534 39804 22714
rect 39960 21978 39988 22918
rect 40052 22817 40080 23054
rect 40144 22982 40172 24074
rect 40132 22976 40184 22982
rect 40132 22918 40184 22924
rect 40038 22808 40094 22817
rect 40236 22794 40264 26200
rect 40960 24948 41012 24954
rect 40960 24890 41012 24896
rect 40408 24880 40460 24886
rect 40408 24822 40460 24828
rect 40316 24268 40368 24274
rect 40316 24210 40368 24216
rect 40038 22743 40094 22752
rect 40144 22766 40264 22794
rect 40144 22438 40172 22766
rect 40224 22636 40276 22642
rect 40224 22578 40276 22584
rect 40040 22432 40092 22438
rect 40040 22374 40092 22380
rect 40132 22432 40184 22438
rect 40132 22374 40184 22380
rect 39868 21950 39988 21978
rect 39868 21894 39896 21950
rect 39856 21888 39908 21894
rect 39856 21830 39908 21836
rect 39948 21888 40000 21894
rect 39948 21830 40000 21836
rect 39868 21690 39896 21830
rect 39856 21684 39908 21690
rect 39856 21626 39908 21632
rect 39764 20528 39816 20534
rect 39764 20470 39816 20476
rect 39672 20460 39724 20466
rect 39672 20402 39724 20408
rect 39580 19712 39632 19718
rect 39580 19654 39632 19660
rect 39592 19514 39620 19654
rect 39580 19508 39632 19514
rect 39580 19450 39632 19456
rect 39488 19440 39540 19446
rect 39684 19417 39712 20402
rect 39854 20224 39910 20233
rect 39854 20159 39910 20168
rect 39868 19417 39896 20159
rect 39960 20058 39988 21830
rect 40052 21486 40080 22374
rect 40040 21480 40092 21486
rect 40040 21422 40092 21428
rect 40236 20806 40264 22578
rect 40328 21146 40356 24210
rect 40316 21140 40368 21146
rect 40316 21082 40368 21088
rect 40224 20800 40276 20806
rect 40224 20742 40276 20748
rect 40236 20584 40264 20742
rect 40236 20556 40356 20584
rect 40132 20392 40184 20398
rect 40132 20334 40184 20340
rect 39948 20052 40000 20058
rect 39948 19994 40000 20000
rect 40040 19780 40092 19786
rect 40040 19722 40092 19728
rect 40052 19514 40080 19722
rect 40040 19508 40092 19514
rect 40040 19450 40092 19456
rect 39488 19382 39540 19388
rect 39670 19408 39726 19417
rect 39670 19343 39726 19352
rect 39854 19408 39910 19417
rect 39854 19343 39910 19352
rect 39396 19304 39448 19310
rect 39396 19246 39448 19252
rect 39408 18970 39436 19246
rect 40040 19168 40092 19174
rect 40040 19110 40092 19116
rect 39396 18964 39448 18970
rect 39396 18906 39448 18912
rect 38568 18828 38620 18834
rect 38568 18770 38620 18776
rect 38580 16454 38608 18770
rect 40052 18766 40080 19110
rect 40040 18760 40092 18766
rect 40040 18702 40092 18708
rect 39764 18692 39816 18698
rect 39764 18634 39816 18640
rect 39776 18290 39804 18634
rect 39948 18624 40000 18630
rect 39948 18566 40000 18572
rect 39764 18284 39816 18290
rect 39764 18226 39816 18232
rect 39960 17882 39988 18566
rect 40052 18086 40080 18702
rect 40144 18630 40172 20334
rect 40224 19848 40276 19854
rect 40224 19790 40276 19796
rect 40236 19242 40264 19790
rect 40224 19236 40276 19242
rect 40224 19178 40276 19184
rect 40132 18624 40184 18630
rect 40132 18566 40184 18572
rect 40224 18624 40276 18630
rect 40224 18566 40276 18572
rect 40040 18080 40092 18086
rect 40040 18022 40092 18028
rect 39948 17876 40000 17882
rect 39948 17818 40000 17824
rect 40052 17746 40080 18022
rect 40040 17740 40092 17746
rect 40040 17682 40092 17688
rect 38660 17672 38712 17678
rect 38660 17614 38712 17620
rect 38844 17672 38896 17678
rect 38844 17614 38896 17620
rect 38672 17270 38700 17614
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 38672 16522 38700 17206
rect 38856 16998 38884 17614
rect 38936 17536 38988 17542
rect 38936 17478 38988 17484
rect 38948 17202 38976 17478
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 38844 16992 38896 16998
rect 38844 16934 38896 16940
rect 38856 16658 38884 16934
rect 38844 16652 38896 16658
rect 38844 16594 38896 16600
rect 38660 16516 38712 16522
rect 38660 16458 38712 16464
rect 38568 16448 38620 16454
rect 38568 16390 38620 16396
rect 38580 16182 38608 16390
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38672 15450 38700 16458
rect 38672 15434 38792 15450
rect 38660 15428 38792 15434
rect 38712 15422 38792 15428
rect 38660 15370 38712 15376
rect 38488 15286 38700 15314
rect 38672 15162 38700 15286
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38764 15094 38792 15422
rect 38752 15088 38804 15094
rect 38752 15030 38804 15036
rect 37832 14952 37884 14958
rect 37832 14894 37884 14900
rect 38292 14952 38344 14958
rect 38292 14894 38344 14900
rect 37556 14544 37608 14550
rect 37556 14486 37608 14492
rect 37280 14476 37332 14482
rect 37280 14418 37332 14424
rect 37372 14476 37424 14482
rect 37372 14418 37424 14424
rect 37292 12434 37320 14418
rect 38304 14346 38332 14894
rect 38764 14770 38792 15030
rect 38672 14742 38792 14770
rect 38292 14340 38344 14346
rect 38292 14282 38344 14288
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 38672 14006 38700 14742
rect 38752 14612 38804 14618
rect 38752 14554 38804 14560
rect 38660 14000 38712 14006
rect 38660 13942 38712 13948
rect 38200 13796 38252 13802
rect 38200 13738 38252 13744
rect 38212 13530 38240 13738
rect 38200 13524 38252 13530
rect 38200 13466 38252 13472
rect 38212 13274 38240 13466
rect 38212 13246 38332 13274
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37648 13184 37700 13190
rect 37648 13126 37700 13132
rect 37476 12850 37504 13126
rect 37660 12918 37688 13126
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37648 12912 37700 12918
rect 37648 12854 37700 12860
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 37292 12406 37412 12434
rect 37384 12306 37412 12406
rect 37372 12300 37424 12306
rect 37372 12242 37424 12248
rect 37372 11824 37424 11830
rect 37372 11766 37424 11772
rect 37188 11620 37240 11626
rect 37188 11562 37240 11568
rect 37200 11082 37228 11562
rect 37384 11218 37412 11766
rect 37476 11218 37504 12786
rect 38304 12782 38332 13246
rect 38292 12776 38344 12782
rect 38292 12718 38344 12724
rect 38764 12306 38792 14554
rect 38844 14000 38896 14006
rect 38844 13942 38896 13948
rect 38856 13530 38884 13942
rect 38844 13524 38896 13530
rect 38844 13466 38896 13472
rect 38856 12850 38884 13466
rect 38844 12844 38896 12850
rect 38844 12786 38896 12792
rect 38856 12442 38884 12786
rect 38844 12436 38896 12442
rect 38844 12378 38896 12384
rect 38384 12300 38436 12306
rect 38384 12242 38436 12248
rect 38752 12300 38804 12306
rect 38752 12242 38804 12248
rect 37556 12096 37608 12102
rect 37556 12038 37608 12044
rect 37372 11212 37424 11218
rect 37372 11154 37424 11160
rect 37464 11212 37516 11218
rect 37464 11154 37516 11160
rect 37188 11076 37240 11082
rect 37188 11018 37240 11024
rect 37568 10538 37596 12038
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 38396 11082 38424 12242
rect 38660 12096 38712 12102
rect 38660 12038 38712 12044
rect 38672 11898 38700 12038
rect 38660 11892 38712 11898
rect 38660 11834 38712 11840
rect 38856 11286 38884 12378
rect 38844 11280 38896 11286
rect 38844 11222 38896 11228
rect 38384 11076 38436 11082
rect 38384 11018 38436 11024
rect 38568 11008 38620 11014
rect 38568 10950 38620 10956
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 38580 10742 38608 10950
rect 38568 10736 38620 10742
rect 38568 10678 38620 10684
rect 38948 10674 38976 17138
rect 40052 16998 40080 17682
rect 40144 17270 40172 18566
rect 40236 18154 40264 18566
rect 40328 18329 40356 20556
rect 40420 19854 40448 24822
rect 40592 24744 40644 24750
rect 40592 24686 40644 24692
rect 40604 24274 40632 24686
rect 40592 24268 40644 24274
rect 40592 24210 40644 24216
rect 40776 24064 40828 24070
rect 40776 24006 40828 24012
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 40696 23497 40724 23598
rect 40682 23488 40738 23497
rect 40604 23446 40682 23474
rect 40500 22976 40552 22982
rect 40500 22918 40552 22924
rect 40512 22234 40540 22918
rect 40500 22228 40552 22234
rect 40500 22170 40552 22176
rect 40500 22092 40552 22098
rect 40604 22094 40632 23446
rect 40682 23423 40738 23432
rect 40682 23216 40738 23225
rect 40682 23151 40684 23160
rect 40736 23151 40738 23160
rect 40684 23122 40736 23128
rect 40604 22066 40724 22094
rect 40500 22034 40552 22040
rect 40512 21865 40540 22034
rect 40498 21856 40554 21865
rect 40498 21791 40554 21800
rect 40512 21457 40540 21791
rect 40592 21616 40644 21622
rect 40592 21558 40644 21564
rect 40498 21448 40554 21457
rect 40498 21383 40554 21392
rect 40512 20058 40540 21383
rect 40604 20924 40632 21558
rect 40696 21078 40724 22066
rect 40788 21622 40816 24006
rect 40972 23746 41000 24890
rect 41234 24848 41290 24857
rect 41234 24783 41290 24792
rect 41052 24676 41104 24682
rect 41052 24618 41104 24624
rect 41064 24410 41092 24618
rect 41052 24404 41104 24410
rect 41052 24346 41104 24352
rect 41064 23866 41092 24346
rect 41248 24138 41276 24783
rect 42524 24404 42576 24410
rect 42524 24346 42576 24352
rect 41236 24132 41288 24138
rect 41236 24074 41288 24080
rect 41052 23860 41104 23866
rect 41052 23802 41104 23808
rect 40972 23718 41092 23746
rect 40960 23656 41012 23662
rect 40960 23598 41012 23604
rect 40868 22976 40920 22982
rect 40866 22944 40868 22953
rect 40920 22944 40922 22953
rect 40866 22879 40922 22888
rect 40868 22704 40920 22710
rect 40868 22646 40920 22652
rect 40880 22438 40908 22646
rect 40868 22432 40920 22438
rect 40868 22374 40920 22380
rect 40972 22098 41000 23598
rect 40960 22092 41012 22098
rect 40960 22034 41012 22040
rect 40866 21992 40922 22001
rect 40866 21927 40922 21936
rect 40960 21956 41012 21962
rect 40880 21622 40908 21927
rect 40960 21898 41012 21904
rect 40776 21616 40828 21622
rect 40776 21558 40828 21564
rect 40868 21616 40920 21622
rect 40868 21558 40920 21564
rect 40880 21486 40908 21558
rect 40868 21480 40920 21486
rect 40868 21422 40920 21428
rect 40972 21418 41000 21898
rect 40960 21412 41012 21418
rect 40960 21354 41012 21360
rect 40868 21344 40920 21350
rect 40868 21286 40920 21292
rect 40684 21072 40736 21078
rect 40684 21014 40736 21020
rect 40684 20936 40736 20942
rect 40604 20896 40684 20924
rect 40684 20878 40736 20884
rect 40880 20806 40908 21286
rect 40868 20800 40920 20806
rect 40868 20742 40920 20748
rect 41064 20398 41092 23718
rect 42064 23588 42116 23594
rect 42064 23530 42116 23536
rect 41328 23112 41380 23118
rect 41328 23054 41380 23060
rect 41340 22642 41368 23054
rect 41418 22808 41474 22817
rect 41418 22743 41474 22752
rect 41328 22636 41380 22642
rect 41328 22578 41380 22584
rect 41236 22432 41288 22438
rect 41236 22374 41288 22380
rect 41144 22092 41196 22098
rect 41144 22034 41196 22040
rect 41052 20392 41104 20398
rect 41052 20334 41104 20340
rect 40684 20256 40736 20262
rect 40684 20198 40736 20204
rect 40500 20052 40552 20058
rect 40500 19994 40552 20000
rect 40512 19922 40540 19994
rect 40500 19916 40552 19922
rect 40500 19858 40552 19864
rect 40408 19848 40460 19854
rect 40408 19790 40460 19796
rect 40314 18320 40370 18329
rect 40314 18255 40370 18264
rect 40224 18148 40276 18154
rect 40224 18090 40276 18096
rect 40222 17912 40278 17921
rect 40222 17847 40278 17856
rect 40592 17876 40644 17882
rect 40132 17264 40184 17270
rect 40132 17206 40184 17212
rect 40040 16992 40092 16998
rect 39960 16952 40040 16980
rect 39488 16584 39540 16590
rect 39488 16526 39540 16532
rect 39212 16040 39264 16046
rect 39212 15982 39264 15988
rect 39224 15434 39252 15982
rect 39500 15570 39528 16526
rect 39960 16182 39988 16952
rect 40040 16934 40092 16940
rect 40236 16794 40264 17847
rect 40592 17818 40644 17824
rect 40604 17338 40632 17818
rect 40696 17746 40724 20198
rect 40868 19712 40920 19718
rect 40868 19654 40920 19660
rect 40880 18426 40908 19654
rect 41064 19514 41092 20334
rect 41052 19508 41104 19514
rect 41052 19450 41104 19456
rect 41052 19304 41104 19310
rect 41052 19246 41104 19252
rect 41064 19174 41092 19246
rect 41052 19168 41104 19174
rect 41052 19110 41104 19116
rect 40868 18420 40920 18426
rect 40868 18362 40920 18368
rect 41156 18193 41184 22034
rect 41248 20913 41276 22374
rect 41340 21706 41368 22578
rect 41432 22234 41460 22743
rect 42076 22642 42104 23530
rect 42432 23520 42484 23526
rect 42430 23488 42432 23497
rect 42484 23488 42486 23497
rect 42430 23423 42486 23432
rect 42444 23225 42472 23423
rect 42430 23216 42486 23225
rect 42430 23151 42486 23160
rect 42064 22636 42116 22642
rect 42064 22578 42116 22584
rect 41880 22432 41932 22438
rect 41878 22400 41880 22409
rect 41932 22400 41934 22409
rect 41878 22335 41934 22344
rect 41420 22228 41472 22234
rect 41420 22170 41472 22176
rect 42064 22160 42116 22166
rect 42064 22102 42116 22108
rect 41880 22092 41932 22098
rect 41880 22034 41932 22040
rect 41512 22024 41564 22030
rect 41512 21966 41564 21972
rect 41524 21894 41552 21966
rect 41512 21888 41564 21894
rect 41512 21830 41564 21836
rect 41340 21678 41460 21706
rect 41432 21350 41460 21678
rect 41892 21486 41920 22034
rect 42076 21690 42104 22102
rect 42156 22092 42208 22098
rect 42156 22034 42208 22040
rect 42168 21894 42196 22034
rect 42536 22030 42564 24346
rect 42720 24290 42748 26302
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26200 45430 27000
rect 46018 26330 46074 27000
rect 46018 26302 46336 26330
rect 46018 26200 46074 26302
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 42720 24262 42840 24290
rect 42812 24206 42840 24262
rect 42800 24200 42852 24206
rect 42800 24142 42852 24148
rect 43352 24200 43404 24206
rect 43352 24142 43404 24148
rect 42800 23656 42852 23662
rect 42800 23598 42852 23604
rect 42812 23338 42840 23598
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42720 23310 42840 23338
rect 42720 23050 42748 23310
rect 42800 23180 42852 23186
rect 42800 23122 42852 23128
rect 42708 23044 42760 23050
rect 42708 22986 42760 22992
rect 42614 22672 42670 22681
rect 42614 22607 42616 22616
rect 42668 22607 42670 22616
rect 42616 22578 42668 22584
rect 42720 22166 42748 22986
rect 42708 22160 42760 22166
rect 42708 22102 42760 22108
rect 42524 22024 42576 22030
rect 42524 21966 42576 21972
rect 42156 21888 42208 21894
rect 42156 21830 42208 21836
rect 42248 21888 42300 21894
rect 42248 21830 42300 21836
rect 42064 21684 42116 21690
rect 42064 21626 42116 21632
rect 41512 21480 41564 21486
rect 41512 21422 41564 21428
rect 41880 21480 41932 21486
rect 41880 21422 41932 21428
rect 41420 21344 41472 21350
rect 41420 21286 41472 21292
rect 41328 20936 41380 20942
rect 41234 20904 41290 20913
rect 41328 20878 41380 20884
rect 41234 20839 41290 20848
rect 41234 19136 41290 19145
rect 41234 19071 41290 19080
rect 41142 18184 41198 18193
rect 41142 18119 41198 18128
rect 40868 17808 40920 17814
rect 40868 17750 40920 17756
rect 40684 17740 40736 17746
rect 40684 17682 40736 17688
rect 40592 17332 40644 17338
rect 40592 17274 40644 17280
rect 40684 17128 40736 17134
rect 40684 17070 40736 17076
rect 40224 16788 40276 16794
rect 40224 16730 40276 16736
rect 40236 16522 40264 16730
rect 40316 16652 40368 16658
rect 40316 16594 40368 16600
rect 40224 16516 40276 16522
rect 40224 16458 40276 16464
rect 39948 16176 40000 16182
rect 39948 16118 40000 16124
rect 39488 15564 39540 15570
rect 39488 15506 39540 15512
rect 39302 15464 39358 15473
rect 39212 15428 39264 15434
rect 39960 15434 39988 16118
rect 40328 15910 40356 16594
rect 40696 16590 40724 17070
rect 40684 16584 40736 16590
rect 40684 16526 40736 16532
rect 40316 15904 40368 15910
rect 40316 15846 40368 15852
rect 40328 15570 40356 15846
rect 40316 15564 40368 15570
rect 40316 15506 40368 15512
rect 39302 15399 39358 15408
rect 39948 15428 40000 15434
rect 39212 15370 39264 15376
rect 39224 13462 39252 15370
rect 39316 14414 39344 15399
rect 39948 15370 40000 15376
rect 39396 14952 39448 14958
rect 39396 14894 39448 14900
rect 39304 14408 39356 14414
rect 39304 14350 39356 14356
rect 39408 14278 39436 14894
rect 39960 14618 39988 15370
rect 40880 15026 40908 17750
rect 41052 16992 41104 16998
rect 41052 16934 41104 16940
rect 41064 16794 41092 16934
rect 41248 16794 41276 19071
rect 41052 16788 41104 16794
rect 41052 16730 41104 16736
rect 41236 16788 41288 16794
rect 41236 16730 41288 16736
rect 41064 16658 41092 16730
rect 41052 16652 41104 16658
rect 41052 16594 41104 16600
rect 41248 16522 41276 16730
rect 41236 16516 41288 16522
rect 41236 16458 41288 16464
rect 40960 16448 41012 16454
rect 40960 16390 41012 16396
rect 40972 16250 41000 16390
rect 40960 16244 41012 16250
rect 40960 16186 41012 16192
rect 41340 15609 41368 20878
rect 41524 20097 41552 21422
rect 41602 21176 41658 21185
rect 42260 21146 42288 21830
rect 42536 21690 42564 21966
rect 42524 21684 42576 21690
rect 42524 21626 42576 21632
rect 42812 21146 42840 23122
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42982 22128 43038 22137
rect 42982 22063 43038 22072
rect 43260 22092 43312 22098
rect 42996 22030 43024 22063
rect 43260 22034 43312 22040
rect 42984 22024 43036 22030
rect 42984 21966 43036 21972
rect 43272 21894 43300 22034
rect 43260 21888 43312 21894
rect 43260 21830 43312 21836
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 43364 21146 43392 24142
rect 43628 24064 43680 24070
rect 43628 24006 43680 24012
rect 43720 24064 43772 24070
rect 43720 24006 43772 24012
rect 43536 23520 43588 23526
rect 43536 23462 43588 23468
rect 43548 23050 43576 23462
rect 43536 23044 43588 23050
rect 43536 22986 43588 22992
rect 43444 22500 43496 22506
rect 43444 22442 43496 22448
rect 43456 21593 43484 22442
rect 43536 22432 43588 22438
rect 43536 22374 43588 22380
rect 43548 22234 43576 22374
rect 43536 22228 43588 22234
rect 43536 22170 43588 22176
rect 43548 21865 43576 22170
rect 43534 21856 43590 21865
rect 43534 21791 43590 21800
rect 43442 21584 43498 21593
rect 43442 21519 43498 21528
rect 43444 21344 43496 21350
rect 43444 21286 43496 21292
rect 41602 21111 41658 21120
rect 42248 21140 42300 21146
rect 41616 20942 41644 21111
rect 42248 21082 42300 21088
rect 42800 21140 42852 21146
rect 42800 21082 42852 21088
rect 43352 21140 43404 21146
rect 43352 21082 43404 21088
rect 42708 21072 42760 21078
rect 42708 21014 42760 21020
rect 41972 21004 42024 21010
rect 41708 20964 41972 20992
rect 41604 20936 41656 20942
rect 41604 20878 41656 20884
rect 41604 20800 41656 20806
rect 41708 20788 41736 20964
rect 41972 20946 42024 20952
rect 41788 20868 41840 20874
rect 41788 20810 41840 20816
rect 42064 20868 42116 20874
rect 42064 20810 42116 20816
rect 41656 20760 41736 20788
rect 41604 20742 41656 20748
rect 41800 20618 41828 20810
rect 42076 20754 42104 20810
rect 41984 20726 42104 20754
rect 41984 20618 42012 20726
rect 41800 20590 42012 20618
rect 41510 20088 41566 20097
rect 41510 20023 41566 20032
rect 42720 19854 42748 21014
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 43456 19990 43484 21286
rect 43640 20806 43668 24006
rect 43732 23769 43760 24006
rect 43718 23760 43774 23769
rect 43718 23695 43774 23704
rect 43996 23724 44048 23730
rect 43996 23666 44048 23672
rect 44008 23322 44036 23666
rect 43996 23316 44048 23322
rect 43996 23258 44048 23264
rect 43994 23216 44050 23225
rect 43994 23151 43996 23160
rect 44048 23151 44050 23160
rect 43996 23122 44048 23128
rect 43720 22976 43772 22982
rect 43720 22918 43772 22924
rect 43732 22710 43760 22918
rect 44100 22710 44128 26200
rect 44364 24812 44416 24818
rect 44364 24754 44416 24760
rect 44376 24070 44404 24754
rect 44548 24608 44600 24614
rect 44548 24550 44600 24556
rect 44560 24206 44588 24550
rect 44548 24200 44600 24206
rect 44548 24142 44600 24148
rect 44364 24064 44416 24070
rect 44364 24006 44416 24012
rect 44560 23662 44588 24142
rect 44548 23656 44600 23662
rect 44548 23598 44600 23604
rect 44744 23050 44772 26200
rect 45388 24698 45416 26200
rect 45744 25016 45796 25022
rect 45744 24958 45796 24964
rect 45388 24670 45600 24698
rect 45572 23798 45600 24670
rect 45560 23792 45612 23798
rect 45560 23734 45612 23740
rect 44732 23044 44784 23050
rect 44732 22986 44784 22992
rect 45376 23044 45428 23050
rect 45376 22986 45428 22992
rect 43720 22704 43772 22710
rect 43720 22646 43772 22652
rect 44088 22704 44140 22710
rect 44088 22646 44140 22652
rect 44272 22704 44324 22710
rect 44272 22646 44324 22652
rect 44454 22672 44510 22681
rect 43720 22568 43772 22574
rect 43720 22510 43772 22516
rect 43732 22094 43760 22510
rect 43732 22066 43944 22094
rect 43720 22024 43772 22030
rect 43720 21966 43772 21972
rect 43812 22024 43864 22030
rect 43812 21966 43864 21972
rect 43732 21690 43760 21966
rect 43720 21684 43772 21690
rect 43720 21626 43772 21632
rect 43824 21486 43852 21966
rect 43812 21480 43864 21486
rect 43812 21422 43864 21428
rect 43628 20800 43680 20806
rect 43628 20742 43680 20748
rect 43444 19984 43496 19990
rect 43444 19926 43496 19932
rect 42708 19848 42760 19854
rect 42708 19790 42760 19796
rect 42064 19304 42116 19310
rect 42064 19246 42116 19252
rect 42076 18970 42104 19246
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42064 18964 42116 18970
rect 42064 18906 42116 18912
rect 42708 18896 42760 18902
rect 42708 18838 42760 18844
rect 41970 17776 42026 17785
rect 41970 17711 42026 17720
rect 41984 16726 42012 17711
rect 42720 17241 42748 18838
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42706 17232 42762 17241
rect 42706 17167 42762 17176
rect 43916 17066 43944 22066
rect 44088 22024 44140 22030
rect 44088 21966 44140 21972
rect 44100 18737 44128 21966
rect 44284 21690 44312 22646
rect 44454 22607 44510 22616
rect 45192 22636 45244 22642
rect 44468 21690 44496 22607
rect 45192 22578 45244 22584
rect 45204 22234 45232 22578
rect 45388 22234 45416 22986
rect 45756 22642 45784 24958
rect 46308 24682 46336 26302
rect 46662 26200 46718 27000
rect 47306 26330 47362 27000
rect 47228 26302 47362 26330
rect 46296 24676 46348 24682
rect 46296 24618 46348 24624
rect 46480 24336 46532 24342
rect 46480 24278 46532 24284
rect 46020 24064 46072 24070
rect 46020 24006 46072 24012
rect 45928 23724 45980 23730
rect 45928 23666 45980 23672
rect 45744 22636 45796 22642
rect 45744 22578 45796 22584
rect 45558 22536 45614 22545
rect 45558 22471 45560 22480
rect 45612 22471 45614 22480
rect 45560 22442 45612 22448
rect 45756 22234 45784 22578
rect 45192 22228 45244 22234
rect 45192 22170 45244 22176
rect 45376 22228 45428 22234
rect 45376 22170 45428 22176
rect 45744 22228 45796 22234
rect 45744 22170 45796 22176
rect 45100 22092 45152 22098
rect 45100 22034 45152 22040
rect 45112 21894 45140 22034
rect 45100 21888 45152 21894
rect 45100 21830 45152 21836
rect 45940 21690 45968 23666
rect 46032 23050 46060 24006
rect 46112 23520 46164 23526
rect 46110 23488 46112 23497
rect 46164 23488 46166 23497
rect 46110 23423 46166 23432
rect 46492 23118 46520 24278
rect 46572 24064 46624 24070
rect 46572 24006 46624 24012
rect 46584 23186 46612 24006
rect 46572 23180 46624 23186
rect 46572 23122 46624 23128
rect 46676 23118 46704 26200
rect 47030 24304 47086 24313
rect 47030 24239 47086 24248
rect 46756 23860 46808 23866
rect 46756 23802 46808 23808
rect 46768 23254 46796 23802
rect 46756 23248 46808 23254
rect 46756 23190 46808 23196
rect 46480 23112 46532 23118
rect 46480 23054 46532 23060
rect 46664 23112 46716 23118
rect 46664 23054 46716 23060
rect 46846 23080 46902 23089
rect 46020 23044 46072 23050
rect 46846 23015 46902 23024
rect 46020 22986 46072 22992
rect 44272 21684 44324 21690
rect 44272 21626 44324 21632
rect 44456 21684 44508 21690
rect 44456 21626 44508 21632
rect 45928 21684 45980 21690
rect 45928 21626 45980 21632
rect 46032 20874 46060 22986
rect 46860 22234 46888 23015
rect 46940 22976 46992 22982
rect 46940 22918 46992 22924
rect 46848 22228 46900 22234
rect 46848 22170 46900 22176
rect 46112 22024 46164 22030
rect 46112 21966 46164 21972
rect 46124 21486 46152 21966
rect 46112 21480 46164 21486
rect 46112 21422 46164 21428
rect 46020 20868 46072 20874
rect 46020 20810 46072 20816
rect 46952 20369 46980 22918
rect 47044 22778 47072 24239
rect 47124 24132 47176 24138
rect 47124 24074 47176 24080
rect 47136 23866 47164 24074
rect 47124 23860 47176 23866
rect 47124 23802 47176 23808
rect 47122 23624 47178 23633
rect 47122 23559 47178 23568
rect 47032 22772 47084 22778
rect 47032 22714 47084 22720
rect 47136 20942 47164 23559
rect 47228 22642 47256 26302
rect 47306 26200 47362 26302
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 49238 26200 49294 27000
rect 47490 25120 47546 25129
rect 47490 25055 47546 25064
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 47320 23050 47348 23802
rect 47400 23588 47452 23594
rect 47400 23530 47452 23536
rect 47308 23044 47360 23050
rect 47308 22986 47360 22992
rect 47216 22636 47268 22642
rect 47216 22578 47268 22584
rect 47412 21554 47440 23530
rect 47504 22030 47532 25055
rect 47582 24712 47638 24721
rect 47582 24647 47638 24656
rect 47768 24676 47820 24682
rect 47596 23633 47624 24647
rect 47768 24618 47820 24624
rect 47780 24138 47808 24618
rect 47964 24154 47992 26200
rect 47768 24132 47820 24138
rect 47768 24074 47820 24080
rect 47872 24126 47992 24154
rect 47780 23798 47808 24074
rect 47768 23792 47820 23798
rect 47768 23734 47820 23740
rect 47582 23624 47638 23633
rect 47582 23559 47638 23568
rect 47766 23624 47822 23633
rect 47766 23559 47822 23568
rect 47676 23520 47728 23526
rect 47582 23488 47638 23497
rect 47676 23462 47728 23468
rect 47582 23423 47638 23432
rect 47596 22234 47624 23423
rect 47688 23118 47716 23462
rect 47676 23112 47728 23118
rect 47676 23054 47728 23060
rect 47676 22976 47728 22982
rect 47676 22918 47728 22924
rect 47688 22658 47716 22918
rect 47780 22778 47808 23559
rect 47768 22772 47820 22778
rect 47768 22714 47820 22720
rect 47688 22630 47808 22658
rect 47676 22568 47728 22574
rect 47676 22510 47728 22516
rect 47584 22228 47636 22234
rect 47584 22170 47636 22176
rect 47492 22024 47544 22030
rect 47492 21966 47544 21972
rect 47596 21962 47624 22170
rect 47584 21956 47636 21962
rect 47584 21898 47636 21904
rect 47688 21622 47716 22510
rect 47676 21616 47728 21622
rect 47676 21558 47728 21564
rect 47400 21548 47452 21554
rect 47400 21490 47452 21496
rect 47780 21146 47808 22630
rect 47872 21962 47900 24126
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 48608 23866 48636 26200
rect 49054 25528 49110 25537
rect 49054 25463 49110 25472
rect 49068 24206 49096 25463
rect 49252 24698 49280 26200
rect 49252 24670 49372 24698
rect 49238 24304 49294 24313
rect 49238 24239 49294 24248
rect 49056 24200 49108 24206
rect 49056 24142 49108 24148
rect 49146 24168 49202 24177
rect 48596 23860 48648 23866
rect 48596 23802 48648 23808
rect 48780 23724 48832 23730
rect 48780 23666 48832 23672
rect 47952 23520 48004 23526
rect 47952 23462 48004 23468
rect 47964 22982 47992 23462
rect 48792 23322 48820 23666
rect 49068 23526 49096 24142
rect 49146 24103 49202 24112
rect 49160 24070 49188 24103
rect 49148 24064 49200 24070
rect 49148 24006 49200 24012
rect 49056 23520 49108 23526
rect 49056 23462 49108 23468
rect 49252 23322 49280 24239
rect 49344 24070 49372 24670
rect 49332 24064 49384 24070
rect 49332 24006 49384 24012
rect 49344 23866 49372 24006
rect 49332 23860 49384 23866
rect 49332 23802 49384 23808
rect 48780 23316 48832 23322
rect 48780 23258 48832 23264
rect 49240 23316 49292 23322
rect 49240 23258 49292 23264
rect 48594 23080 48650 23089
rect 48594 23015 48596 23024
rect 48648 23015 48650 23024
rect 48596 22986 48648 22992
rect 47952 22976 48004 22982
rect 47952 22918 48004 22924
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48608 22778 48636 22986
rect 48596 22772 48648 22778
rect 48596 22714 48648 22720
rect 48226 22672 48282 22681
rect 49252 22642 49280 23258
rect 49332 22976 49384 22982
rect 49332 22918 49384 22924
rect 48226 22607 48282 22616
rect 49240 22636 49292 22642
rect 47860 21956 47912 21962
rect 48240 21944 48268 22607
rect 49240 22578 49292 22584
rect 48412 22432 48464 22438
rect 48412 22374 48464 22380
rect 48504 22432 48556 22438
rect 48504 22374 48556 22380
rect 48240 21916 48360 21944
rect 47860 21898 47912 21904
rect 47872 21690 47900 21898
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47860 21684 47912 21690
rect 47860 21626 47912 21632
rect 48332 21570 48360 21916
rect 48240 21554 48360 21570
rect 48228 21548 48360 21554
rect 48280 21542 48360 21548
rect 48228 21490 48280 21496
rect 48320 21344 48372 21350
rect 48320 21286 48372 21292
rect 47768 21140 47820 21146
rect 47768 21082 47820 21088
rect 47124 20936 47176 20942
rect 47124 20878 47176 20884
rect 47860 20936 47912 20942
rect 47860 20878 47912 20884
rect 47872 20602 47900 20878
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47860 20596 47912 20602
rect 47860 20538 47912 20544
rect 46938 20360 46994 20369
rect 46938 20295 46994 20304
rect 48332 20262 48360 21286
rect 48424 20346 48452 22374
rect 48516 22094 48544 22374
rect 48516 22066 48636 22094
rect 48424 20318 48544 20346
rect 48320 20256 48372 20262
rect 48320 20198 48372 20204
rect 48412 20256 48464 20262
rect 48412 20198 48464 20204
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 48424 19446 48452 20198
rect 48516 19961 48544 20318
rect 48502 19952 48558 19961
rect 48502 19887 48558 19896
rect 48412 19440 48464 19446
rect 48412 19382 48464 19388
rect 48608 18873 48636 22066
rect 49240 21956 49292 21962
rect 49240 21898 49292 21904
rect 48780 21888 48832 21894
rect 48778 21856 48780 21865
rect 48872 21888 48924 21894
rect 48832 21856 48834 21865
rect 48872 21830 48924 21836
rect 48778 21791 48834 21800
rect 48792 20942 48820 21791
rect 48780 20936 48832 20942
rect 48780 20878 48832 20884
rect 48780 20460 48832 20466
rect 48780 20402 48832 20408
rect 48792 20233 48820 20402
rect 48778 20224 48834 20233
rect 48778 20159 48834 20168
rect 48792 20058 48820 20159
rect 48780 20052 48832 20058
rect 48780 19994 48832 20000
rect 48884 19417 48912 21830
rect 49252 21486 49280 21898
rect 49344 21554 49372 22918
rect 49424 22568 49476 22574
rect 49424 22510 49476 22516
rect 49436 22273 49464 22510
rect 49422 22264 49478 22273
rect 49422 22199 49478 22208
rect 49332 21548 49384 21554
rect 49332 21490 49384 21496
rect 49240 21480 49292 21486
rect 49238 21448 49240 21457
rect 49292 21448 49294 21457
rect 49238 21383 49294 21392
rect 49344 21049 49372 21490
rect 49330 21040 49386 21049
rect 49330 20975 49386 20984
rect 49332 20936 49384 20942
rect 49332 20878 49384 20884
rect 49344 20641 49372 20878
rect 49330 20632 49386 20641
rect 49330 20567 49386 20576
rect 49424 20460 49476 20466
rect 49424 20402 49476 20408
rect 49436 19825 49464 20402
rect 49422 19816 49478 19825
rect 49332 19780 49384 19786
rect 49422 19751 49478 19760
rect 49332 19722 49384 19728
rect 49148 19712 49200 19718
rect 49148 19654 49200 19660
rect 48870 19408 48926 19417
rect 48870 19343 48926 19352
rect 49160 19281 49188 19654
rect 49344 19417 49372 19722
rect 49330 19408 49386 19417
rect 49240 19372 49292 19378
rect 49330 19343 49386 19352
rect 49240 19314 49292 19320
rect 49146 19272 49202 19281
rect 49146 19207 49202 19216
rect 49252 19009 49280 19314
rect 49424 19168 49476 19174
rect 49424 19110 49476 19116
rect 49238 19000 49294 19009
rect 49238 18935 49294 18944
rect 48594 18864 48650 18873
rect 48594 18799 48650 18808
rect 49436 18766 49464 19110
rect 48780 18760 48832 18766
rect 44086 18728 44142 18737
rect 48780 18702 48832 18708
rect 49424 18760 49476 18766
rect 49424 18702 49476 18708
rect 44086 18663 44142 18672
rect 48412 18624 48464 18630
rect 48792 18601 48820 18702
rect 48412 18566 48464 18572
rect 48778 18592 48834 18601
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 48424 18358 48452 18566
rect 48778 18527 48834 18536
rect 48792 18426 48820 18527
rect 48780 18420 48832 18426
rect 48780 18362 48832 18368
rect 48412 18352 48464 18358
rect 48412 18294 48464 18300
rect 49332 18284 49384 18290
rect 49332 18226 49384 18232
rect 49148 18080 49200 18086
rect 49148 18022 49200 18028
rect 49160 17882 49188 18022
rect 49148 17876 49200 17882
rect 49148 17818 49200 17824
rect 49344 17785 49372 18226
rect 49436 18193 49464 18702
rect 49422 18184 49478 18193
rect 49422 18119 49478 18128
rect 49330 17776 49386 17785
rect 49330 17711 49386 17720
rect 49332 17672 49384 17678
rect 49332 17614 49384 17620
rect 48412 17604 48464 17610
rect 48412 17546 48464 17552
rect 49240 17604 49292 17610
rect 49240 17546 49292 17552
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48424 17338 48452 17546
rect 49148 17536 49200 17542
rect 49148 17478 49200 17484
rect 48412 17332 48464 17338
rect 48412 17274 48464 17280
rect 48780 17196 48832 17202
rect 48780 17138 48832 17144
rect 43904 17060 43956 17066
rect 43904 17002 43956 17008
rect 48792 16969 48820 17138
rect 49056 17128 49108 17134
rect 49054 17096 49056 17105
rect 49108 17096 49110 17105
rect 49054 17031 49110 17040
rect 48778 16960 48834 16969
rect 42950 16892 43258 16901
rect 48778 16895 48834 16904
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 48792 16794 48820 16895
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 41972 16720 42024 16726
rect 49160 16697 49188 17478
rect 49252 17218 49280 17546
rect 49344 17377 49372 17614
rect 49330 17368 49386 17377
rect 49330 17303 49386 17312
rect 49252 17202 49372 17218
rect 49252 17196 49384 17202
rect 49252 17190 49332 17196
rect 49332 17138 49384 17144
rect 41972 16662 42024 16668
rect 49146 16688 49202 16697
rect 49146 16623 49202 16632
rect 41604 16584 41656 16590
rect 49344 16561 49372 17138
rect 49424 16584 49476 16590
rect 41604 16526 41656 16532
rect 49146 16552 49202 16561
rect 41616 15910 41644 16526
rect 49146 16487 49202 16496
rect 49330 16552 49386 16561
rect 49424 16526 49476 16532
rect 49330 16487 49386 16496
rect 49160 16454 49188 16487
rect 49148 16448 49200 16454
rect 49148 16390 49200 16396
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 49436 16153 49464 16526
rect 49422 16144 49478 16153
rect 48688 16108 48740 16114
rect 48688 16050 48740 16056
rect 49332 16108 49384 16114
rect 49422 16079 49478 16088
rect 49332 16050 49384 16056
rect 41788 16040 41840 16046
rect 41788 15982 41840 15988
rect 41604 15904 41656 15910
rect 41604 15846 41656 15852
rect 41800 15706 41828 15982
rect 42064 15904 42116 15910
rect 42064 15846 42116 15852
rect 42076 15706 42104 15846
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 48700 15706 48728 16050
rect 49146 16008 49202 16017
rect 49146 15943 49148 15952
rect 49200 15943 49202 15952
rect 49148 15914 49200 15920
rect 49344 15745 49372 16050
rect 49330 15736 49386 15745
rect 41788 15700 41840 15706
rect 41788 15642 41840 15648
rect 42064 15700 42116 15706
rect 42064 15642 42116 15648
rect 48688 15700 48740 15706
rect 49330 15671 49386 15680
rect 48688 15642 48740 15648
rect 41326 15600 41382 15609
rect 41326 15535 41382 15544
rect 49332 15496 49384 15502
rect 49332 15438 49384 15444
rect 49344 15337 49372 15438
rect 49330 15328 49386 15337
rect 47950 15260 48258 15269
rect 49330 15263 49386 15272
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 48412 15088 48464 15094
rect 48412 15030 48464 15036
rect 48870 15056 48926 15065
rect 40868 15020 40920 15026
rect 40868 14962 40920 14968
rect 45652 14816 45704 14822
rect 45652 14758 45704 14764
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 39948 14612 40000 14618
rect 39948 14554 40000 14560
rect 39396 14272 39448 14278
rect 39396 14214 39448 14220
rect 39488 14272 39540 14278
rect 39488 14214 39540 14220
rect 39500 14006 39528 14214
rect 41328 14068 41380 14074
rect 41328 14010 41380 14016
rect 39488 14000 39540 14006
rect 39488 13942 39540 13948
rect 39212 13456 39264 13462
rect 39212 13398 39264 13404
rect 39488 13388 39540 13394
rect 39488 13330 39540 13336
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39316 12782 39344 13126
rect 39304 12776 39356 12782
rect 39304 12718 39356 12724
rect 39120 12640 39172 12646
rect 39120 12582 39172 12588
rect 39132 11898 39160 12582
rect 39316 12442 39344 12718
rect 39304 12436 39356 12442
rect 39304 12378 39356 12384
rect 39120 11892 39172 11898
rect 39120 11834 39172 11840
rect 39028 11756 39080 11762
rect 39028 11698 39080 11704
rect 38936 10668 38988 10674
rect 38936 10610 38988 10616
rect 37556 10532 37608 10538
rect 37556 10474 37608 10480
rect 38948 10062 38976 10610
rect 38936 10056 38988 10062
rect 38936 9998 38988 10004
rect 37464 9988 37516 9994
rect 37464 9930 37516 9936
rect 37096 9172 37148 9178
rect 37096 9114 37148 9120
rect 37108 8906 37136 9114
rect 37096 8900 37148 8906
rect 37096 8842 37148 8848
rect 37476 8498 37504 9930
rect 38384 9920 38436 9926
rect 38384 9862 38436 9868
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 38396 9722 38424 9862
rect 38384 9716 38436 9722
rect 38384 9658 38436 9664
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 37464 8492 37516 8498
rect 37464 8434 37516 8440
rect 38752 8424 38804 8430
rect 38752 8366 38804 8372
rect 38764 7886 38792 8366
rect 38936 8356 38988 8362
rect 38936 8298 38988 8304
rect 38752 7880 38804 7886
rect 38752 7822 38804 7828
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 38672 7546 38700 7686
rect 38660 7540 38712 7546
rect 38660 7482 38712 7488
rect 38476 7336 38528 7342
rect 38476 7278 38528 7284
rect 37280 7268 37332 7274
rect 37280 7210 37332 7216
rect 37292 5370 37320 7210
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 37936 6934 37964 7142
rect 37924 6928 37976 6934
rect 37924 6870 37976 6876
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37740 6248 37792 6254
rect 37740 6190 37792 6196
rect 37648 6112 37700 6118
rect 37648 6054 37700 6060
rect 37660 5914 37688 6054
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37280 5364 37332 5370
rect 37280 5306 37332 5312
rect 37004 4684 37056 4690
rect 37004 4626 37056 4632
rect 37752 4622 37780 6190
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 38488 5302 38516 7278
rect 38476 5296 38528 5302
rect 38476 5238 38528 5244
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 37844 4826 37872 4966
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 38948 4758 38976 8298
rect 39040 8022 39068 11698
rect 39500 11286 39528 13330
rect 41340 13326 41368 14010
rect 45664 13938 45692 14758
rect 48320 14272 48372 14278
rect 48320 14214 48372 14220
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47860 14068 47912 14074
rect 48332 14056 48360 14214
rect 48424 14074 48452 15030
rect 48870 14991 48926 15000
rect 49332 15020 49384 15026
rect 48884 14074 48912 14991
rect 49332 14962 49384 14968
rect 49344 14929 49372 14962
rect 49146 14920 49202 14929
rect 49146 14855 49148 14864
rect 49200 14855 49202 14864
rect 49330 14920 49386 14929
rect 49330 14855 49386 14864
rect 49148 14826 49200 14832
rect 49056 14544 49108 14550
rect 49054 14512 49056 14521
rect 49108 14512 49110 14521
rect 49054 14447 49110 14456
rect 49238 14512 49294 14521
rect 49238 14447 49294 14456
rect 49252 14414 49280 14447
rect 49240 14408 49292 14414
rect 49240 14350 49292 14356
rect 49238 14104 49294 14113
rect 47860 14010 47912 14016
rect 48240 14028 48360 14056
rect 48412 14068 48464 14074
rect 45652 13932 45704 13938
rect 45652 13874 45704 13880
rect 46572 13864 46624 13870
rect 46572 13806 46624 13812
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 46584 13326 46612 13806
rect 41328 13320 41380 13326
rect 41328 13262 41380 13268
rect 46572 13320 46624 13326
rect 46572 13262 46624 13268
rect 45928 13184 45980 13190
rect 45928 13126 45980 13132
rect 40316 12980 40368 12986
rect 40316 12922 40368 12928
rect 40040 12844 40092 12850
rect 40040 12786 40092 12792
rect 40052 12753 40080 12786
rect 40038 12744 40094 12753
rect 40038 12679 40094 12688
rect 40224 11552 40276 11558
rect 40224 11494 40276 11500
rect 39488 11280 39540 11286
rect 39488 11222 39540 11228
rect 40236 11150 40264 11494
rect 40224 11144 40276 11150
rect 40224 11086 40276 11092
rect 39948 9104 40000 9110
rect 39948 9046 40000 9052
rect 39764 8832 39816 8838
rect 39764 8774 39816 8780
rect 39776 8566 39804 8774
rect 39764 8560 39816 8566
rect 39764 8502 39816 8508
rect 39028 8016 39080 8022
rect 39028 7958 39080 7964
rect 39960 5710 39988 9046
rect 40328 8498 40356 12922
rect 45940 12850 45968 13126
rect 47872 12850 47900 14010
rect 48240 13938 48268 14028
rect 48412 14010 48464 14016
rect 48872 14068 48924 14074
rect 49238 14039 49294 14048
rect 48872 14010 48924 14016
rect 49252 14006 49280 14039
rect 49240 14000 49292 14006
rect 49240 13942 49292 13948
rect 48228 13932 48280 13938
rect 48228 13874 48280 13880
rect 48240 13705 48268 13874
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 49148 13320 49200 13326
rect 49146 13288 49148 13297
rect 49200 13288 49202 13297
rect 49146 13223 49202 13232
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 49146 12880 49202 12889
rect 45928 12844 45980 12850
rect 45928 12786 45980 12792
rect 47860 12844 47912 12850
rect 49146 12815 49148 12824
rect 47860 12786 47912 12792
rect 49200 12815 49202 12824
rect 49148 12786 49200 12792
rect 46756 12708 46808 12714
rect 46756 12650 46808 12656
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 40408 12164 40460 12170
rect 40408 12106 40460 12112
rect 40420 11801 40448 12106
rect 40960 12096 41012 12102
rect 40960 12038 41012 12044
rect 46112 12096 46164 12102
rect 46112 12038 46164 12044
rect 40972 11830 41000 12038
rect 40960 11824 41012 11830
rect 40406 11792 40462 11801
rect 40960 11766 41012 11772
rect 46124 11762 46152 12038
rect 40406 11727 40408 11736
rect 40460 11727 40462 11736
rect 46112 11756 46164 11762
rect 40408 11698 40460 11704
rect 46112 11698 46164 11704
rect 46572 11620 46624 11626
rect 46572 11562 46624 11568
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 44364 11348 44416 11354
rect 44364 11290 44416 11296
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 44376 9994 44404 11290
rect 46112 11008 46164 11014
rect 46112 10950 46164 10956
rect 46124 10062 46152 10950
rect 46584 10062 46612 11562
rect 46768 11150 46796 12650
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 47216 12368 47268 12374
rect 47216 12310 47268 12316
rect 47032 11552 47084 11558
rect 47032 11494 47084 11500
rect 46756 11144 46808 11150
rect 46756 11086 46808 11092
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10674 46980 11018
rect 46940 10668 46992 10674
rect 46940 10610 46992 10616
rect 45836 10056 45888 10062
rect 45836 9998 45888 10004
rect 46112 10056 46164 10062
rect 46112 9998 46164 10004
rect 46572 10056 46624 10062
rect 46572 9998 46624 10004
rect 44364 9988 44416 9994
rect 44364 9930 44416 9936
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 41420 8628 41472 8634
rect 41420 8570 41472 8576
rect 40316 8492 40368 8498
rect 40316 8434 40368 8440
rect 41328 7812 41380 7818
rect 41328 7754 41380 7760
rect 41340 6798 41368 7754
rect 41328 6792 41380 6798
rect 41328 6734 41380 6740
rect 41432 6390 41460 8570
rect 45848 8498 45876 9998
rect 46756 9988 46808 9994
rect 46756 9930 46808 9936
rect 46768 8498 46796 9930
rect 46940 9716 46992 9722
rect 46940 9658 46992 9664
rect 45836 8492 45888 8498
rect 45836 8434 45888 8440
rect 46756 8492 46808 8498
rect 46756 8434 46808 8440
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 44916 8356 44968 8362
rect 44916 8298 44968 8304
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 44928 7478 44956 8298
rect 46860 7993 46888 8366
rect 46846 7984 46902 7993
rect 46846 7919 46902 7928
rect 44916 7472 44968 7478
rect 44916 7414 44968 7420
rect 46952 7410 46980 9658
rect 47044 8974 47072 11494
rect 47124 10532 47176 10538
rect 47124 10474 47176 10480
rect 47032 8968 47084 8974
rect 47032 8910 47084 8916
rect 47136 7886 47164 10474
rect 47228 9586 47256 12310
rect 47964 12238 47992 12582
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49160 12306 49188 12407
rect 49148 12300 49200 12306
rect 49148 12242 49200 12248
rect 47952 12232 48004 12238
rect 47952 12174 48004 12180
rect 49146 12064 49202 12073
rect 47950 11996 48258 12005
rect 49146 11999 49202 12008
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 49160 11830 49188 11999
rect 49148 11824 49200 11830
rect 49148 11766 49200 11772
rect 49146 11656 49202 11665
rect 49146 11591 49202 11600
rect 49160 11218 49188 11591
rect 49238 11248 49294 11257
rect 49148 11212 49200 11218
rect 49238 11183 49294 11192
rect 49148 11154 49200 11160
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 49146 10840 49202 10849
rect 49146 10775 49202 10784
rect 49160 10130 49188 10775
rect 49252 10742 49280 11183
rect 49240 10736 49292 10742
rect 49240 10678 49292 10684
rect 49238 10432 49294 10441
rect 49238 10367 49294 10376
rect 49148 10124 49200 10130
rect 49148 10066 49200 10072
rect 47308 9988 47360 9994
rect 47308 9930 47360 9936
rect 47320 9625 47348 9930
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 49252 9654 49280 10367
rect 49330 10024 49386 10033
rect 49330 9959 49386 9968
rect 49240 9648 49292 9654
rect 47306 9616 47362 9625
rect 47216 9580 47268 9586
rect 49240 9590 49292 9596
rect 47306 9551 47362 9560
rect 47216 9522 47268 9528
rect 49146 9208 49202 9217
rect 49146 9143 49202 9152
rect 47584 8900 47636 8906
rect 47584 8842 47636 8848
rect 47124 7880 47176 7886
rect 47124 7822 47176 7828
rect 47308 7540 47360 7546
rect 47308 7482 47360 7488
rect 46940 7404 46992 7410
rect 46940 7346 46992 7352
rect 45836 7200 45888 7206
rect 45836 7142 45888 7148
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 41420 6384 41472 6390
rect 41420 6326 41472 6332
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 39948 5704 40000 5710
rect 39948 5646 40000 5652
rect 45744 5636 45796 5642
rect 45744 5578 45796 5584
rect 41328 5092 41380 5098
rect 41328 5034 41380 5040
rect 38936 4752 38988 4758
rect 38936 4694 38988 4700
rect 36820 4616 36872 4622
rect 36820 4558 36872 4564
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 39948 4548 40000 4554
rect 39948 4490 40000 4496
rect 37372 4480 37424 4486
rect 37372 4422 37424 4428
rect 37384 4282 37412 4422
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 36452 3460 36504 3466
rect 36452 3402 36504 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 32772 2576 32824 2582
rect 32772 2518 32824 2524
rect 34336 2576 34388 2582
rect 34336 2518 34388 2524
rect 37752 2514 37780 3130
rect 38292 2916 38344 2922
rect 38292 2858 38344 2864
rect 37740 2508 37792 2514
rect 37740 2450 37792 2456
rect 38304 2446 38332 2858
rect 27160 2440 27212 2446
rect 29000 2440 29052 2446
rect 27160 2382 27212 2388
rect 28920 2388 29000 2394
rect 28920 2382 29052 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 38292 2440 38344 2446
rect 38292 2382 38344 2388
rect 28920 2366 29040 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28644 870 28764 898
rect 28644 800 28672 870
rect 18156 734 18368 762
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 28736 762 28764 870
rect 28920 762 28948 2366
rect 30760 800 30788 2382
rect 33152 1578 33180 2382
rect 32876 1550 33180 1578
rect 32876 800 32904 1550
rect 34992 800 35020 2382
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37108 800 37136 2246
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 39224 800 39252 3470
rect 39960 3058 39988 4490
rect 41340 3738 41368 5034
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 45652 4276 45704 4282
rect 45652 4218 45704 4224
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 41328 3732 41380 3738
rect 41328 3674 41380 3680
rect 45560 3460 45612 3466
rect 45560 3402 45612 3408
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 800 41368 2450
rect 43444 2304 43496 2310
rect 43444 2246 43496 2252
rect 43456 800 43484 2246
rect 45572 800 45600 3402
rect 45664 2446 45692 4218
rect 45756 3058 45784 5578
rect 45848 5234 45876 7142
rect 46940 6928 46992 6934
rect 46940 6870 46992 6876
rect 45836 5228 45888 5234
rect 45836 5170 45888 5176
rect 46952 4146 46980 6870
rect 47032 6180 47084 6186
rect 47032 6122 47084 6128
rect 45836 4140 45888 4146
rect 45836 4082 45888 4088
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 45848 3534 45876 4082
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45836 3528 45888 3534
rect 45836 3470 45888 3476
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 45652 2440 45704 2446
rect 45652 2382 45704 2388
rect 46676 1465 46704 4014
rect 47044 3534 47072 6122
rect 47216 5908 47268 5914
rect 47216 5850 47268 5856
rect 47124 4820 47176 4826
rect 47124 4762 47176 4768
rect 47032 3528 47084 3534
rect 47032 3470 47084 3476
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46768 1873 46796 2926
rect 46860 2689 46888 2926
rect 46846 2680 46902 2689
rect 46846 2615 46902 2624
rect 47136 2446 47164 4762
rect 47228 3058 47256 5850
rect 47320 4622 47348 7482
rect 47596 6322 47624 8842
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 49160 8566 49188 9143
rect 49344 9042 49372 9959
rect 49332 9036 49384 9042
rect 49332 8978 49384 8984
rect 49238 8800 49294 8809
rect 49238 8735 49294 8744
rect 47860 8560 47912 8566
rect 47860 8502 47912 8508
rect 49148 8560 49200 8566
rect 49148 8502 49200 8508
rect 47676 8356 47728 8362
rect 47676 8298 47728 8304
rect 47584 6316 47636 6322
rect 47584 6258 47636 6264
rect 47688 5710 47716 8298
rect 47768 7268 47820 7274
rect 47768 7210 47820 7216
rect 47676 5704 47728 5710
rect 47676 5646 47728 5652
rect 47780 5234 47808 7210
rect 47872 6798 47900 8502
rect 49252 7954 49280 8735
rect 49330 8392 49386 8401
rect 49330 8327 49386 8336
rect 49240 7948 49292 7954
rect 49240 7890 49292 7896
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49146 7576 49202 7585
rect 49146 7511 49202 7520
rect 49160 6866 49188 7511
rect 49344 7478 49372 8327
rect 49332 7472 49384 7478
rect 49332 7414 49384 7420
rect 49422 7168 49478 7177
rect 49422 7103 49478 7112
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 47860 6792 47912 6798
rect 47860 6734 47912 6740
rect 49238 6760 49294 6769
rect 48688 6724 48740 6730
rect 49238 6695 49294 6704
rect 48688 6666 48740 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48700 6361 48728 6666
rect 48686 6352 48742 6361
rect 48686 6287 48742 6296
rect 49146 5944 49202 5953
rect 49146 5879 49202 5888
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49160 5302 49188 5879
rect 49252 5778 49280 6695
rect 49436 6390 49464 7103
rect 49424 6384 49476 6390
rect 49424 6326 49476 6332
rect 49240 5772 49292 5778
rect 49240 5714 49292 5720
rect 49422 5536 49478 5545
rect 49422 5471 49478 5480
rect 49148 5296 49200 5302
rect 49148 5238 49200 5244
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 49330 5128 49386 5137
rect 48332 4729 48360 5102
rect 49330 5063 49386 5072
rect 48318 4720 48374 4729
rect 48318 4655 48374 4664
rect 47308 4616 47360 4622
rect 47308 4558 47360 4564
rect 47676 4548 47728 4554
rect 47676 4490 47728 4496
rect 47688 3942 47716 4490
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 47676 3936 47728 3942
rect 47676 3878 47728 3884
rect 47216 3052 47268 3058
rect 47216 2994 47268 3000
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 46754 1864 46810 1873
rect 46754 1799 46810 1808
rect 46662 1456 46718 1465
rect 46662 1391 46718 1400
rect 47688 800 47716 3878
rect 49160 3602 49188 4247
rect 49344 4146 49372 5063
rect 49436 4690 49464 5471
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49792 4480 49844 4486
rect 49792 4422 49844 4428
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49238 3904 49294 3913
rect 49238 3839 49294 3848
rect 49148 3596 49200 3602
rect 49148 3538 49200 3544
rect 49146 3496 49202 3505
rect 48688 3460 48740 3466
rect 49146 3431 49202 3440
rect 48688 3402 48740 3408
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48700 3097 48728 3402
rect 48686 3088 48742 3097
rect 48686 3023 48742 3032
rect 49160 2514 49188 3431
rect 49252 3126 49280 3839
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 2281 48544 2314
rect 48502 2272 48558 2281
rect 47950 2204 48258 2213
rect 48502 2207 48558 2216
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49804 800 49832 4422
rect 28736 734 28948 762
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< via2 >>
rect 3146 25608 3202 25664
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2778 24384 2834 24440
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2962 23160 3018 23216
rect 1766 21528 1822 21584
rect 1030 20712 1086 20768
rect 1306 20304 1362 20360
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3238 21956 3294 21992
rect 3238 21936 3240 21956
rect 3240 21936 3292 21956
rect 3292 21936 3294 21956
rect 3790 25200 3846 25256
rect 3514 23976 3570 24032
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2778 21120 2834 21176
rect 1766 19896 1822 19952
rect 1490 18672 1546 18728
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2870 19488 2926 19544
rect 2778 19080 2834 19136
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3882 24812 3938 24848
rect 3882 24792 3884 24812
rect 3884 24792 3936 24812
rect 3936 24792 3938 24812
rect 3974 23588 4030 23624
rect 3974 23568 3976 23588
rect 3976 23568 4028 23588
rect 4028 23568 4030 23588
rect 3974 22752 4030 22808
rect 1766 18264 1822 18320
rect 4158 22072 4214 22128
rect 1398 17856 1454 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 1766 17448 1822 17504
rect 1030 17040 1086 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 938 16632 994 16688
rect 1030 16224 1086 16280
rect 5354 18808 5410 18864
rect 6550 21548 6606 21584
rect 6550 21528 6552 21548
rect 6552 21528 6604 21548
rect 6604 21528 6606 21548
rect 7470 24248 7526 24304
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8390 20884 8392 20904
rect 8392 20884 8444 20904
rect 8444 20884 8446 20904
rect 8390 20848 8446 20884
rect 9586 21548 9642 21584
rect 9586 21528 9588 21548
rect 9588 21528 9640 21548
rect 9640 21528 9642 21548
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 1030 15816 1086 15872
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 938 15428 994 15464
rect 938 15408 940 15428
rect 940 15408 992 15428
rect 992 15408 994 15428
rect 938 15020 994 15056
rect 938 15000 940 15020
rect 940 15000 992 15020
rect 992 15000 994 15020
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 938 14592 994 14648
rect 1030 14184 1086 14240
rect 1766 13776 1822 13832
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3514 13368 3570 13424
rect 1306 12960 1362 13016
rect 1214 12552 1270 12608
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 1214 12144 1270 12200
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 9862 20460 9918 20496
rect 9862 20440 9864 20460
rect 9864 20440 9916 20460
rect 9916 20440 9918 20460
rect 9954 19352 10010 19408
rect 11334 23024 11390 23080
rect 10782 20324 10838 20360
rect 10782 20304 10784 20324
rect 10784 20304 10836 20324
rect 10836 20304 10838 20324
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 10506 17196 10562 17232
rect 10506 17176 10508 17196
rect 10508 17176 10560 17196
rect 10560 17176 10562 17196
rect 11058 19216 11114 19272
rect 10874 16632 10930 16688
rect 11702 21936 11758 21992
rect 11242 18808 11298 18864
rect 10782 15544 10838 15600
rect 10506 15272 10562 15328
rect 10414 14340 10470 14376
rect 10414 14320 10416 14340
rect 10416 14320 10468 14340
rect 10468 14320 10470 14340
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 1306 11736 1362 11792
rect 1306 11328 1362 11384
rect 1582 10920 1638 10976
rect 1306 10512 1362 10568
rect 1214 10104 1270 10160
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 1306 9716 1362 9752
rect 1306 9696 1308 9716
rect 1308 9696 1360 9716
rect 1360 9696 1362 9716
rect 1766 9444 1822 9480
rect 1766 9424 1768 9444
rect 1768 9424 1820 9444
rect 1820 9424 1822 9444
rect 1306 9288 1362 9344
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 1306 8900 1362 8936
rect 1306 8880 1308 8900
rect 1308 8880 1360 8900
rect 1360 8880 1362 8900
rect 1214 8472 1270 8528
rect 1306 8084 1362 8120
rect 1306 8064 1308 8084
rect 1308 8064 1360 8084
rect 1360 8064 1362 8084
rect 1306 7656 1362 7712
rect 1306 7248 1362 7304
rect 1214 6840 1270 6896
rect 1306 6432 1362 6488
rect 1306 6024 1362 6080
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 1306 4820 1362 4856
rect 1306 4800 1308 4820
rect 1308 4800 1360 4820
rect 1360 4800 1362 4820
rect 1306 4392 1362 4448
rect 1398 3984 1454 4040
rect 1306 3576 1362 3632
rect 1122 3440 1178 3496
rect 1306 3188 1362 3224
rect 1306 3168 1308 3188
rect 1308 3168 1360 3188
rect 1360 3168 1362 3188
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2778 5208 2834 5264
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 11886 19624 11942 19680
rect 11610 16496 11666 16552
rect 11242 13948 11244 13968
rect 11244 13948 11296 13968
rect 11296 13948 11298 13968
rect 11242 13912 11298 13948
rect 11150 13096 11206 13152
rect 11150 12824 11206 12880
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12806 20984 12862 21040
rect 12162 18808 12218 18864
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 11886 17040 11942 17096
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13634 19896 13690 19952
rect 13818 19760 13874 19816
rect 13726 19352 13782 19408
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13174 15952 13230 16008
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 11610 10648 11666 10704
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 5354 3984 5410 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1306 2760 1362 2816
rect 1306 2388 1308 2408
rect 1308 2388 1360 2408
rect 1360 2388 1362 2408
rect 1306 2352 1362 2388
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 1214 1944 1270 2000
rect 1306 1536 1362 1592
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 13910 18264 13966 18320
rect 14278 19488 14334 19544
rect 14922 20304 14978 20360
rect 15474 21528 15530 21584
rect 15290 20304 15346 20360
rect 15198 19372 15254 19408
rect 15198 19352 15200 19372
rect 15200 19352 15252 19372
rect 15252 19352 15254 19372
rect 15566 19252 15568 19272
rect 15568 19252 15620 19272
rect 15620 19252 15622 19272
rect 15566 19216 15622 19252
rect 14462 16768 14518 16824
rect 14002 14456 14058 14512
rect 13450 12688 13506 12744
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13358 11892 13414 11928
rect 13358 11872 13360 11892
rect 13360 11872 13412 11892
rect 13412 11872 13414 11892
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13266 10548 13268 10568
rect 13268 10548 13320 10568
rect 13320 10548 13322 10568
rect 13266 10512 13322 10548
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13726 12688 13782 12744
rect 13818 12144 13874 12200
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 14278 16088 14334 16144
rect 15106 16632 15162 16688
rect 14554 15952 14610 16008
rect 14370 13640 14426 13696
rect 14462 13096 14518 13152
rect 14738 13404 14740 13424
rect 14740 13404 14792 13424
rect 14792 13404 14794 13424
rect 14738 13368 14794 13404
rect 15842 19624 15898 19680
rect 16210 19372 16266 19408
rect 16210 19352 16212 19372
rect 16212 19352 16264 19372
rect 16264 19352 16266 19372
rect 15842 16088 15898 16144
rect 16394 16496 16450 16552
rect 16210 15544 16266 15600
rect 15842 12824 15898 12880
rect 14646 10004 14648 10024
rect 14648 10004 14700 10024
rect 14700 10004 14702 10024
rect 14646 9968 14702 10004
rect 15106 9968 15162 10024
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 16578 14456 16634 14512
rect 16486 13776 16542 13832
rect 16210 12688 16266 12744
rect 17406 20440 17462 20496
rect 17406 18692 17462 18728
rect 17406 18672 17408 18692
rect 17408 18672 17460 18692
rect 17460 18672 17462 18692
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17866 20440 17922 20496
rect 17774 17992 17830 18048
rect 16854 15408 16910 15464
rect 17314 15272 17370 15328
rect 17130 13640 17186 13696
rect 17130 13368 17186 13424
rect 17314 13776 17370 13832
rect 17314 13640 17370 13696
rect 17222 11872 17278 11928
rect 16486 10648 16542 10704
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18694 21936 18750 21992
rect 19798 22616 19854 22672
rect 18602 18808 18658 18864
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18418 15580 18420 15600
rect 18420 15580 18472 15600
rect 18472 15580 18474 15600
rect 18418 15544 18474 15580
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 19338 18692 19394 18728
rect 19338 18672 19340 18692
rect 19340 18672 19392 18692
rect 19392 18672 19394 18692
rect 19338 17992 19394 18048
rect 18970 16768 19026 16824
rect 18510 11076 18566 11112
rect 18510 11056 18512 11076
rect 18512 11056 18564 11076
rect 18564 11056 18566 11076
rect 18786 13232 18842 13288
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 19522 17720 19578 17776
rect 21086 22072 21142 22128
rect 20718 18808 20774 18864
rect 19614 14592 19670 14648
rect 19890 14456 19946 14512
rect 19614 13912 19670 13968
rect 18970 10668 19026 10704
rect 18970 10648 18972 10668
rect 18972 10648 19024 10668
rect 19024 10648 19026 10668
rect 19982 12008 20038 12064
rect 21362 21392 21418 21448
rect 21270 20984 21326 21040
rect 20718 12824 20774 12880
rect 20534 11872 20590 11928
rect 20534 11756 20590 11792
rect 20534 11736 20536 11756
rect 20536 11736 20588 11756
rect 20588 11736 20590 11756
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 21546 20576 21602 20632
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23294 23024 23350 23080
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23754 22208 23810 22264
rect 25778 24284 25780 24304
rect 25780 24284 25832 24304
rect 25832 24284 25834 24304
rect 25778 24248 25834 24284
rect 24214 22072 24270 22128
rect 24766 22480 24822 22536
rect 25318 22924 25320 22944
rect 25320 22924 25372 22944
rect 25372 22924 25374 22944
rect 25318 22888 25374 22924
rect 25134 22344 25190 22400
rect 24858 22108 24860 22128
rect 24860 22108 24912 22128
rect 24912 22108 24914 22128
rect 24858 22072 24914 22108
rect 24858 21936 24914 21992
rect 23754 20848 23810 20904
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23018 19896 23074 19952
rect 21454 15408 21510 15464
rect 21178 14320 21234 14376
rect 21822 15408 21878 15464
rect 22006 14592 22062 14648
rect 22374 17312 22430 17368
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22834 17720 22890 17776
rect 21730 12824 21786 12880
rect 22374 15136 22430 15192
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23846 19916 23902 19952
rect 23846 19896 23848 19916
rect 23848 19896 23900 19916
rect 23900 19896 23902 19916
rect 23662 17992 23718 18048
rect 23662 17176 23718 17232
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22558 14456 22614 14512
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22374 12164 22430 12200
rect 22374 12144 22376 12164
rect 22376 12144 22428 12164
rect 22428 12144 22430 12164
rect 22466 12008 22522 12064
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22466 11056 22522 11112
rect 22926 12980 22982 13016
rect 22926 12960 22928 12980
rect 22928 12960 22980 12980
rect 22980 12960 22982 12980
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23846 14864 23902 14920
rect 25134 20984 25190 21040
rect 25410 20576 25466 20632
rect 25318 20168 25374 20224
rect 25134 19760 25190 19816
rect 25042 19080 25098 19136
rect 25134 18284 25190 18320
rect 25134 18264 25136 18284
rect 25136 18264 25188 18284
rect 25188 18264 25190 18284
rect 25042 18128 25098 18184
rect 24950 16360 25006 16416
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23846 11056 23902 11112
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 25778 21936 25834 21992
rect 25778 20984 25834 21040
rect 26606 24132 26662 24168
rect 26606 24112 26608 24132
rect 26608 24112 26660 24132
rect 26660 24112 26662 24132
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 26606 22092 26662 22128
rect 26606 22072 26608 22092
rect 26608 22072 26660 22092
rect 26660 22072 26662 22092
rect 26422 21412 26478 21448
rect 26422 21392 26424 21412
rect 26424 21392 26476 21412
rect 26476 21392 26478 21412
rect 26054 20324 26110 20360
rect 26054 20304 26056 20324
rect 26056 20304 26108 20324
rect 26108 20304 26110 20324
rect 25962 18264 26018 18320
rect 25962 16632 26018 16688
rect 25962 16496 26018 16552
rect 26238 18128 26294 18184
rect 26238 16396 26240 16416
rect 26240 16396 26292 16416
rect 26292 16396 26294 16416
rect 26238 16360 26294 16396
rect 26238 15020 26294 15056
rect 26238 15000 26240 15020
rect 26240 15000 26292 15020
rect 26292 15000 26294 15020
rect 24950 11736 25006 11792
rect 26422 12980 26478 13016
rect 26422 12960 26424 12980
rect 26424 12960 26476 12980
rect 26476 12960 26478 12980
rect 26054 12824 26110 12880
rect 27434 20884 27436 20904
rect 27436 20884 27488 20904
rect 27488 20884 27490 20904
rect 27434 20848 27490 20884
rect 27618 21972 27620 21992
rect 27620 21972 27672 21992
rect 27672 21972 27674 21992
rect 27618 21936 27674 21972
rect 28262 22208 28318 22264
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 26974 15408 27030 15464
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 28446 19896 28502 19952
rect 27710 18944 27766 19000
rect 27250 16088 27306 16144
rect 27250 15020 27306 15056
rect 27250 15000 27252 15020
rect 27252 15000 27304 15020
rect 27304 15000 27306 15020
rect 27710 17332 27766 17368
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 29918 23840 29974 23896
rect 30010 23704 30066 23760
rect 28814 21528 28870 21584
rect 28354 18672 28410 18728
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27710 17312 27712 17332
rect 27712 17312 27764 17332
rect 27764 17312 27766 17332
rect 27986 17040 28042 17096
rect 28078 16652 28134 16688
rect 28078 16632 28080 16652
rect 28080 16632 28132 16652
rect 28132 16632 28134 16652
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27526 15156 27582 15192
rect 27526 15136 27528 15156
rect 27528 15136 27580 15156
rect 27580 15136 27582 15156
rect 28538 19080 28594 19136
rect 28446 18128 28502 18184
rect 28354 15544 28410 15600
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 28630 18944 28686 19000
rect 28998 18844 29000 18864
rect 29000 18844 29052 18864
rect 29052 18844 29054 18864
rect 28998 18808 29054 18844
rect 28630 16768 28686 16824
rect 27986 14764 27988 14784
rect 27988 14764 28040 14784
rect 28040 14764 28042 14784
rect 27986 14728 28042 14764
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27434 11872 27490 11928
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27710 11056 27766 11112
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 29642 22616 29698 22672
rect 29734 22344 29790 22400
rect 29918 21664 29974 21720
rect 30010 20984 30066 21040
rect 29826 20848 29882 20904
rect 29642 19488 29698 19544
rect 28538 12688 28594 12744
rect 30194 21936 30250 21992
rect 31114 23704 31170 23760
rect 30654 22636 30710 22672
rect 30654 22616 30656 22636
rect 30656 22616 30708 22636
rect 30708 22616 30710 22636
rect 32494 24792 32550 24848
rect 30378 21528 30434 21584
rect 29918 19216 29974 19272
rect 30102 19352 30158 19408
rect 30102 19116 30104 19136
rect 30104 19116 30156 19136
rect 30156 19116 30158 19136
rect 30102 19080 30158 19116
rect 30010 18808 30066 18864
rect 29642 15952 29698 16008
rect 30102 18128 30158 18184
rect 30010 17448 30066 17504
rect 30102 15952 30158 16008
rect 30378 19624 30434 19680
rect 30378 17448 30434 17504
rect 29642 11736 29698 11792
rect 30378 14764 30380 14784
rect 30380 14764 30432 14784
rect 30432 14764 30434 14784
rect 30378 14728 30434 14764
rect 31206 21564 31208 21584
rect 31208 21564 31260 21584
rect 31260 21564 31262 21584
rect 31206 21528 31262 21564
rect 31114 20984 31170 21040
rect 31482 22480 31538 22536
rect 30562 16360 30618 16416
rect 30930 19352 30986 19408
rect 30930 18672 30986 18728
rect 30930 18572 30932 18592
rect 30932 18572 30984 18592
rect 30984 18572 30986 18592
rect 30930 18536 30986 18572
rect 31850 24248 31906 24304
rect 33782 24656 33838 24712
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 31666 23568 31722 23624
rect 33598 23840 33654 23896
rect 32126 22072 32182 22128
rect 31666 20984 31722 21040
rect 31482 19080 31538 19136
rect 31022 17312 31078 17368
rect 30654 15156 30710 15192
rect 30654 15136 30656 15156
rect 30656 15136 30708 15156
rect 30708 15136 30710 15156
rect 31758 20868 31814 20904
rect 31758 20848 31760 20868
rect 31760 20848 31812 20868
rect 31812 20848 31814 20868
rect 32954 23704 33010 23760
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33230 23160 33286 23216
rect 33414 22344 33470 22400
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32586 20848 32642 20904
rect 31942 20324 31998 20360
rect 31942 20304 31944 20324
rect 31944 20304 31996 20324
rect 31996 20304 31998 20324
rect 30562 13232 30618 13288
rect 30102 12144 30158 12200
rect 24858 4020 24860 4040
rect 24860 4020 24912 4040
rect 24912 4020 24914 4040
rect 24858 3984 24914 4020
rect 25778 3440 25834 3496
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 31942 18400 31998 18456
rect 31850 17312 31906 17368
rect 31666 13368 31722 13424
rect 31390 11076 31446 11112
rect 31390 11056 31392 11076
rect 31392 11056 31444 11076
rect 31444 11056 31446 11076
rect 33506 21548 33562 21584
rect 33506 21528 33508 21548
rect 33508 21528 33560 21548
rect 33560 21528 33562 21548
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32402 17312 32458 17368
rect 32402 16360 32458 16416
rect 32310 11056 32366 11112
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32954 18828 33010 18864
rect 32954 18808 32956 18828
rect 32956 18808 33008 18828
rect 33008 18808 33010 18828
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 33598 18844 33600 18864
rect 33600 18844 33652 18864
rect 33652 18844 33654 18864
rect 33598 18808 33654 18844
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 34426 21936 34482 21992
rect 34794 23704 34850 23760
rect 34794 22616 34850 22672
rect 35438 24012 35440 24032
rect 35440 24012 35492 24032
rect 35492 24012 35494 24032
rect 35438 23976 35494 24012
rect 35070 23432 35126 23488
rect 35162 23024 35218 23080
rect 34886 22072 34942 22128
rect 35070 20576 35126 20632
rect 34518 20168 34574 20224
rect 34242 18844 34244 18864
rect 34244 18844 34296 18864
rect 34296 18844 34298 18864
rect 34242 18808 34298 18844
rect 34058 17332 34114 17368
rect 34058 17312 34060 17332
rect 34060 17312 34112 17332
rect 34112 17312 34114 17332
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 34610 15408 34666 15464
rect 35346 22344 35402 22400
rect 35254 20440 35310 20496
rect 35714 22616 35770 22672
rect 36082 23568 36138 23624
rect 36910 24384 36966 24440
rect 35990 21664 36046 21720
rect 34978 18944 35034 19000
rect 35254 18944 35310 19000
rect 34886 16088 34942 16144
rect 33690 9424 33746 9480
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 34426 9560 34482 9616
rect 35162 13252 35218 13288
rect 35162 13232 35164 13252
rect 35164 13232 35216 13252
rect 35216 13232 35218 13252
rect 34702 9596 34704 9616
rect 34704 9596 34756 9616
rect 34756 9596 34758 9616
rect 34702 9560 34758 9596
rect 35530 20576 35586 20632
rect 35530 17484 35532 17504
rect 35532 17484 35584 17504
rect 35584 17484 35586 17504
rect 35530 17448 35586 17484
rect 35714 15952 35770 16008
rect 35438 15272 35494 15328
rect 35438 14184 35494 14240
rect 35898 18400 35954 18456
rect 36726 20576 36782 20632
rect 35714 14320 35770 14376
rect 36634 20032 36690 20088
rect 36634 19488 36690 19544
rect 37094 22208 37150 22264
rect 37646 23976 37702 24032
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37462 22480 37518 22536
rect 37278 21392 37334 21448
rect 36910 18944 36966 19000
rect 36174 14592 36230 14648
rect 36358 14612 36414 14648
rect 36358 14592 36360 14612
rect 36360 14592 36412 14612
rect 36412 14592 36414 14612
rect 35806 13368 35862 13424
rect 36634 14184 36690 14240
rect 37370 18944 37426 19000
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 38658 23296 38714 23352
rect 38290 21120 38346 21176
rect 38842 23160 38898 23216
rect 40038 24656 40094 24712
rect 39394 24248 39450 24304
rect 39026 23160 39082 23216
rect 39118 22888 39174 22944
rect 39302 23024 39358 23080
rect 39578 23024 39634 23080
rect 38750 20984 38806 21040
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 38198 19796 38200 19816
rect 38200 19796 38252 19816
rect 38252 19796 38254 19816
rect 38198 19760 38254 19796
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37646 18944 37702 19000
rect 37370 17856 37426 17912
rect 37002 15136 37058 15192
rect 34978 10512 35034 10568
rect 38014 19216 38070 19272
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 39762 23296 39818 23352
rect 40038 22752 40094 22808
rect 39854 20168 39910 20224
rect 39670 19352 39726 19408
rect 39854 19352 39910 19408
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 40682 23432 40738 23488
rect 40682 23180 40738 23216
rect 40682 23160 40684 23180
rect 40684 23160 40736 23180
rect 40736 23160 40738 23180
rect 40498 21800 40554 21856
rect 40498 21392 40554 21448
rect 41234 24792 41290 24848
rect 40866 22924 40868 22944
rect 40868 22924 40920 22944
rect 40920 22924 40922 22944
rect 40866 22888 40922 22924
rect 40866 21936 40922 21992
rect 41418 22752 41474 22808
rect 40314 18264 40370 18320
rect 40222 17856 40278 17912
rect 42430 23468 42432 23488
rect 42432 23468 42484 23488
rect 42484 23468 42486 23488
rect 42430 23432 42486 23468
rect 42430 23160 42486 23216
rect 41878 22380 41880 22400
rect 41880 22380 41932 22400
rect 41932 22380 41934 22400
rect 41878 22344 41934 22380
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42614 22636 42670 22672
rect 42614 22616 42616 22636
rect 42616 22616 42668 22636
rect 42668 22616 42670 22636
rect 41234 20848 41290 20904
rect 41234 19080 41290 19136
rect 41142 18128 41198 18184
rect 39302 15408 39358 15464
rect 41602 21120 41658 21176
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42982 22072 43038 22128
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 43534 21800 43590 21856
rect 43442 21528 43498 21584
rect 41510 20032 41566 20088
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 43718 23704 43774 23760
rect 43994 23180 44050 23216
rect 43994 23160 43996 23180
rect 43996 23160 44048 23180
rect 44048 23160 44050 23180
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 41970 17720 42026 17776
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42706 17176 42762 17232
rect 44454 22616 44510 22672
rect 45558 22500 45614 22536
rect 45558 22480 45560 22500
rect 45560 22480 45612 22500
rect 45612 22480 45614 22500
rect 46110 23468 46112 23488
rect 46112 23468 46164 23488
rect 46164 23468 46166 23488
rect 46110 23432 46166 23468
rect 47030 24248 47086 24304
rect 46846 23024 46902 23080
rect 47122 23568 47178 23624
rect 47490 25064 47546 25120
rect 47582 24656 47638 24712
rect 47582 23568 47638 23624
rect 47766 23568 47822 23624
rect 47582 23432 47638 23488
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 49054 25472 49110 25528
rect 49238 24248 49294 24304
rect 49146 24112 49202 24168
rect 48594 23044 48650 23080
rect 48594 23024 48596 23044
rect 48596 23024 48648 23044
rect 48648 23024 48650 23044
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 48226 22616 48282 22672
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 46938 20304 46994 20360
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 48502 19896 48558 19952
rect 48778 21836 48780 21856
rect 48780 21836 48832 21856
rect 48832 21836 48834 21856
rect 48778 21800 48834 21836
rect 48778 20168 48834 20224
rect 49422 22208 49478 22264
rect 49238 21428 49240 21448
rect 49240 21428 49292 21448
rect 49292 21428 49294 21448
rect 49238 21392 49294 21428
rect 49330 20984 49386 21040
rect 49330 20576 49386 20632
rect 49422 19760 49478 19816
rect 48870 19352 48926 19408
rect 49330 19352 49386 19408
rect 49146 19216 49202 19272
rect 49238 18944 49294 19000
rect 48594 18808 48650 18864
rect 44086 18672 44142 18728
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 48778 18536 48834 18592
rect 49422 18128 49478 18184
rect 49330 17720 49386 17776
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49054 17076 49056 17096
rect 49056 17076 49108 17096
rect 49108 17076 49110 17096
rect 49054 17040 49110 17076
rect 48778 16904 48834 16960
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 49330 17312 49386 17368
rect 49146 16632 49202 16688
rect 49146 16496 49202 16552
rect 49330 16496 49386 16552
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 49422 16088 49478 16144
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 49146 15972 49202 16008
rect 49146 15952 49148 15972
rect 49148 15952 49200 15972
rect 49200 15952 49202 15972
rect 49330 15680 49386 15736
rect 41326 15544 41382 15600
rect 49330 15272 49386 15328
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 48870 15000 48926 15056
rect 49146 14884 49202 14920
rect 49146 14864 49148 14884
rect 49148 14864 49200 14884
rect 49200 14864 49202 14884
rect 49330 14864 49386 14920
rect 49054 14492 49056 14512
rect 49056 14492 49108 14512
rect 49108 14492 49110 14512
rect 49054 14456 49110 14492
rect 49238 14456 49294 14512
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 40038 12688 40094 12744
rect 49238 14048 49294 14104
rect 48226 13640 48282 13696
rect 49146 13268 49148 13288
rect 49148 13268 49200 13288
rect 49200 13268 49202 13288
rect 49146 13232 49202 13268
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 49146 12844 49202 12880
rect 49146 12824 49148 12844
rect 49148 12824 49200 12844
rect 49200 12824 49202 12844
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 40406 11756 40462 11792
rect 40406 11736 40408 11756
rect 40408 11736 40460 11756
rect 40460 11736 40462 11756
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 46846 7928 46902 7984
rect 49146 12416 49202 12472
rect 49146 12008 49202 12064
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 49146 11600 49202 11656
rect 49238 11192 49294 11248
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49146 10784 49202 10840
rect 49238 10376 49294 10432
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 49330 9968 49386 10024
rect 47306 9560 47362 9616
rect 49146 9152 49202 9208
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 46846 2624 46902 2680
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 49238 8744 49294 8800
rect 49330 8336 49386 8392
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7520 49202 7576
rect 49422 7112 49478 7168
rect 49238 6704 49294 6760
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 48686 6296 48742 6352
rect 49146 5888 49202 5944
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 49422 5480 49478 5536
rect 49330 5072 49386 5128
rect 48318 4664 48374 4720
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 4256 49202 4312
rect 46754 1808 46810 1864
rect 46662 1400 46718 1456
rect 49238 3848 49294 3904
rect 49146 3440 49202 3496
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 48686 3032 48742 3088
rect 48502 2216 48558 2272
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3141 25666 3207 25669
rect 0 25664 3207 25666
rect 0 25608 3146 25664
rect 3202 25608 3207 25664
rect 0 25606 3207 25608
rect 0 25576 800 25606
rect 3141 25603 3207 25606
rect 49049 25530 49115 25533
rect 50200 25530 51000 25560
rect 49049 25528 51000 25530
rect 49049 25472 49054 25528
rect 49110 25472 51000 25528
rect 49049 25470 51000 25472
rect 49049 25467 49115 25470
rect 50200 25440 51000 25470
rect 0 25258 800 25288
rect 3785 25258 3851 25261
rect 0 25256 3851 25258
rect 0 25200 3790 25256
rect 3846 25200 3851 25256
rect 0 25198 3851 25200
rect 0 25168 800 25198
rect 3785 25195 3851 25198
rect 47485 25122 47551 25125
rect 50200 25122 51000 25152
rect 47485 25120 51000 25122
rect 47485 25064 47490 25120
rect 47546 25064 51000 25120
rect 47485 25062 51000 25064
rect 47485 25059 47551 25062
rect 50200 25032 51000 25062
rect 0 24850 800 24880
rect 3877 24850 3943 24853
rect 0 24848 3943 24850
rect 0 24792 3882 24848
rect 3938 24792 3943 24848
rect 0 24790 3943 24792
rect 0 24760 800 24790
rect 3877 24787 3943 24790
rect 32489 24850 32555 24853
rect 41229 24850 41295 24853
rect 32489 24848 41295 24850
rect 32489 24792 32494 24848
rect 32550 24792 41234 24848
rect 41290 24792 41295 24848
rect 32489 24790 41295 24792
rect 32489 24787 32555 24790
rect 41229 24787 41295 24790
rect 33777 24714 33843 24717
rect 40033 24714 40099 24717
rect 33777 24712 40099 24714
rect 33777 24656 33782 24712
rect 33838 24656 40038 24712
rect 40094 24656 40099 24712
rect 33777 24654 40099 24656
rect 33777 24651 33843 24654
rect 40033 24651 40099 24654
rect 47577 24714 47643 24717
rect 50200 24714 51000 24744
rect 47577 24712 51000 24714
rect 47577 24656 47582 24712
rect 47638 24656 51000 24712
rect 47577 24654 51000 24656
rect 47577 24651 47643 24654
rect 50200 24624 51000 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 36905 24442 36971 24445
rect 36905 24440 41430 24442
rect 36905 24384 36910 24440
rect 36966 24384 41430 24440
rect 36905 24382 41430 24384
rect 36905 24379 36971 24382
rect 7465 24306 7531 24309
rect 25773 24306 25839 24309
rect 7465 24304 25839 24306
rect 7465 24248 7470 24304
rect 7526 24248 25778 24304
rect 25834 24248 25839 24304
rect 7465 24246 25839 24248
rect 7465 24243 7531 24246
rect 25773 24243 25839 24246
rect 31845 24306 31911 24309
rect 39389 24306 39455 24309
rect 31845 24304 39455 24306
rect 31845 24248 31850 24304
rect 31906 24248 39394 24304
rect 39450 24248 39455 24304
rect 31845 24246 39455 24248
rect 41370 24306 41430 24382
rect 47025 24306 47091 24309
rect 41370 24304 47091 24306
rect 41370 24248 47030 24304
rect 47086 24248 47091 24304
rect 41370 24246 47091 24248
rect 31845 24243 31911 24246
rect 39389 24243 39455 24246
rect 47025 24243 47091 24246
rect 49233 24306 49299 24309
rect 50200 24306 51000 24336
rect 49233 24304 51000 24306
rect 49233 24248 49238 24304
rect 49294 24248 51000 24304
rect 49233 24246 51000 24248
rect 49233 24243 49299 24246
rect 50200 24216 51000 24246
rect 26601 24170 26667 24173
rect 49141 24170 49207 24173
rect 26601 24168 49207 24170
rect 26601 24112 26606 24168
rect 26662 24112 49146 24168
rect 49202 24112 49207 24168
rect 26601 24110 49207 24112
rect 26601 24107 26667 24110
rect 49141 24107 49207 24110
rect 0 24034 800 24064
rect 3509 24034 3575 24037
rect 0 24032 3575 24034
rect 0 23976 3514 24032
rect 3570 23976 3575 24032
rect 0 23974 3575 23976
rect 0 23944 800 23974
rect 3509 23971 3575 23974
rect 35433 24034 35499 24037
rect 37641 24034 37707 24037
rect 35433 24032 37707 24034
rect 35433 23976 35438 24032
rect 35494 23976 37646 24032
rect 37702 23976 37707 24032
rect 35433 23974 37707 23976
rect 35433 23971 35499 23974
rect 37641 23971 37707 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 29913 23898 29979 23901
rect 33593 23898 33659 23901
rect 50200 23898 51000 23928
rect 29913 23896 33659 23898
rect 29913 23840 29918 23896
rect 29974 23840 33598 23896
rect 33654 23840 33659 23896
rect 29913 23838 33659 23840
rect 29913 23835 29979 23838
rect 33593 23835 33659 23838
rect 48454 23838 51000 23898
rect 30005 23762 30071 23765
rect 31109 23762 31175 23765
rect 32949 23762 33015 23765
rect 30005 23760 33015 23762
rect 30005 23704 30010 23760
rect 30066 23704 31114 23760
rect 31170 23704 32954 23760
rect 33010 23704 33015 23760
rect 30005 23702 33015 23704
rect 30005 23699 30071 23702
rect 31109 23699 31175 23702
rect 32949 23699 33015 23702
rect 34789 23762 34855 23765
rect 43713 23762 43779 23765
rect 34789 23760 43779 23762
rect 34789 23704 34794 23760
rect 34850 23704 43718 23760
rect 43774 23704 43779 23760
rect 34789 23702 43779 23704
rect 34789 23699 34855 23702
rect 43713 23699 43779 23702
rect 0 23626 800 23656
rect 3969 23626 4035 23629
rect 0 23624 4035 23626
rect 0 23568 3974 23624
rect 4030 23568 4035 23624
rect 0 23566 4035 23568
rect 0 23536 800 23566
rect 3969 23563 4035 23566
rect 31661 23626 31727 23629
rect 36077 23626 36143 23629
rect 31661 23624 36143 23626
rect 31661 23568 31666 23624
rect 31722 23568 36082 23624
rect 36138 23568 36143 23624
rect 31661 23566 36143 23568
rect 31661 23563 31727 23566
rect 36077 23563 36143 23566
rect 47117 23626 47183 23629
rect 47577 23626 47643 23629
rect 47117 23624 47643 23626
rect 47117 23568 47122 23624
rect 47178 23568 47582 23624
rect 47638 23568 47643 23624
rect 47117 23566 47643 23568
rect 47117 23563 47183 23566
rect 47577 23563 47643 23566
rect 47761 23626 47827 23629
rect 48454 23626 48514 23838
rect 50200 23808 51000 23838
rect 47761 23624 48514 23626
rect 47761 23568 47766 23624
rect 47822 23568 48514 23624
rect 47761 23566 48514 23568
rect 47761 23563 47827 23566
rect 35065 23490 35131 23493
rect 40677 23490 40743 23493
rect 42425 23490 42491 23493
rect 46105 23492 46171 23493
rect 46054 23490 46060 23492
rect 35065 23488 40743 23490
rect 35065 23432 35070 23488
rect 35126 23432 40682 23488
rect 40738 23432 40743 23488
rect 35065 23430 40743 23432
rect 35065 23427 35131 23430
rect 40677 23427 40743 23430
rect 41370 23488 42491 23490
rect 41370 23432 42430 23488
rect 42486 23432 42491 23488
rect 41370 23430 42491 23432
rect 46014 23430 46060 23490
rect 46124 23488 46171 23492
rect 46166 23432 46171 23488
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 38653 23354 38719 23357
rect 39757 23354 39823 23357
rect 41370 23354 41430 23430
rect 42425 23427 42491 23430
rect 46054 23428 46060 23430
rect 46124 23428 46171 23432
rect 46105 23427 46171 23428
rect 47577 23490 47643 23493
rect 50200 23490 51000 23520
rect 47577 23488 51000 23490
rect 47577 23432 47582 23488
rect 47638 23432 51000 23488
rect 47577 23430 51000 23432
rect 47577 23427 47643 23430
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 50200 23400 51000 23430
rect 42946 23359 43262 23360
rect 38653 23352 41430 23354
rect 38653 23296 38658 23352
rect 38714 23296 39762 23352
rect 39818 23296 41430 23352
rect 38653 23294 41430 23296
rect 38653 23291 38719 23294
rect 39757 23291 39823 23294
rect 0 23218 800 23248
rect 2957 23218 3023 23221
rect 0 23216 3023 23218
rect 0 23160 2962 23216
rect 3018 23160 3023 23216
rect 0 23158 3023 23160
rect 0 23128 800 23158
rect 2957 23155 3023 23158
rect 33225 23218 33291 23221
rect 38837 23218 38903 23221
rect 33225 23216 38903 23218
rect 33225 23160 33230 23216
rect 33286 23160 38842 23216
rect 38898 23160 38903 23216
rect 33225 23158 38903 23160
rect 33225 23155 33291 23158
rect 38837 23155 38903 23158
rect 39021 23218 39087 23221
rect 40677 23218 40743 23221
rect 39021 23216 40743 23218
rect 39021 23160 39026 23216
rect 39082 23160 40682 23216
rect 40738 23160 40743 23216
rect 39021 23158 40743 23160
rect 39021 23155 39087 23158
rect 40677 23155 40743 23158
rect 42425 23218 42491 23221
rect 43989 23218 44055 23221
rect 42425 23216 44055 23218
rect 42425 23160 42430 23216
rect 42486 23160 43994 23216
rect 44050 23160 44055 23216
rect 42425 23158 44055 23160
rect 42425 23155 42491 23158
rect 43989 23155 44055 23158
rect 11329 23082 11395 23085
rect 23289 23082 23355 23085
rect 11329 23080 23355 23082
rect 11329 23024 11334 23080
rect 11390 23024 23294 23080
rect 23350 23024 23355 23080
rect 11329 23022 23355 23024
rect 11329 23019 11395 23022
rect 23289 23019 23355 23022
rect 35157 23082 35223 23085
rect 39297 23082 39363 23085
rect 35157 23080 39363 23082
rect 35157 23024 35162 23080
rect 35218 23024 39302 23080
rect 39358 23024 39363 23080
rect 35157 23022 39363 23024
rect 35157 23019 35223 23022
rect 39297 23019 39363 23022
rect 39573 23082 39639 23085
rect 46841 23082 46907 23085
rect 39573 23080 46907 23082
rect 39573 23024 39578 23080
rect 39634 23024 46846 23080
rect 46902 23024 46907 23080
rect 39573 23022 46907 23024
rect 39573 23019 39639 23022
rect 46841 23019 46907 23022
rect 48589 23082 48655 23085
rect 50200 23082 51000 23112
rect 48589 23080 51000 23082
rect 48589 23024 48594 23080
rect 48650 23024 51000 23080
rect 48589 23022 51000 23024
rect 48589 23019 48655 23022
rect 50200 22992 51000 23022
rect 25313 22948 25379 22949
rect 25262 22884 25268 22948
rect 25332 22946 25379 22948
rect 39113 22946 39179 22949
rect 40861 22946 40927 22949
rect 25332 22944 25424 22946
rect 25374 22888 25424 22944
rect 25332 22886 25424 22888
rect 39113 22944 40927 22946
rect 39113 22888 39118 22944
rect 39174 22888 40866 22944
rect 40922 22888 40927 22944
rect 39113 22886 40927 22888
rect 25332 22884 25379 22886
rect 25313 22883 25379 22884
rect 39113 22883 39179 22886
rect 40861 22883 40927 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 3969 22810 4035 22813
rect 0 22808 4035 22810
rect 0 22752 3974 22808
rect 4030 22752 4035 22808
rect 0 22750 4035 22752
rect 0 22720 800 22750
rect 3969 22747 4035 22750
rect 40033 22810 40099 22813
rect 41413 22810 41479 22813
rect 40033 22808 41479 22810
rect 40033 22752 40038 22808
rect 40094 22752 41418 22808
rect 41474 22752 41479 22808
rect 40033 22750 41479 22752
rect 40033 22747 40099 22750
rect 41413 22747 41479 22750
rect 19793 22674 19859 22677
rect 29637 22674 29703 22677
rect 19793 22672 29703 22674
rect 19793 22616 19798 22672
rect 19854 22616 29642 22672
rect 29698 22616 29703 22672
rect 19793 22614 29703 22616
rect 19793 22611 19859 22614
rect 29637 22611 29703 22614
rect 30649 22674 30715 22677
rect 34789 22674 34855 22677
rect 30649 22672 34855 22674
rect 30649 22616 30654 22672
rect 30710 22616 34794 22672
rect 34850 22616 34855 22672
rect 30649 22614 34855 22616
rect 30649 22611 30715 22614
rect 34789 22611 34855 22614
rect 35709 22674 35775 22677
rect 42609 22674 42675 22677
rect 44449 22674 44515 22677
rect 35709 22672 44515 22674
rect 35709 22616 35714 22672
rect 35770 22616 42614 22672
rect 42670 22616 44454 22672
rect 44510 22616 44515 22672
rect 35709 22614 44515 22616
rect 35709 22611 35775 22614
rect 42609 22611 42675 22614
rect 44449 22611 44515 22614
rect 48221 22674 48287 22677
rect 50200 22674 51000 22704
rect 48221 22672 51000 22674
rect 48221 22616 48226 22672
rect 48282 22616 51000 22672
rect 48221 22614 51000 22616
rect 48221 22611 48287 22614
rect 50200 22584 51000 22614
rect 24761 22538 24827 22541
rect 31477 22538 31543 22541
rect 24761 22536 31543 22538
rect 24761 22480 24766 22536
rect 24822 22480 31482 22536
rect 31538 22480 31543 22536
rect 24761 22478 31543 22480
rect 24761 22475 24827 22478
rect 31477 22475 31543 22478
rect 37457 22538 37523 22541
rect 45553 22538 45619 22541
rect 37457 22536 45619 22538
rect 37457 22480 37462 22536
rect 37518 22480 45558 22536
rect 45614 22480 45619 22536
rect 37457 22478 45619 22480
rect 37457 22475 37523 22478
rect 45553 22475 45619 22478
rect 0 22402 800 22432
rect 25129 22402 25195 22405
rect 29729 22402 29795 22405
rect 0 22342 2146 22402
rect 0 22312 800 22342
rect 2086 22130 2146 22342
rect 25129 22400 29795 22402
rect 25129 22344 25134 22400
rect 25190 22344 29734 22400
rect 29790 22344 29795 22400
rect 25129 22342 29795 22344
rect 25129 22339 25195 22342
rect 29729 22339 29795 22342
rect 33409 22402 33475 22405
rect 35341 22402 35407 22405
rect 41873 22402 41939 22405
rect 33409 22400 41939 22402
rect 33409 22344 33414 22400
rect 33470 22344 35346 22400
rect 35402 22344 41878 22400
rect 41934 22344 41939 22400
rect 33409 22342 41939 22344
rect 33409 22339 33475 22342
rect 35341 22339 35407 22342
rect 41873 22339 41939 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 23749 22266 23815 22269
rect 28257 22266 28323 22269
rect 23749 22264 28323 22266
rect 23749 22208 23754 22264
rect 23810 22208 28262 22264
rect 28318 22208 28323 22264
rect 23749 22206 28323 22208
rect 23749 22203 23815 22206
rect 28257 22203 28323 22206
rect 37089 22266 37155 22269
rect 49417 22266 49483 22269
rect 50200 22266 51000 22296
rect 37089 22264 41430 22266
rect 37089 22208 37094 22264
rect 37150 22208 41430 22264
rect 37089 22206 41430 22208
rect 37089 22203 37155 22206
rect 4153 22130 4219 22133
rect 2086 22128 4219 22130
rect 2086 22072 4158 22128
rect 4214 22072 4219 22128
rect 2086 22070 4219 22072
rect 4153 22067 4219 22070
rect 21081 22130 21147 22133
rect 24209 22130 24275 22133
rect 21081 22128 24275 22130
rect 21081 22072 21086 22128
rect 21142 22072 24214 22128
rect 24270 22072 24275 22128
rect 21081 22070 24275 22072
rect 21081 22067 21147 22070
rect 24209 22067 24275 22070
rect 24853 22130 24919 22133
rect 26601 22130 26667 22133
rect 24853 22128 26667 22130
rect 24853 22072 24858 22128
rect 24914 22072 26606 22128
rect 26662 22072 26667 22128
rect 24853 22070 26667 22072
rect 24853 22067 24919 22070
rect 26601 22067 26667 22070
rect 32121 22130 32187 22133
rect 34881 22130 34947 22133
rect 32121 22128 34947 22130
rect 32121 22072 32126 22128
rect 32182 22072 34886 22128
rect 34942 22072 34947 22128
rect 32121 22070 34947 22072
rect 41370 22130 41430 22206
rect 49417 22264 51000 22266
rect 49417 22208 49422 22264
rect 49478 22208 51000 22264
rect 49417 22206 51000 22208
rect 49417 22203 49483 22206
rect 50200 22176 51000 22206
rect 42977 22130 43043 22133
rect 41370 22128 43043 22130
rect 41370 22072 42982 22128
rect 43038 22072 43043 22128
rect 41370 22070 43043 22072
rect 32121 22067 32187 22070
rect 34881 22067 34947 22070
rect 42977 22067 43043 22070
rect 0 21994 800 22024
rect 3233 21994 3299 21997
rect 0 21992 3299 21994
rect 0 21936 3238 21992
rect 3294 21936 3299 21992
rect 0 21934 3299 21936
rect 0 21904 800 21934
rect 3233 21931 3299 21934
rect 11697 21994 11763 21997
rect 18689 21994 18755 21997
rect 24853 21994 24919 21997
rect 25773 21994 25839 21997
rect 11697 21992 25839 21994
rect 11697 21936 11702 21992
rect 11758 21936 18694 21992
rect 18750 21936 24858 21992
rect 24914 21936 25778 21992
rect 25834 21936 25839 21992
rect 11697 21934 25839 21936
rect 11697 21931 11763 21934
rect 18689 21931 18755 21934
rect 24853 21931 24919 21934
rect 25773 21931 25839 21934
rect 27613 21994 27679 21997
rect 30189 21994 30255 21997
rect 27613 21992 30255 21994
rect 27613 21936 27618 21992
rect 27674 21936 30194 21992
rect 30250 21936 30255 21992
rect 27613 21934 30255 21936
rect 27613 21931 27679 21934
rect 30189 21931 30255 21934
rect 34421 21994 34487 21997
rect 40861 21994 40927 21997
rect 34421 21992 40927 21994
rect 34421 21936 34426 21992
rect 34482 21936 40866 21992
rect 40922 21936 40927 21992
rect 34421 21934 40927 21936
rect 34421 21931 34487 21934
rect 40861 21931 40927 21934
rect 40493 21858 40559 21861
rect 43529 21858 43595 21861
rect 40493 21856 43595 21858
rect 40493 21800 40498 21856
rect 40554 21800 43534 21856
rect 43590 21800 43595 21856
rect 40493 21798 43595 21800
rect 40493 21795 40559 21798
rect 43529 21795 43595 21798
rect 48773 21858 48839 21861
rect 50200 21858 51000 21888
rect 48773 21856 51000 21858
rect 48773 21800 48778 21856
rect 48834 21800 51000 21856
rect 48773 21798 51000 21800
rect 48773 21795 48839 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 50200 21768 51000 21798
rect 47946 21727 48262 21728
rect 29913 21722 29979 21725
rect 35985 21722 36051 21725
rect 29913 21720 36051 21722
rect 29913 21664 29918 21720
rect 29974 21664 35990 21720
rect 36046 21664 36051 21720
rect 29913 21662 36051 21664
rect 29913 21659 29979 21662
rect 35985 21659 36051 21662
rect 0 21586 800 21616
rect 1761 21586 1827 21589
rect 0 21584 1827 21586
rect 0 21528 1766 21584
rect 1822 21528 1827 21584
rect 0 21526 1827 21528
rect 0 21496 800 21526
rect 1761 21523 1827 21526
rect 6545 21586 6611 21589
rect 9581 21586 9647 21589
rect 6545 21584 9647 21586
rect 6545 21528 6550 21584
rect 6606 21528 9586 21584
rect 9642 21528 9647 21584
rect 6545 21526 9647 21528
rect 6545 21523 6611 21526
rect 9581 21523 9647 21526
rect 15469 21586 15535 21589
rect 28809 21586 28875 21589
rect 30373 21588 30439 21589
rect 30373 21586 30420 21588
rect 15469 21584 30420 21586
rect 30484 21586 30490 21588
rect 31201 21586 31267 21589
rect 33501 21586 33567 21589
rect 43437 21586 43503 21589
rect 15469 21528 15474 21584
rect 15530 21528 28814 21584
rect 28870 21528 30378 21584
rect 15469 21526 30420 21528
rect 15469 21523 15535 21526
rect 28809 21523 28875 21526
rect 30373 21524 30420 21526
rect 30484 21526 30566 21586
rect 31201 21584 43503 21586
rect 31201 21528 31206 21584
rect 31262 21528 33506 21584
rect 33562 21528 43442 21584
rect 43498 21528 43503 21584
rect 31201 21526 43503 21528
rect 30484 21524 30490 21526
rect 30373 21523 30439 21524
rect 31201 21523 31267 21526
rect 33501 21523 33567 21526
rect 43437 21523 43503 21526
rect 21357 21450 21423 21453
rect 26417 21450 26483 21453
rect 21357 21448 26483 21450
rect 21357 21392 21362 21448
rect 21418 21392 26422 21448
rect 26478 21392 26483 21448
rect 21357 21390 26483 21392
rect 21357 21387 21423 21390
rect 26417 21387 26483 21390
rect 37273 21450 37339 21453
rect 40493 21450 40559 21453
rect 37273 21448 40559 21450
rect 37273 21392 37278 21448
rect 37334 21392 40498 21448
rect 40554 21392 40559 21448
rect 37273 21390 40559 21392
rect 37273 21387 37339 21390
rect 40493 21387 40559 21390
rect 49233 21450 49299 21453
rect 50200 21450 51000 21480
rect 49233 21448 51000 21450
rect 49233 21392 49238 21448
rect 49294 21392 51000 21448
rect 49233 21390 51000 21392
rect 49233 21387 49299 21390
rect 50200 21360 51000 21390
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 38285 21178 38351 21181
rect 41597 21178 41663 21181
rect 38285 21176 41663 21178
rect 38285 21120 38290 21176
rect 38346 21120 41602 21176
rect 41658 21120 41663 21176
rect 38285 21118 41663 21120
rect 38285 21115 38351 21118
rect 41597 21115 41663 21118
rect 12801 21042 12867 21045
rect 21265 21042 21331 21045
rect 25129 21042 25195 21045
rect 12801 21040 25195 21042
rect 12801 20984 12806 21040
rect 12862 20984 21270 21040
rect 21326 20984 25134 21040
rect 25190 20984 25195 21040
rect 12801 20982 25195 20984
rect 12801 20979 12867 20982
rect 21265 20979 21331 20982
rect 25129 20979 25195 20982
rect 25773 21042 25839 21045
rect 30005 21042 30071 21045
rect 25773 21040 30071 21042
rect 25773 20984 25778 21040
rect 25834 20984 30010 21040
rect 30066 20984 30071 21040
rect 25773 20982 30071 20984
rect 25773 20979 25839 20982
rect 30005 20979 30071 20982
rect 31109 21042 31175 21045
rect 31661 21042 31727 21045
rect 38745 21042 38811 21045
rect 31109 21040 38811 21042
rect 31109 20984 31114 21040
rect 31170 20984 31666 21040
rect 31722 20984 38750 21040
rect 38806 20984 38811 21040
rect 31109 20982 38811 20984
rect 31109 20979 31175 20982
rect 31661 20979 31727 20982
rect 38745 20979 38811 20982
rect 49325 21042 49391 21045
rect 50200 21042 51000 21072
rect 49325 21040 51000 21042
rect 49325 20984 49330 21040
rect 49386 20984 51000 21040
rect 49325 20982 51000 20984
rect 49325 20979 49391 20982
rect 50200 20952 51000 20982
rect 8385 20906 8451 20909
rect 23749 20906 23815 20909
rect 8385 20904 23815 20906
rect 8385 20848 8390 20904
rect 8446 20848 23754 20904
rect 23810 20848 23815 20904
rect 8385 20846 23815 20848
rect 8385 20843 8451 20846
rect 23749 20843 23815 20846
rect 27429 20906 27495 20909
rect 29821 20906 29887 20909
rect 27429 20904 29887 20906
rect 27429 20848 27434 20904
rect 27490 20848 29826 20904
rect 29882 20848 29887 20904
rect 27429 20846 29887 20848
rect 27429 20843 27495 20846
rect 29821 20843 29887 20846
rect 31753 20906 31819 20909
rect 32581 20906 32647 20909
rect 41229 20906 41295 20909
rect 31753 20904 41295 20906
rect 31753 20848 31758 20904
rect 31814 20848 32586 20904
rect 32642 20848 41234 20904
rect 41290 20848 41295 20904
rect 31753 20846 41295 20848
rect 31753 20843 31819 20846
rect 32581 20843 32647 20846
rect 41229 20843 41295 20846
rect 0 20770 800 20800
rect 1025 20770 1091 20773
rect 0 20768 1091 20770
rect 0 20712 1030 20768
rect 1086 20712 1091 20768
rect 0 20710 1091 20712
rect 0 20680 800 20710
rect 1025 20707 1091 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 21541 20634 21607 20637
rect 25405 20634 25471 20637
rect 21541 20632 25471 20634
rect 21541 20576 21546 20632
rect 21602 20576 25410 20632
rect 25466 20576 25471 20632
rect 21541 20574 25471 20576
rect 21541 20571 21607 20574
rect 25405 20571 25471 20574
rect 35065 20634 35131 20637
rect 35525 20634 35591 20637
rect 36721 20634 36787 20637
rect 35065 20632 36787 20634
rect 35065 20576 35070 20632
rect 35126 20576 35530 20632
rect 35586 20576 36726 20632
rect 36782 20576 36787 20632
rect 35065 20574 36787 20576
rect 35065 20571 35131 20574
rect 35525 20571 35591 20574
rect 36721 20571 36787 20574
rect 49325 20634 49391 20637
rect 50200 20634 51000 20664
rect 49325 20632 51000 20634
rect 49325 20576 49330 20632
rect 49386 20576 51000 20632
rect 49325 20574 51000 20576
rect 49325 20571 49391 20574
rect 50200 20544 51000 20574
rect 9857 20498 9923 20501
rect 17401 20498 17467 20501
rect 9857 20496 17467 20498
rect 9857 20440 9862 20496
rect 9918 20440 17406 20496
rect 17462 20440 17467 20496
rect 9857 20438 17467 20440
rect 9857 20435 9923 20438
rect 17401 20435 17467 20438
rect 17861 20498 17927 20501
rect 35249 20498 35315 20501
rect 17861 20496 35315 20498
rect 17861 20440 17866 20496
rect 17922 20440 35254 20496
rect 35310 20440 35315 20496
rect 17861 20438 35315 20440
rect 17861 20435 17927 20438
rect 35249 20435 35315 20438
rect 0 20362 800 20392
rect 1301 20362 1367 20365
rect 0 20360 1367 20362
rect 0 20304 1306 20360
rect 1362 20304 1367 20360
rect 0 20302 1367 20304
rect 0 20272 800 20302
rect 1301 20299 1367 20302
rect 10777 20362 10843 20365
rect 14917 20362 14983 20365
rect 10777 20360 14983 20362
rect 10777 20304 10782 20360
rect 10838 20304 14922 20360
rect 14978 20304 14983 20360
rect 10777 20302 14983 20304
rect 10777 20299 10843 20302
rect 14917 20299 14983 20302
rect 15285 20362 15351 20365
rect 26049 20362 26115 20365
rect 31937 20362 32003 20365
rect 46933 20362 46999 20365
rect 15285 20360 26115 20362
rect 15285 20304 15290 20360
rect 15346 20304 26054 20360
rect 26110 20304 26115 20360
rect 15285 20302 26115 20304
rect 15285 20299 15351 20302
rect 26049 20299 26115 20302
rect 31710 20360 46999 20362
rect 31710 20304 31942 20360
rect 31998 20304 46938 20360
rect 46994 20304 46999 20360
rect 31710 20302 46999 20304
rect 25313 20226 25379 20229
rect 31710 20226 31770 20302
rect 31937 20299 32003 20302
rect 46933 20299 46999 20302
rect 25313 20224 31770 20226
rect 25313 20168 25318 20224
rect 25374 20168 31770 20224
rect 25313 20166 31770 20168
rect 34513 20226 34579 20229
rect 39849 20226 39915 20229
rect 34513 20224 39915 20226
rect 34513 20168 34518 20224
rect 34574 20168 39854 20224
rect 39910 20168 39915 20224
rect 34513 20166 39915 20168
rect 25313 20163 25379 20166
rect 34513 20163 34579 20166
rect 39849 20163 39915 20166
rect 48773 20226 48839 20229
rect 50200 20226 51000 20256
rect 48773 20224 51000 20226
rect 48773 20168 48778 20224
rect 48834 20168 51000 20224
rect 48773 20166 51000 20168
rect 48773 20163 48839 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 50200 20136 51000 20166
rect 42946 20095 43262 20096
rect 36629 20090 36695 20093
rect 41505 20090 41571 20093
rect 36629 20088 41571 20090
rect 36629 20032 36634 20088
rect 36690 20032 41510 20088
rect 41566 20032 41571 20088
rect 36629 20030 41571 20032
rect 36629 20027 36695 20030
rect 41505 20027 41571 20030
rect 0 19954 800 19984
rect 1761 19954 1827 19957
rect 0 19952 1827 19954
rect 0 19896 1766 19952
rect 1822 19896 1827 19952
rect 0 19894 1827 19896
rect 0 19864 800 19894
rect 1761 19891 1827 19894
rect 13629 19954 13695 19957
rect 23013 19954 23079 19957
rect 23841 19954 23907 19957
rect 28441 19954 28507 19957
rect 48497 19954 48563 19957
rect 13629 19952 48563 19954
rect 13629 19896 13634 19952
rect 13690 19896 23018 19952
rect 23074 19896 23846 19952
rect 23902 19896 28446 19952
rect 28502 19896 48502 19952
rect 48558 19896 48563 19952
rect 13629 19894 48563 19896
rect 13629 19891 13695 19894
rect 23013 19891 23079 19894
rect 23841 19891 23907 19894
rect 28441 19891 28507 19894
rect 48497 19891 48563 19894
rect 13813 19818 13879 19821
rect 25129 19818 25195 19821
rect 13813 19816 25195 19818
rect 13813 19760 13818 19816
rect 13874 19760 25134 19816
rect 25190 19760 25195 19816
rect 13813 19758 25195 19760
rect 13813 19755 13879 19758
rect 25129 19755 25195 19758
rect 30414 19756 30420 19820
rect 30484 19818 30490 19820
rect 38193 19818 38259 19821
rect 30484 19816 38259 19818
rect 30484 19760 38198 19816
rect 38254 19760 38259 19816
rect 30484 19758 38259 19760
rect 30484 19756 30490 19758
rect 38193 19755 38259 19758
rect 49417 19818 49483 19821
rect 50200 19818 51000 19848
rect 49417 19816 51000 19818
rect 49417 19760 49422 19816
rect 49478 19760 51000 19816
rect 49417 19758 51000 19760
rect 49417 19755 49483 19758
rect 50200 19728 51000 19758
rect 11881 19682 11947 19685
rect 15837 19682 15903 19685
rect 11881 19680 15903 19682
rect 11881 19624 11886 19680
rect 11942 19624 15842 19680
rect 15898 19624 15903 19680
rect 11881 19622 15903 19624
rect 11881 19619 11947 19622
rect 15837 19619 15903 19622
rect 30373 19682 30439 19685
rect 30373 19680 37842 19682
rect 30373 19624 30378 19680
rect 30434 19624 37842 19680
rect 30373 19622 37842 19624
rect 30373 19619 30439 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 2865 19546 2931 19549
rect 0 19544 2931 19546
rect 0 19488 2870 19544
rect 2926 19488 2931 19544
rect 0 19486 2931 19488
rect 0 19456 800 19486
rect 2865 19483 2931 19486
rect 14273 19546 14339 19549
rect 16430 19546 16436 19548
rect 14273 19544 16436 19546
rect 14273 19488 14278 19544
rect 14334 19488 16436 19544
rect 14273 19486 16436 19488
rect 14273 19483 14339 19486
rect 16430 19484 16436 19486
rect 16500 19484 16506 19548
rect 29637 19546 29703 19549
rect 36629 19546 36695 19549
rect 29637 19544 36695 19546
rect 29637 19488 29642 19544
rect 29698 19488 36634 19544
rect 36690 19488 36695 19544
rect 29637 19486 36695 19488
rect 29637 19483 29703 19486
rect 36629 19483 36695 19486
rect 9949 19410 10015 19413
rect 13721 19410 13787 19413
rect 9949 19408 13787 19410
rect 9949 19352 9954 19408
rect 10010 19352 13726 19408
rect 13782 19352 13787 19408
rect 9949 19350 13787 19352
rect 9949 19347 10015 19350
rect 13721 19347 13787 19350
rect 15193 19410 15259 19413
rect 16205 19410 16271 19413
rect 30097 19410 30163 19413
rect 30925 19410 30991 19413
rect 15193 19408 30991 19410
rect 15193 19352 15198 19408
rect 15254 19352 16210 19408
rect 16266 19352 30102 19408
rect 30158 19352 30930 19408
rect 30986 19352 30991 19408
rect 15193 19350 30991 19352
rect 37782 19410 37842 19622
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 39665 19410 39731 19413
rect 37782 19408 39731 19410
rect 37782 19352 39670 19408
rect 39726 19352 39731 19408
rect 37782 19350 39731 19352
rect 15193 19347 15259 19350
rect 16205 19347 16271 19350
rect 30097 19347 30163 19350
rect 30925 19347 30991 19350
rect 39665 19347 39731 19350
rect 39849 19410 39915 19413
rect 48865 19410 48931 19413
rect 39849 19408 48931 19410
rect 39849 19352 39854 19408
rect 39910 19352 48870 19408
rect 48926 19352 48931 19408
rect 39849 19350 48931 19352
rect 39849 19347 39915 19350
rect 48865 19347 48931 19350
rect 49325 19410 49391 19413
rect 50200 19410 51000 19440
rect 49325 19408 51000 19410
rect 49325 19352 49330 19408
rect 49386 19352 51000 19408
rect 49325 19350 51000 19352
rect 49325 19347 49391 19350
rect 50200 19320 51000 19350
rect 11053 19274 11119 19277
rect 15561 19274 15627 19277
rect 11053 19272 15627 19274
rect 11053 19216 11058 19272
rect 11114 19216 15566 19272
rect 15622 19216 15627 19272
rect 11053 19214 15627 19216
rect 11053 19211 11119 19214
rect 15561 19211 15627 19214
rect 29913 19274 29979 19277
rect 38009 19274 38075 19277
rect 49141 19274 49207 19277
rect 29913 19272 38075 19274
rect 29913 19216 29918 19272
rect 29974 19216 38014 19272
rect 38070 19216 38075 19272
rect 29913 19214 38075 19216
rect 29913 19211 29979 19214
rect 38009 19211 38075 19214
rect 41370 19272 49207 19274
rect 41370 19216 49146 19272
rect 49202 19216 49207 19272
rect 41370 19214 49207 19216
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 25037 19138 25103 19141
rect 28533 19138 28599 19141
rect 25037 19136 28599 19138
rect 25037 19080 25042 19136
rect 25098 19080 28538 19136
rect 28594 19080 28599 19136
rect 25037 19078 28599 19080
rect 25037 19075 25103 19078
rect 28533 19075 28599 19078
rect 30097 19138 30163 19141
rect 31477 19138 31543 19141
rect 41229 19138 41295 19141
rect 41370 19138 41430 19214
rect 49141 19211 49207 19214
rect 30097 19136 31543 19138
rect 30097 19080 30102 19136
rect 30158 19080 31482 19136
rect 31538 19080 31543 19136
rect 30097 19078 31543 19080
rect 30097 19075 30163 19078
rect 31477 19075 31543 19078
rect 34102 19136 41430 19138
rect 34102 19080 41234 19136
rect 41290 19080 41430 19136
rect 34102 19078 41430 19080
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 27705 19002 27771 19005
rect 28625 19002 28691 19005
rect 27705 19000 28691 19002
rect 27705 18944 27710 19000
rect 27766 18944 28630 19000
rect 28686 18944 28691 19000
rect 27705 18942 28691 18944
rect 27705 18939 27771 18942
rect 28625 18939 28691 18942
rect 5349 18866 5415 18869
rect 11237 18866 11303 18869
rect 5349 18864 11303 18866
rect 5349 18808 5354 18864
rect 5410 18808 11242 18864
rect 11298 18808 11303 18864
rect 5349 18806 11303 18808
rect 5349 18803 5415 18806
rect 11237 18803 11303 18806
rect 12157 18866 12223 18869
rect 18597 18866 18663 18869
rect 12157 18864 18663 18866
rect 12157 18808 12162 18864
rect 12218 18808 18602 18864
rect 18658 18808 18663 18864
rect 12157 18806 18663 18808
rect 12157 18803 12223 18806
rect 18597 18803 18663 18806
rect 20713 18866 20779 18869
rect 28993 18866 29059 18869
rect 20713 18864 29059 18866
rect 20713 18808 20718 18864
rect 20774 18808 28998 18864
rect 29054 18808 29059 18864
rect 20713 18806 29059 18808
rect 20713 18803 20779 18806
rect 28993 18803 29059 18806
rect 30005 18866 30071 18869
rect 32949 18866 33015 18869
rect 33593 18866 33659 18869
rect 30005 18864 33659 18866
rect 30005 18808 30010 18864
rect 30066 18808 32954 18864
rect 33010 18808 33598 18864
rect 33654 18808 33659 18864
rect 30005 18806 33659 18808
rect 30005 18803 30071 18806
rect 32949 18803 33015 18806
rect 33593 18803 33659 18806
rect 0 18730 800 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 800 18670
rect 1485 18667 1551 18670
rect 17401 18730 17467 18733
rect 19333 18730 19399 18733
rect 28349 18730 28415 18733
rect 17401 18728 28415 18730
rect 17401 18672 17406 18728
rect 17462 18672 19338 18728
rect 19394 18672 28354 18728
rect 28410 18672 28415 18728
rect 17401 18670 28415 18672
rect 17401 18667 17467 18670
rect 19333 18667 19399 18670
rect 28349 18667 28415 18670
rect 30925 18730 30991 18733
rect 34102 18730 34162 19078
rect 41229 19075 41295 19078
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 34973 19002 35039 19005
rect 35249 19002 35315 19005
rect 36905 19002 36971 19005
rect 37365 19002 37431 19005
rect 37641 19002 37707 19005
rect 34973 19000 37707 19002
rect 34973 18944 34978 19000
rect 35034 18944 35254 19000
rect 35310 18944 36910 19000
rect 36966 18944 37370 19000
rect 37426 18944 37646 19000
rect 37702 18944 37707 19000
rect 34973 18942 37707 18944
rect 34973 18939 35039 18942
rect 35249 18939 35315 18942
rect 36905 18939 36971 18942
rect 37365 18939 37431 18942
rect 37641 18939 37707 18942
rect 49233 19002 49299 19005
rect 50200 19002 51000 19032
rect 49233 19000 51000 19002
rect 49233 18944 49238 19000
rect 49294 18944 51000 19000
rect 49233 18942 51000 18944
rect 49233 18939 49299 18942
rect 50200 18912 51000 18942
rect 34237 18866 34303 18869
rect 48589 18866 48655 18869
rect 34237 18864 48655 18866
rect 34237 18808 34242 18864
rect 34298 18808 48594 18864
rect 48650 18808 48655 18864
rect 34237 18806 48655 18808
rect 34237 18803 34303 18806
rect 48589 18803 48655 18806
rect 44081 18730 44147 18733
rect 30925 18728 34162 18730
rect 30925 18672 30930 18728
rect 30986 18672 34162 18728
rect 30925 18670 34162 18672
rect 36494 18728 44147 18730
rect 36494 18672 44086 18728
rect 44142 18672 44147 18728
rect 36494 18670 44147 18672
rect 30925 18667 30991 18670
rect 30925 18594 30991 18597
rect 36494 18594 36554 18670
rect 44081 18667 44147 18670
rect 30925 18592 36554 18594
rect 30925 18536 30930 18592
rect 30986 18536 36554 18592
rect 30925 18534 36554 18536
rect 48773 18594 48839 18597
rect 50200 18594 51000 18624
rect 48773 18592 51000 18594
rect 48773 18536 48778 18592
rect 48834 18536 51000 18592
rect 48773 18534 51000 18536
rect 30925 18531 30991 18534
rect 48773 18531 48839 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 31937 18458 32003 18461
rect 35893 18458 35959 18461
rect 31937 18456 35959 18458
rect 31937 18400 31942 18456
rect 31998 18400 35898 18456
rect 35954 18400 35959 18456
rect 31937 18398 35959 18400
rect 31937 18395 32003 18398
rect 35893 18395 35959 18398
rect 0 18322 800 18352
rect 1761 18322 1827 18325
rect 0 18320 1827 18322
rect 0 18264 1766 18320
rect 1822 18264 1827 18320
rect 0 18262 1827 18264
rect 0 18232 800 18262
rect 1761 18259 1827 18262
rect 13905 18322 13971 18325
rect 25129 18322 25195 18325
rect 25957 18322 26023 18325
rect 40309 18322 40375 18325
rect 13905 18320 22110 18322
rect 13905 18264 13910 18320
rect 13966 18264 22110 18320
rect 13905 18262 22110 18264
rect 13905 18259 13971 18262
rect 22050 18186 22110 18262
rect 25129 18320 40375 18322
rect 25129 18264 25134 18320
rect 25190 18264 25962 18320
rect 26018 18264 40314 18320
rect 40370 18264 40375 18320
rect 25129 18262 40375 18264
rect 25129 18259 25195 18262
rect 25957 18259 26023 18262
rect 40309 18259 40375 18262
rect 25037 18186 25103 18189
rect 26233 18186 26299 18189
rect 22050 18184 26299 18186
rect 22050 18128 25042 18184
rect 25098 18128 26238 18184
rect 26294 18128 26299 18184
rect 22050 18126 26299 18128
rect 25037 18123 25103 18126
rect 26233 18123 26299 18126
rect 27654 18124 27660 18188
rect 27724 18186 27730 18188
rect 28441 18186 28507 18189
rect 27724 18184 28507 18186
rect 27724 18128 28446 18184
rect 28502 18128 28507 18184
rect 27724 18126 28507 18128
rect 27724 18124 27730 18126
rect 28441 18123 28507 18126
rect 30097 18186 30163 18189
rect 41137 18186 41203 18189
rect 30097 18184 41203 18186
rect 30097 18128 30102 18184
rect 30158 18128 41142 18184
rect 41198 18128 41203 18184
rect 30097 18126 41203 18128
rect 30097 18123 30163 18126
rect 41137 18123 41203 18126
rect 49417 18186 49483 18189
rect 50200 18186 51000 18216
rect 49417 18184 51000 18186
rect 49417 18128 49422 18184
rect 49478 18128 51000 18184
rect 49417 18126 51000 18128
rect 49417 18123 49483 18126
rect 50200 18096 51000 18126
rect 17769 18050 17835 18053
rect 19333 18050 19399 18053
rect 17769 18048 19399 18050
rect 17769 17992 17774 18048
rect 17830 17992 19338 18048
rect 19394 17992 19399 18048
rect 17769 17990 19399 17992
rect 17769 17987 17835 17990
rect 19333 17987 19399 17990
rect 23657 18050 23723 18053
rect 25262 18050 25268 18052
rect 23657 18048 25268 18050
rect 23657 17992 23662 18048
rect 23718 17992 25268 18048
rect 23657 17990 25268 17992
rect 23657 17987 23723 17990
rect 25262 17988 25268 17990
rect 25332 17988 25338 18052
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 37365 17914 37431 17917
rect 40217 17914 40283 17917
rect 37365 17912 40283 17914
rect 37365 17856 37370 17912
rect 37426 17856 40222 17912
rect 40278 17856 40283 17912
rect 37365 17854 40283 17856
rect 37365 17851 37431 17854
rect 40217 17851 40283 17854
rect 19517 17778 19583 17781
rect 22829 17778 22895 17781
rect 19517 17776 22895 17778
rect 19517 17720 19522 17776
rect 19578 17720 22834 17776
rect 22890 17720 22895 17776
rect 19517 17718 22895 17720
rect 19517 17715 19583 17718
rect 22829 17715 22895 17718
rect 41965 17778 42031 17781
rect 46054 17778 46060 17780
rect 41965 17776 46060 17778
rect 41965 17720 41970 17776
rect 42026 17720 46060 17776
rect 41965 17718 46060 17720
rect 41965 17715 42031 17718
rect 46054 17716 46060 17718
rect 46124 17716 46130 17780
rect 49325 17778 49391 17781
rect 50200 17778 51000 17808
rect 49325 17776 51000 17778
rect 49325 17720 49330 17776
rect 49386 17720 51000 17776
rect 49325 17718 51000 17720
rect 49325 17715 49391 17718
rect 50200 17688 51000 17718
rect 0 17506 800 17536
rect 1761 17506 1827 17509
rect 0 17504 1827 17506
rect 0 17448 1766 17504
rect 1822 17448 1827 17504
rect 0 17446 1827 17448
rect 0 17416 800 17446
rect 1761 17443 1827 17446
rect 30005 17506 30071 17509
rect 30373 17506 30439 17509
rect 35525 17506 35591 17509
rect 30005 17504 35591 17506
rect 30005 17448 30010 17504
rect 30066 17448 30378 17504
rect 30434 17448 35530 17504
rect 35586 17448 35591 17504
rect 30005 17446 35591 17448
rect 30005 17443 30071 17446
rect 30373 17443 30439 17446
rect 35525 17443 35591 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 22369 17370 22435 17373
rect 27705 17370 27771 17373
rect 22369 17368 27771 17370
rect 22369 17312 22374 17368
rect 22430 17312 27710 17368
rect 27766 17312 27771 17368
rect 22369 17310 27771 17312
rect 22369 17307 22435 17310
rect 10501 17234 10567 17237
rect 23657 17234 23723 17237
rect 10501 17232 23723 17234
rect 10501 17176 10506 17232
rect 10562 17176 23662 17232
rect 23718 17176 23723 17232
rect 10501 17174 23723 17176
rect 10501 17171 10567 17174
rect 23657 17171 23723 17174
rect 27478 17234 27538 17310
rect 27705 17307 27771 17310
rect 31017 17370 31083 17373
rect 31845 17370 31911 17373
rect 31017 17368 31911 17370
rect 31017 17312 31022 17368
rect 31078 17312 31850 17368
rect 31906 17312 31911 17368
rect 31017 17310 31911 17312
rect 31017 17307 31083 17310
rect 31845 17307 31911 17310
rect 32397 17370 32463 17373
rect 34053 17370 34119 17373
rect 32397 17368 34119 17370
rect 32397 17312 32402 17368
rect 32458 17312 34058 17368
rect 34114 17312 34119 17368
rect 32397 17310 34119 17312
rect 32397 17307 32463 17310
rect 34053 17307 34119 17310
rect 49325 17370 49391 17373
rect 50200 17370 51000 17400
rect 49325 17368 51000 17370
rect 49325 17312 49330 17368
rect 49386 17312 51000 17368
rect 49325 17310 51000 17312
rect 49325 17307 49391 17310
rect 50200 17280 51000 17310
rect 42701 17234 42767 17237
rect 27478 17232 42767 17234
rect 27478 17176 42706 17232
rect 42762 17176 42767 17232
rect 27478 17174 42767 17176
rect 0 17098 800 17128
rect 1025 17098 1091 17101
rect 0 17096 1091 17098
rect 0 17040 1030 17096
rect 1086 17040 1091 17096
rect 0 17038 1091 17040
rect 0 17008 800 17038
rect 1025 17035 1091 17038
rect 11881 17098 11947 17101
rect 14222 17098 14228 17100
rect 11881 17096 14228 17098
rect 11881 17040 11886 17096
rect 11942 17040 14228 17096
rect 11881 17038 14228 17040
rect 11881 17035 11947 17038
rect 14222 17036 14228 17038
rect 14292 17036 14298 17100
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 14457 16826 14523 16829
rect 18965 16826 19031 16829
rect 27478 16826 27538 17174
rect 42701 17171 42767 17174
rect 27981 17098 28047 17101
rect 49049 17098 49115 17101
rect 27981 17096 49115 17098
rect 27981 17040 27986 17096
rect 28042 17040 49054 17096
rect 49110 17040 49115 17096
rect 27981 17038 49115 17040
rect 27981 17035 28047 17038
rect 49049 17035 49115 17038
rect 48773 16962 48839 16965
rect 50200 16962 51000 16992
rect 48773 16960 51000 16962
rect 48773 16904 48778 16960
rect 48834 16904 51000 16960
rect 48773 16902 51000 16904
rect 48773 16899 48839 16902
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 50200 16872 51000 16902
rect 42946 16831 43262 16832
rect 28625 16826 28691 16829
rect 14457 16824 22110 16826
rect 14457 16768 14462 16824
rect 14518 16768 18970 16824
rect 19026 16768 22110 16824
rect 14457 16766 22110 16768
rect 27478 16824 28691 16826
rect 27478 16768 28630 16824
rect 28686 16768 28691 16824
rect 27478 16766 28691 16768
rect 14457 16763 14523 16766
rect 18965 16763 19031 16766
rect 0 16690 800 16720
rect 933 16690 999 16693
rect 0 16688 999 16690
rect 0 16632 938 16688
rect 994 16632 999 16688
rect 0 16630 999 16632
rect 0 16600 800 16630
rect 933 16627 999 16630
rect 10869 16690 10935 16693
rect 15101 16690 15167 16693
rect 10869 16688 15167 16690
rect 10869 16632 10874 16688
rect 10930 16632 15106 16688
rect 15162 16632 15167 16688
rect 10869 16630 15167 16632
rect 22050 16690 22110 16766
rect 28625 16763 28691 16766
rect 25957 16690 26023 16693
rect 22050 16688 26023 16690
rect 22050 16632 25962 16688
rect 26018 16632 26023 16688
rect 22050 16630 26023 16632
rect 10869 16627 10935 16630
rect 15101 16627 15167 16630
rect 25957 16627 26023 16630
rect 28073 16690 28139 16693
rect 49141 16690 49207 16693
rect 28073 16688 49207 16690
rect 28073 16632 28078 16688
rect 28134 16632 49146 16688
rect 49202 16632 49207 16688
rect 28073 16630 49207 16632
rect 28073 16627 28139 16630
rect 49141 16627 49207 16630
rect 11605 16554 11671 16557
rect 16389 16554 16455 16557
rect 11605 16552 16455 16554
rect 11605 16496 11610 16552
rect 11666 16496 16394 16552
rect 16450 16496 16455 16552
rect 11605 16494 16455 16496
rect 11605 16491 11671 16494
rect 16389 16491 16455 16494
rect 25957 16554 26023 16557
rect 49141 16554 49207 16557
rect 25957 16552 49207 16554
rect 25957 16496 25962 16552
rect 26018 16496 49146 16552
rect 49202 16496 49207 16552
rect 25957 16494 49207 16496
rect 25957 16491 26023 16494
rect 49141 16491 49207 16494
rect 49325 16554 49391 16557
rect 50200 16554 51000 16584
rect 49325 16552 51000 16554
rect 49325 16496 49330 16552
rect 49386 16496 51000 16552
rect 49325 16494 51000 16496
rect 49325 16491 49391 16494
rect 50200 16464 51000 16494
rect 24945 16418 25011 16421
rect 26233 16418 26299 16421
rect 24945 16416 26299 16418
rect 24945 16360 24950 16416
rect 25006 16360 26238 16416
rect 26294 16360 26299 16416
rect 24945 16358 26299 16360
rect 24945 16355 25011 16358
rect 26233 16355 26299 16358
rect 30557 16418 30623 16421
rect 32397 16418 32463 16421
rect 30557 16416 32463 16418
rect 30557 16360 30562 16416
rect 30618 16360 32402 16416
rect 32458 16360 32463 16416
rect 30557 16358 32463 16360
rect 30557 16355 30623 16358
rect 32397 16355 32463 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1025 16282 1091 16285
rect 0 16280 1091 16282
rect 0 16224 1030 16280
rect 1086 16224 1091 16280
rect 0 16222 1091 16224
rect 0 16192 800 16222
rect 1025 16219 1091 16222
rect 14273 16146 14339 16149
rect 15837 16146 15903 16149
rect 27245 16146 27311 16149
rect 34881 16146 34947 16149
rect 14273 16144 22110 16146
rect 14273 16088 14278 16144
rect 14334 16088 15842 16144
rect 15898 16088 22110 16144
rect 14273 16086 22110 16088
rect 14273 16083 14339 16086
rect 15837 16083 15903 16086
rect 13169 16010 13235 16013
rect 14549 16010 14615 16013
rect 13169 16008 14615 16010
rect 13169 15952 13174 16008
rect 13230 15952 14554 16008
rect 14610 15952 14615 16008
rect 13169 15950 14615 15952
rect 22050 16010 22110 16086
rect 27245 16144 34947 16146
rect 27245 16088 27250 16144
rect 27306 16088 34886 16144
rect 34942 16088 34947 16144
rect 27245 16086 34947 16088
rect 27245 16083 27311 16086
rect 34881 16083 34947 16086
rect 49417 16146 49483 16149
rect 50200 16146 51000 16176
rect 49417 16144 51000 16146
rect 49417 16088 49422 16144
rect 49478 16088 51000 16144
rect 49417 16086 51000 16088
rect 49417 16083 49483 16086
rect 50200 16056 51000 16086
rect 29637 16010 29703 16013
rect 30097 16010 30163 16013
rect 22050 16008 30163 16010
rect 22050 15952 29642 16008
rect 29698 15952 30102 16008
rect 30158 15952 30163 16008
rect 22050 15950 30163 15952
rect 13169 15947 13235 15950
rect 14549 15947 14615 15950
rect 29637 15947 29703 15950
rect 30097 15947 30163 15950
rect 35709 16010 35775 16013
rect 49141 16010 49207 16013
rect 35709 16008 49207 16010
rect 35709 15952 35714 16008
rect 35770 15952 49146 16008
rect 49202 15952 49207 16008
rect 35709 15950 49207 15952
rect 35709 15947 35775 15950
rect 49141 15947 49207 15950
rect 0 15874 800 15904
rect 1025 15874 1091 15877
rect 0 15872 1091 15874
rect 0 15816 1030 15872
rect 1086 15816 1091 15872
rect 0 15814 1091 15816
rect 0 15784 800 15814
rect 1025 15811 1091 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 49325 15738 49391 15741
rect 50200 15738 51000 15768
rect 49325 15736 51000 15738
rect 49325 15680 49330 15736
rect 49386 15680 51000 15736
rect 49325 15678 51000 15680
rect 49325 15675 49391 15678
rect 50200 15648 51000 15678
rect 10777 15602 10843 15605
rect 16205 15602 16271 15605
rect 18413 15602 18479 15605
rect 10777 15600 18479 15602
rect 10777 15544 10782 15600
rect 10838 15544 16210 15600
rect 16266 15544 18418 15600
rect 18474 15544 18479 15600
rect 10777 15542 18479 15544
rect 10777 15539 10843 15542
rect 16205 15539 16271 15542
rect 18413 15539 18479 15542
rect 28349 15602 28415 15605
rect 41321 15602 41387 15605
rect 28349 15600 41387 15602
rect 28349 15544 28354 15600
rect 28410 15544 41326 15600
rect 41382 15544 41387 15600
rect 28349 15542 41387 15544
rect 28349 15539 28415 15542
rect 41321 15539 41387 15542
rect 0 15466 800 15496
rect 933 15466 999 15469
rect 0 15464 999 15466
rect 0 15408 938 15464
rect 994 15408 999 15464
rect 0 15406 999 15408
rect 0 15376 800 15406
rect 933 15403 999 15406
rect 16849 15466 16915 15469
rect 21449 15466 21515 15469
rect 21817 15466 21883 15469
rect 16849 15464 21883 15466
rect 16849 15408 16854 15464
rect 16910 15408 21454 15464
rect 21510 15408 21822 15464
rect 21878 15408 21883 15464
rect 16849 15406 21883 15408
rect 16849 15403 16915 15406
rect 21449 15403 21515 15406
rect 21817 15403 21883 15406
rect 26969 15466 27035 15469
rect 34605 15466 34671 15469
rect 39297 15466 39363 15469
rect 26969 15464 31770 15466
rect 26969 15408 26974 15464
rect 27030 15408 31770 15464
rect 26969 15406 31770 15408
rect 26969 15403 27035 15406
rect 10501 15330 10567 15333
rect 17309 15330 17375 15333
rect 10501 15328 17375 15330
rect 10501 15272 10506 15328
rect 10562 15272 17314 15328
rect 17370 15272 17375 15328
rect 10501 15270 17375 15272
rect 31710 15330 31770 15406
rect 34605 15464 39363 15466
rect 34605 15408 34610 15464
rect 34666 15408 39302 15464
rect 39358 15408 39363 15464
rect 34605 15406 39363 15408
rect 34605 15403 34671 15406
rect 39297 15403 39363 15406
rect 35433 15330 35499 15333
rect 31710 15328 35499 15330
rect 31710 15272 35438 15328
rect 35494 15272 35499 15328
rect 31710 15270 35499 15272
rect 10501 15267 10567 15270
rect 17309 15267 17375 15270
rect 35433 15267 35499 15270
rect 49325 15330 49391 15333
rect 50200 15330 51000 15360
rect 49325 15328 51000 15330
rect 49325 15272 49330 15328
rect 49386 15272 51000 15328
rect 49325 15270 51000 15272
rect 49325 15267 49391 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 50200 15240 51000 15270
rect 47946 15199 48262 15200
rect 22369 15194 22435 15197
rect 27521 15194 27587 15197
rect 27654 15194 27660 15196
rect 22369 15192 27660 15194
rect 22369 15136 22374 15192
rect 22430 15136 27526 15192
rect 27582 15136 27660 15192
rect 22369 15134 27660 15136
rect 22369 15131 22435 15134
rect 27521 15131 27587 15134
rect 27654 15132 27660 15134
rect 27724 15132 27730 15196
rect 30649 15194 30715 15197
rect 36997 15194 37063 15197
rect 30649 15192 37063 15194
rect 30649 15136 30654 15192
rect 30710 15136 37002 15192
rect 37058 15136 37063 15192
rect 30649 15134 37063 15136
rect 30649 15131 30715 15134
rect 36997 15131 37063 15134
rect 0 15058 800 15088
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14968 800 14998
rect 933 14995 999 14998
rect 26233 15058 26299 15061
rect 27245 15058 27311 15061
rect 48865 15058 48931 15061
rect 26233 15056 48931 15058
rect 26233 15000 26238 15056
rect 26294 15000 27250 15056
rect 27306 15000 48870 15056
rect 48926 15000 48931 15056
rect 26233 14998 48931 15000
rect 26233 14995 26299 14998
rect 27245 14995 27311 14998
rect 48865 14995 48931 14998
rect 23841 14922 23907 14925
rect 49141 14922 49207 14925
rect 23841 14920 49207 14922
rect 23841 14864 23846 14920
rect 23902 14864 49146 14920
rect 49202 14864 49207 14920
rect 23841 14862 49207 14864
rect 23841 14859 23907 14862
rect 49141 14859 49207 14862
rect 49325 14922 49391 14925
rect 50200 14922 51000 14952
rect 49325 14920 51000 14922
rect 49325 14864 49330 14920
rect 49386 14864 51000 14920
rect 49325 14862 51000 14864
rect 49325 14859 49391 14862
rect 50200 14832 51000 14862
rect 27981 14786 28047 14789
rect 30373 14786 30439 14789
rect 27981 14784 30439 14786
rect 27981 14728 27986 14784
rect 28042 14728 30378 14784
rect 30434 14728 30439 14784
rect 27981 14726 30439 14728
rect 27981 14723 28047 14726
rect 30373 14723 30439 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 933 14650 999 14653
rect 0 14648 999 14650
rect 0 14592 938 14648
rect 994 14592 999 14648
rect 0 14590 999 14592
rect 0 14560 800 14590
rect 933 14587 999 14590
rect 19609 14650 19675 14653
rect 22001 14650 22067 14653
rect 36169 14650 36235 14653
rect 36353 14650 36419 14653
rect 19609 14648 22754 14650
rect 19609 14592 19614 14648
rect 19670 14592 22006 14648
rect 22062 14592 22754 14648
rect 19609 14590 22754 14592
rect 19609 14587 19675 14590
rect 22001 14587 22067 14590
rect 13997 14514 14063 14517
rect 16573 14514 16639 14517
rect 13997 14512 16639 14514
rect 13997 14456 14002 14512
rect 14058 14456 16578 14512
rect 16634 14456 16639 14512
rect 13997 14454 16639 14456
rect 13997 14451 14063 14454
rect 16573 14451 16639 14454
rect 19885 14514 19951 14517
rect 22553 14514 22619 14517
rect 19885 14512 22619 14514
rect 19885 14456 19890 14512
rect 19946 14456 22558 14512
rect 22614 14456 22619 14512
rect 19885 14454 22619 14456
rect 22694 14514 22754 14590
rect 36169 14648 36419 14650
rect 36169 14592 36174 14648
rect 36230 14592 36358 14648
rect 36414 14592 36419 14648
rect 36169 14590 36419 14592
rect 36169 14587 36235 14590
rect 36353 14587 36419 14590
rect 49049 14514 49115 14517
rect 22694 14512 49115 14514
rect 22694 14456 49054 14512
rect 49110 14456 49115 14512
rect 22694 14454 49115 14456
rect 19885 14451 19951 14454
rect 22553 14451 22619 14454
rect 49049 14451 49115 14454
rect 49233 14514 49299 14517
rect 50200 14514 51000 14544
rect 49233 14512 51000 14514
rect 49233 14456 49238 14512
rect 49294 14456 51000 14512
rect 49233 14454 51000 14456
rect 49233 14451 49299 14454
rect 50200 14424 51000 14454
rect 10409 14378 10475 14381
rect 21173 14378 21239 14381
rect 35709 14378 35775 14381
rect 10409 14376 35775 14378
rect 10409 14320 10414 14376
rect 10470 14320 21178 14376
rect 21234 14320 35714 14376
rect 35770 14320 35775 14376
rect 10409 14318 35775 14320
rect 10409 14315 10475 14318
rect 21173 14315 21239 14318
rect 35709 14315 35775 14318
rect 0 14242 800 14272
rect 1025 14242 1091 14245
rect 0 14240 1091 14242
rect 0 14184 1030 14240
rect 1086 14184 1091 14240
rect 0 14182 1091 14184
rect 0 14152 800 14182
rect 1025 14179 1091 14182
rect 35433 14242 35499 14245
rect 36629 14242 36695 14245
rect 35433 14240 36695 14242
rect 35433 14184 35438 14240
rect 35494 14184 36634 14240
rect 36690 14184 36695 14240
rect 35433 14182 36695 14184
rect 35433 14179 35499 14182
rect 36629 14179 36695 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 49233 14106 49299 14109
rect 50200 14106 51000 14136
rect 49233 14104 51000 14106
rect 49233 14048 49238 14104
rect 49294 14048 51000 14104
rect 49233 14046 51000 14048
rect 49233 14043 49299 14046
rect 50200 14016 51000 14046
rect 11237 13970 11303 13973
rect 19609 13970 19675 13973
rect 11237 13968 19675 13970
rect 11237 13912 11242 13968
rect 11298 13912 19614 13968
rect 19670 13912 19675 13968
rect 11237 13910 19675 13912
rect 11237 13907 11303 13910
rect 0 13834 800 13864
rect 1761 13834 1827 13837
rect 0 13832 1827 13834
rect 0 13776 1766 13832
rect 1822 13776 1827 13832
rect 0 13774 1827 13776
rect 0 13744 800 13774
rect 1761 13771 1827 13774
rect 16481 13834 16547 13837
rect 17309 13834 17375 13837
rect 16481 13832 17375 13834
rect 16481 13776 16486 13832
rect 16542 13776 17314 13832
rect 17370 13776 17375 13832
rect 16481 13774 17375 13776
rect 16481 13771 16547 13774
rect 17309 13771 17375 13774
rect 14365 13698 14431 13701
rect 17125 13698 17191 13701
rect 14365 13696 17191 13698
rect 14365 13640 14370 13696
rect 14426 13640 17130 13696
rect 17186 13640 17191 13696
rect 14365 13638 17191 13640
rect 14365 13635 14431 13638
rect 17125 13635 17191 13638
rect 17309 13698 17375 13701
rect 17542 13698 17602 13910
rect 19609 13907 19675 13910
rect 17309 13696 17602 13698
rect 17309 13640 17314 13696
rect 17370 13640 17602 13696
rect 17309 13638 17602 13640
rect 48221 13698 48287 13701
rect 50200 13698 51000 13728
rect 48221 13696 51000 13698
rect 48221 13640 48226 13696
rect 48282 13640 51000 13696
rect 48221 13638 51000 13640
rect 17309 13635 17375 13638
rect 48221 13635 48287 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 50200 13608 51000 13638
rect 42946 13567 43262 13568
rect 0 13426 800 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 800 13366
rect 3509 13363 3575 13366
rect 14733 13426 14799 13429
rect 17125 13426 17191 13429
rect 14733 13424 17191 13426
rect 14733 13368 14738 13424
rect 14794 13368 17130 13424
rect 17186 13368 17191 13424
rect 14733 13366 17191 13368
rect 14733 13363 14799 13366
rect 17125 13363 17191 13366
rect 31661 13426 31727 13429
rect 35801 13426 35867 13429
rect 31661 13424 35867 13426
rect 31661 13368 31666 13424
rect 31722 13368 35806 13424
rect 35862 13368 35867 13424
rect 31661 13366 35867 13368
rect 31661 13363 31727 13366
rect 35801 13363 35867 13366
rect 18781 13290 18847 13293
rect 30557 13290 30623 13293
rect 35157 13290 35223 13293
rect 18781 13288 35223 13290
rect 18781 13232 18786 13288
rect 18842 13232 30562 13288
rect 30618 13232 35162 13288
rect 35218 13232 35223 13288
rect 18781 13230 35223 13232
rect 18781 13227 18847 13230
rect 30557 13227 30623 13230
rect 35157 13227 35223 13230
rect 49141 13290 49207 13293
rect 50200 13290 51000 13320
rect 49141 13288 51000 13290
rect 49141 13232 49146 13288
rect 49202 13232 51000 13288
rect 49141 13230 51000 13232
rect 49141 13227 49207 13230
rect 50200 13200 51000 13230
rect 11145 13154 11211 13157
rect 14457 13154 14523 13157
rect 11145 13152 14523 13154
rect 11145 13096 11150 13152
rect 11206 13096 14462 13152
rect 14518 13096 14523 13152
rect 11145 13094 14523 13096
rect 11145 13091 11211 13094
rect 14457 13091 14523 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 22921 13018 22987 13021
rect 26417 13018 26483 13021
rect 22921 13016 26483 13018
rect 22921 12960 22926 13016
rect 22982 12960 26422 13016
rect 26478 12960 26483 13016
rect 22921 12958 26483 12960
rect 22921 12955 22987 12958
rect 26417 12955 26483 12958
rect 11145 12882 11211 12885
rect 15837 12882 15903 12885
rect 11145 12880 15903 12882
rect 11145 12824 11150 12880
rect 11206 12824 15842 12880
rect 15898 12824 15903 12880
rect 11145 12822 15903 12824
rect 11145 12819 11211 12822
rect 15837 12819 15903 12822
rect 16430 12820 16436 12884
rect 16500 12882 16506 12884
rect 20713 12882 20779 12885
rect 16500 12880 20779 12882
rect 16500 12824 20718 12880
rect 20774 12824 20779 12880
rect 16500 12822 20779 12824
rect 16500 12820 16506 12822
rect 20713 12819 20779 12822
rect 21725 12882 21791 12885
rect 26049 12882 26115 12885
rect 21725 12880 26115 12882
rect 21725 12824 21730 12880
rect 21786 12824 26054 12880
rect 26110 12824 26115 12880
rect 21725 12822 26115 12824
rect 21725 12819 21791 12822
rect 26049 12819 26115 12822
rect 49141 12882 49207 12885
rect 50200 12882 51000 12912
rect 49141 12880 51000 12882
rect 49141 12824 49146 12880
rect 49202 12824 51000 12880
rect 49141 12822 51000 12824
rect 49141 12819 49207 12822
rect 50200 12792 51000 12822
rect 13445 12746 13511 12749
rect 13721 12746 13787 12749
rect 13445 12744 13787 12746
rect 13445 12688 13450 12744
rect 13506 12688 13726 12744
rect 13782 12688 13787 12744
rect 13445 12686 13787 12688
rect 13445 12683 13511 12686
rect 13721 12683 13787 12686
rect 14222 12684 14228 12748
rect 14292 12746 14298 12748
rect 16205 12746 16271 12749
rect 14292 12744 16271 12746
rect 14292 12688 16210 12744
rect 16266 12688 16271 12744
rect 14292 12686 16271 12688
rect 14292 12684 14298 12686
rect 16205 12683 16271 12686
rect 28533 12746 28599 12749
rect 40033 12746 40099 12749
rect 28533 12744 40099 12746
rect 28533 12688 28538 12744
rect 28594 12688 40038 12744
rect 40094 12688 40099 12744
rect 28533 12686 40099 12688
rect 28533 12683 28599 12686
rect 40033 12683 40099 12686
rect 0 12610 800 12640
rect 1209 12610 1275 12613
rect 0 12608 1275 12610
rect 0 12552 1214 12608
rect 1270 12552 1275 12608
rect 0 12550 1275 12552
rect 0 12520 800 12550
rect 1209 12547 1275 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 0 12202 800 12232
rect 1209 12202 1275 12205
rect 0 12200 1275 12202
rect 0 12144 1214 12200
rect 1270 12144 1275 12200
rect 0 12142 1275 12144
rect 0 12112 800 12142
rect 1209 12139 1275 12142
rect 13813 12202 13879 12205
rect 22369 12202 22435 12205
rect 30097 12202 30163 12205
rect 13813 12200 19350 12202
rect 13813 12144 13818 12200
rect 13874 12144 19350 12200
rect 13813 12142 19350 12144
rect 13813 12139 13879 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 13353 11930 13419 11933
rect 17217 11930 17283 11933
rect 13353 11928 17283 11930
rect 13353 11872 13358 11928
rect 13414 11872 17222 11928
rect 17278 11872 17283 11928
rect 13353 11870 17283 11872
rect 19290 11930 19350 12142
rect 22369 12200 30163 12202
rect 22369 12144 22374 12200
rect 22430 12144 30102 12200
rect 30158 12144 30163 12200
rect 22369 12142 30163 12144
rect 22369 12139 22435 12142
rect 30097 12139 30163 12142
rect 19977 12066 20043 12069
rect 22461 12066 22527 12069
rect 19977 12064 22527 12066
rect 19977 12008 19982 12064
rect 20038 12008 22466 12064
rect 22522 12008 22527 12064
rect 19977 12006 22527 12008
rect 19977 12003 20043 12006
rect 22461 12003 22527 12006
rect 49141 12066 49207 12069
rect 50200 12066 51000 12096
rect 49141 12064 51000 12066
rect 49141 12008 49146 12064
rect 49202 12008 51000 12064
rect 49141 12006 51000 12008
rect 49141 12003 49207 12006
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 50200 11976 51000 12006
rect 47946 11935 48262 11936
rect 20529 11930 20595 11933
rect 27429 11930 27495 11933
rect 19290 11928 27495 11930
rect 19290 11872 20534 11928
rect 20590 11872 27434 11928
rect 27490 11872 27495 11928
rect 19290 11870 27495 11872
rect 13353 11867 13419 11870
rect 17217 11867 17283 11870
rect 20529 11867 20595 11870
rect 27429 11867 27495 11870
rect 0 11794 800 11824
rect 1301 11794 1367 11797
rect 0 11792 1367 11794
rect 0 11736 1306 11792
rect 1362 11736 1367 11792
rect 0 11734 1367 11736
rect 0 11704 800 11734
rect 1301 11731 1367 11734
rect 20529 11794 20595 11797
rect 24945 11794 25011 11797
rect 20529 11792 25011 11794
rect 20529 11736 20534 11792
rect 20590 11736 24950 11792
rect 25006 11736 25011 11792
rect 20529 11734 25011 11736
rect 20529 11731 20595 11734
rect 24945 11731 25011 11734
rect 29637 11794 29703 11797
rect 40401 11794 40467 11797
rect 29637 11792 40467 11794
rect 29637 11736 29642 11792
rect 29698 11736 40406 11792
rect 40462 11736 40467 11792
rect 29637 11734 40467 11736
rect 29637 11731 29703 11734
rect 40401 11731 40467 11734
rect 49141 11658 49207 11661
rect 50200 11658 51000 11688
rect 49141 11656 51000 11658
rect 49141 11600 49146 11656
rect 49202 11600 51000 11656
rect 49141 11598 51000 11600
rect 49141 11595 49207 11598
rect 50200 11568 51000 11598
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 1301 11386 1367 11389
rect 0 11384 1367 11386
rect 0 11328 1306 11384
rect 1362 11328 1367 11384
rect 0 11326 1367 11328
rect 0 11296 800 11326
rect 1301 11323 1367 11326
rect 49233 11250 49299 11253
rect 50200 11250 51000 11280
rect 49233 11248 51000 11250
rect 49233 11192 49238 11248
rect 49294 11192 51000 11248
rect 49233 11190 51000 11192
rect 49233 11187 49299 11190
rect 50200 11160 51000 11190
rect 18505 11114 18571 11117
rect 22461 11114 22527 11117
rect 18505 11112 22527 11114
rect 18505 11056 18510 11112
rect 18566 11056 22466 11112
rect 22522 11056 22527 11112
rect 18505 11054 22527 11056
rect 18505 11051 18571 11054
rect 22461 11051 22527 11054
rect 23841 11114 23907 11117
rect 27705 11114 27771 11117
rect 23841 11112 27771 11114
rect 23841 11056 23846 11112
rect 23902 11056 27710 11112
rect 27766 11056 27771 11112
rect 23841 11054 27771 11056
rect 23841 11051 23907 11054
rect 27705 11051 27771 11054
rect 31385 11114 31451 11117
rect 32305 11114 32371 11117
rect 31385 11112 32371 11114
rect 31385 11056 31390 11112
rect 31446 11056 32310 11112
rect 32366 11056 32371 11112
rect 31385 11054 32371 11056
rect 31385 11051 31451 11054
rect 32305 11051 32371 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 49141 10842 49207 10845
rect 50200 10842 51000 10872
rect 49141 10840 51000 10842
rect 49141 10784 49146 10840
rect 49202 10784 51000 10840
rect 49141 10782 51000 10784
rect 49141 10779 49207 10782
rect 50200 10752 51000 10782
rect 11605 10706 11671 10709
rect 16481 10706 16547 10709
rect 18965 10706 19031 10709
rect 11605 10704 19031 10706
rect 11605 10648 11610 10704
rect 11666 10648 16486 10704
rect 16542 10648 18970 10704
rect 19026 10648 19031 10704
rect 11605 10646 19031 10648
rect 11605 10643 11671 10646
rect 16481 10643 16547 10646
rect 18965 10643 19031 10646
rect 0 10570 800 10600
rect 1301 10570 1367 10573
rect 0 10568 1367 10570
rect 0 10512 1306 10568
rect 1362 10512 1367 10568
rect 0 10510 1367 10512
rect 0 10480 800 10510
rect 1301 10507 1367 10510
rect 13261 10570 13327 10573
rect 34973 10570 35039 10573
rect 13261 10568 35039 10570
rect 13261 10512 13266 10568
rect 13322 10512 34978 10568
rect 35034 10512 35039 10568
rect 13261 10510 35039 10512
rect 13261 10507 13327 10510
rect 34973 10507 35039 10510
rect 49233 10434 49299 10437
rect 50200 10434 51000 10464
rect 49233 10432 51000 10434
rect 49233 10376 49238 10432
rect 49294 10376 51000 10432
rect 49233 10374 51000 10376
rect 49233 10371 49299 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 1209 10162 1275 10165
rect 0 10160 1275 10162
rect 0 10104 1214 10160
rect 1270 10104 1275 10160
rect 0 10102 1275 10104
rect 0 10072 800 10102
rect 1209 10099 1275 10102
rect 14641 10026 14707 10029
rect 15101 10026 15167 10029
rect 14641 10024 15167 10026
rect 14641 9968 14646 10024
rect 14702 9968 15106 10024
rect 15162 9968 15167 10024
rect 14641 9966 15167 9968
rect 14641 9963 14707 9966
rect 15101 9963 15167 9966
rect 49325 10026 49391 10029
rect 50200 10026 51000 10056
rect 49325 10024 51000 10026
rect 49325 9968 49330 10024
rect 49386 9968 51000 10024
rect 49325 9966 51000 9968
rect 49325 9963 49391 9966
rect 50200 9936 51000 9966
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1301 9754 1367 9757
rect 0 9752 1367 9754
rect 0 9696 1306 9752
rect 1362 9696 1367 9752
rect 0 9694 1367 9696
rect 0 9664 800 9694
rect 1301 9691 1367 9694
rect 34421 9618 34487 9621
rect 34697 9618 34763 9621
rect 34421 9616 34763 9618
rect 34421 9560 34426 9616
rect 34482 9560 34702 9616
rect 34758 9560 34763 9616
rect 34421 9558 34763 9560
rect 34421 9555 34487 9558
rect 34697 9555 34763 9558
rect 47301 9618 47367 9621
rect 50200 9618 51000 9648
rect 47301 9616 51000 9618
rect 47301 9560 47306 9616
rect 47362 9560 51000 9616
rect 47301 9558 51000 9560
rect 47301 9555 47367 9558
rect 50200 9528 51000 9558
rect 1761 9482 1827 9485
rect 33685 9482 33751 9485
rect 1761 9480 33751 9482
rect 1761 9424 1766 9480
rect 1822 9424 33690 9480
rect 33746 9424 33751 9480
rect 1761 9422 33751 9424
rect 1761 9419 1827 9422
rect 33685 9419 33751 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9210 49207 9213
rect 50200 9210 51000 9240
rect 49141 9208 51000 9210
rect 49141 9152 49146 9208
rect 49202 9152 51000 9208
rect 49141 9150 51000 9152
rect 49141 9147 49207 9150
rect 50200 9120 51000 9150
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 49233 8802 49299 8805
rect 50200 8802 51000 8832
rect 49233 8800 51000 8802
rect 49233 8744 49238 8800
rect 49294 8744 51000 8800
rect 49233 8742 51000 8744
rect 49233 8739 49299 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 50200 8712 51000 8742
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 49325 8394 49391 8397
rect 50200 8394 51000 8424
rect 49325 8392 51000 8394
rect 49325 8336 49330 8392
rect 49386 8336 51000 8392
rect 49325 8334 51000 8336
rect 49325 8331 49391 8334
rect 50200 8304 51000 8334
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1301 8122 1367 8125
rect 0 8120 1367 8122
rect 0 8064 1306 8120
rect 1362 8064 1367 8120
rect 0 8062 1367 8064
rect 0 8032 800 8062
rect 1301 8059 1367 8062
rect 46841 7986 46907 7989
rect 50200 7986 51000 8016
rect 46841 7984 51000 7986
rect 46841 7928 46846 7984
rect 46902 7928 51000 7984
rect 46841 7926 51000 7928
rect 46841 7923 46907 7926
rect 50200 7896 51000 7926
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 49141 7578 49207 7581
rect 50200 7578 51000 7608
rect 49141 7576 51000 7578
rect 49141 7520 49146 7576
rect 49202 7520 51000 7576
rect 49141 7518 51000 7520
rect 49141 7515 49207 7518
rect 50200 7488 51000 7518
rect 0 7306 800 7336
rect 1301 7306 1367 7309
rect 0 7304 1367 7306
rect 0 7248 1306 7304
rect 1362 7248 1367 7304
rect 0 7246 1367 7248
rect 0 7216 800 7246
rect 1301 7243 1367 7246
rect 49417 7170 49483 7173
rect 50200 7170 51000 7200
rect 49417 7168 51000 7170
rect 49417 7112 49422 7168
rect 49478 7112 51000 7168
rect 49417 7110 51000 7112
rect 49417 7107 49483 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 50200 7080 51000 7110
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 800 6838
rect 1209 6835 1275 6838
rect 49233 6762 49299 6765
rect 50200 6762 51000 6792
rect 49233 6760 51000 6762
rect 49233 6704 49238 6760
rect 49294 6704 51000 6760
rect 49233 6702 51000 6704
rect 49233 6699 49299 6702
rect 50200 6672 51000 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 48681 6354 48747 6357
rect 50200 6354 51000 6384
rect 48681 6352 51000 6354
rect 48681 6296 48686 6352
rect 48742 6296 51000 6352
rect 48681 6294 51000 6296
rect 48681 6291 48747 6294
rect 50200 6264 51000 6294
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5946 49207 5949
rect 50200 5946 51000 5976
rect 49141 5944 51000 5946
rect 49141 5888 49146 5944
rect 49202 5888 51000 5944
rect 49141 5886 51000 5888
rect 49141 5883 49207 5886
rect 50200 5856 51000 5886
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 49417 5538 49483 5541
rect 50200 5538 51000 5568
rect 49417 5536 51000 5538
rect 49417 5480 49422 5536
rect 49478 5480 51000 5536
rect 49417 5478 51000 5480
rect 49417 5475 49483 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 50200 5448 51000 5478
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 49325 5130 49391 5133
rect 50200 5130 51000 5160
rect 49325 5128 51000 5130
rect 49325 5072 49330 5128
rect 49386 5072 51000 5128
rect 49325 5070 51000 5072
rect 49325 5067 49391 5070
rect 50200 5040 51000 5070
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 48313 4722 48379 4725
rect 50200 4722 51000 4752
rect 48313 4720 51000 4722
rect 48313 4664 48318 4720
rect 48374 4664 51000 4720
rect 48313 4662 51000 4664
rect 48313 4659 48379 4662
rect 50200 4632 51000 4662
rect 0 4450 800 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 800 4390
rect 1301 4387 1367 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 5349 4042 5415 4045
rect 24853 4042 24919 4045
rect 5349 4040 24919 4042
rect 5349 3984 5354 4040
rect 5410 3984 24858 4040
rect 24914 3984 24919 4040
rect 5349 3982 24919 3984
rect 5349 3979 5415 3982
rect 24853 3979 24919 3982
rect 49233 3906 49299 3909
rect 50200 3906 51000 3936
rect 49233 3904 51000 3906
rect 49233 3848 49238 3904
rect 49294 3848 51000 3904
rect 49233 3846 51000 3848
rect 49233 3843 49299 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 50200 3816 51000 3846
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 1117 3498 1183 3501
rect 25773 3498 25839 3501
rect 1117 3496 25839 3498
rect 1117 3440 1122 3496
rect 1178 3440 25778 3496
rect 25834 3440 25839 3496
rect 1117 3438 25839 3440
rect 1117 3435 1183 3438
rect 25773 3435 25839 3438
rect 49141 3498 49207 3501
rect 50200 3498 51000 3528
rect 49141 3496 51000 3498
rect 49141 3440 49146 3496
rect 49202 3440 51000 3496
rect 49141 3438 51000 3440
rect 49141 3435 49207 3438
rect 50200 3408 51000 3438
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 48681 3090 48747 3093
rect 50200 3090 51000 3120
rect 48681 3088 51000 3090
rect 48681 3032 48686 3088
rect 48742 3032 51000 3088
rect 48681 3030 51000 3032
rect 48681 3027 48747 3030
rect 50200 3000 51000 3030
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 46841 2682 46907 2685
rect 50200 2682 51000 2712
rect 46841 2680 51000 2682
rect 46841 2624 46846 2680
rect 46902 2624 51000 2680
rect 46841 2622 51000 2624
rect 46841 2619 46907 2622
rect 50200 2592 51000 2622
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 48497 2274 48563 2277
rect 50200 2274 51000 2304
rect 48497 2272 51000 2274
rect 48497 2216 48502 2272
rect 48558 2216 51000 2272
rect 48497 2214 51000 2216
rect 48497 2211 48563 2214
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 50200 2184 51000 2214
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 46749 1866 46815 1869
rect 50200 1866 51000 1896
rect 46749 1864 51000 1866
rect 46749 1808 46754 1864
rect 46810 1808 51000 1864
rect 46749 1806 51000 1808
rect 46749 1803 46815 1806
rect 50200 1776 51000 1806
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
rect 46657 1458 46723 1461
rect 50200 1458 51000 1488
rect 46657 1456 51000 1458
rect 46657 1400 46662 1456
rect 46718 1400 51000 1456
rect 46657 1398 51000 1400
rect 46657 1395 46723 1398
rect 50200 1368 51000 1398
<< via3 >>
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 46060 23488 46124 23492
rect 46060 23432 46110 23488
rect 46110 23432 46124 23488
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 46060 23428 46124 23432
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 25268 22944 25332 22948
rect 25268 22888 25318 22944
rect 25318 22888 25332 22944
rect 25268 22884 25332 22888
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 30420 21584 30484 21588
rect 30420 21528 30434 21584
rect 30434 21528 30484 21584
rect 30420 21524 30484 21528
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 30420 19756 30484 19820
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 16436 19484 16500 19548
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 27660 18124 27724 18188
rect 25268 17988 25332 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 46060 17716 46124 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 14228 17036 14292 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 27660 15132 27724 15196
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 16436 12820 16500 12884
rect 14228 12684 14292 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 16435 19548 16501 19549
rect 16435 19484 16436 19548
rect 16500 19484 16501 19548
rect 16435 19483 16501 19484
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 14227 17100 14293 17101
rect 14227 17036 14228 17100
rect 14292 17036 14293 17100
rect 14227 17035 14293 17036
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 14230 12749 14290 17035
rect 16438 12885 16498 19483
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 16435 12884 16501 12885
rect 16435 12820 16436 12884
rect 16500 12820 16501 12884
rect 16435 12819 16501 12820
rect 14227 12748 14293 12749
rect 14227 12684 14228 12748
rect 14292 12684 14293 12748
rect 14227 12683 14293 12684
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 25267 22948 25333 22949
rect 25267 22884 25268 22948
rect 25332 22884 25333 22948
rect 25267 22883 25333 22884
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 25270 18053 25330 22883
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 30419 21588 30485 21589
rect 30419 21524 30420 21588
rect 30484 21524 30485 21588
rect 30419 21523 30485 21524
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 30422 19821 30482 21523
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 30419 19820 30485 19821
rect 30419 19756 30420 19820
rect 30484 19756 30485 19820
rect 30419 19755 30485 19756
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27659 18188 27725 18189
rect 27659 18124 27660 18188
rect 27724 18124 27725 18188
rect 27659 18123 27725 18124
rect 25267 18052 25333 18053
rect 25267 17988 25268 18052
rect 25332 17988 25333 18052
rect 25267 17987 25333 17988
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 27662 15197 27722 18123
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27659 15196 27725 15197
rect 27659 15132 27660 15196
rect 27724 15132 27725 15196
rect 27659 15131 27725 15132
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 46059 23492 46125 23493
rect 46059 23428 46060 23492
rect 46124 23428 46125 23492
rect 46059 23427 46125 23428
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 46062 17781 46122 23427
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 46059 17780 46125 17781
rect 46059 17716 46060 17780
rect 46124 17716 46125 17780
rect 46059 17715 46125 17716
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform -1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform -1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform -1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform -1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform -1 0 11224 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform -1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform -1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform -1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform -1 0 11224 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform -1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform -1 0 9476 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform -1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform -1 0 16376 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform -1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform -1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform -1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform -1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform -1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform -1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform -1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform -1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform -1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform -1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform -1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1676037725
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform -1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 37904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 37168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 37628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 44804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 39192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 44068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 39836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 45540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 39928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform -1 0 46184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform -1 0 46184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform -1 0 45908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform -1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform -1 0 5612 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1676037725
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1676037725
transform -1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1676037725
transform -1 0 2392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1676037725
transform -1 0 6808 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1676037725
transform -1 0 4232 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform -1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform -1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1676037725
transform -1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1676037725
transform 1 0 13892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform -1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform -1 0 7544 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform -1 0 23736 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform -1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform -1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1676037725
transform -1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform -1 0 21528 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform -1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform -1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1676037725
transform -1 0 21528 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform -1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1676037725
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform -1 0 21528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform -1 0 26680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1676037725
transform -1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1676037725
transform -1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1676037725
transform -1 0 13984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1676037725
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform -1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1676037725
transform -1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1676037725
transform -1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1676037725
transform -1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1676037725
transform -1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1676037725
transform 1 0 11592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1676037725
transform -1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1676037725
transform -1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1676037725
transform -1 0 11408 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1676037725
transform -1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1676037725
transform -1 0 9384 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1676037725
transform -1 0 37076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1676037725
transform -1 0 38640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1676037725
transform 1 0 36800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1676037725
transform -1 0 39100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1676037725
transform -1 0 38180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform -1 0 39192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 37352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 37536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform -1 0 39376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform -1 0 40940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform -1 0 40020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform -1 0 40756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform -1 0 38916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform -1 0 40388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform -1 0 40756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform -1 0 40572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform -1 0 40664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1676037725
transform -1 0 26496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1676037725
transform -1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19504 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform -1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 16744 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 16376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform -1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform -1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform -1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 28244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 28060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform -1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform -1 0 22724 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 30360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform -1 0 37168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 35328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform -1 0 42964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold10_A
timestamp 1676037725
transform -1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1676037725
transform -1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform -1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform -1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform -1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform -1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform -1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform -1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform -1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform -1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform -1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform -1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform -1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform -1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform -1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform -1 0 2852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform -1 0 2300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform -1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform -1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform -1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform -1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform -1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform -1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform -1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform -1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform -1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform -1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform -1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform -1 0 48852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform -1 0 48668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform -1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform -1 0 48852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform -1 0 48668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform -1 0 48668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform -1 0 48024 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform -1 0 48852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform -1 0 47564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform -1 0 49588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform -1 0 46184 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform -1 0 48208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform -1 0 48852 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform -1 0 46828 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform -1 0 47840 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform -1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 47472 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform -1 0 47748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 49128 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform -1 0 48208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 47656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform -1 0 47380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform -1 0 48668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform -1 0 48852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform -1 0 48944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform -1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform -1 0 48668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform -1 0 48852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform -1 0 48852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform -1 0 48668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform -1 0 27048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform -1 0 29716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform -1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform -1 0 31188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform -1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform -1 0 41952 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform -1 0 34868 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform -1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform -1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform -1 0 42780 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform -1 0 47472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform -1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform -1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform -1 0 42780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform -1 0 44620 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform -1 0 44252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform -1 0 43884 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform -1 0 42964 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1676037725
transform -1 0 44068 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1676037725
transform -1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1676037725
transform -1 0 45724 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1676037725
transform -1 0 45356 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1676037725
transform -1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1676037725
transform -1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1676037725
transform -1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1676037725
transform -1 0 31648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1676037725
transform -1 0 25300 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1676037725
transform -1 0 29164 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1676037725
transform -1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1676037725
transform -1 0 29348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1676037725
transform -1 0 29716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1676037725
transform -1 0 31464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1676037725
transform -1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1676037725
transform -1 0 35696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1676037725
transform -1 0 37168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1676037725
transform -1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1676037725
transform -1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1676037725
transform -1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1676037725
transform -1 0 49220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1676037725
transform -1 0 49588 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1676037725
transform -1 0 47932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1676037725
transform -1 0 47932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1676037725
transform -1 0 48024 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1676037725
transform -1 0 44436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1676037725
transform -1 0 45540 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1676037725
transform -1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 27048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24472 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20516 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23460 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform -1 0 22172 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23184 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 27784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30176 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30728 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21896 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 28152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform -1 0 37076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 38456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 38456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform -1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 38640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 35880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 33488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 33672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 28980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform -1 0 42596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 33304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 36892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 38456 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 39284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 39468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 37076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 37260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 35512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 40388 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 41032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 37628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 39376 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 40204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 40020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 37260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 39192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 37444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 41124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 40020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 40940 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 41032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 41492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 35880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 12328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 12696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 31924 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 28152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 26404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__S
timestamp 1676037725
transform -1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 30176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 30176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 27508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 29440 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26680 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 30544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 25576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 30360 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 36064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 34316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 34500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 27600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__S
timestamp 1676037725
transform -1 0 27968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 34040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 29532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 37444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 37076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1
timestamp 1676037725
transform -1 0 29440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__S
timestamp 1676037725
transform -1 0 31924 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 35880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 34592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 36616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 36800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 32752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__S
timestamp 1676037725
transform -1 0 33488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 34316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 34224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 34316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 34500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 30452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__S
timestamp 1676037725
transform -1 0 32016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 31832 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 32292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 29440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 26036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 29072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 32016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 33764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 33304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 30268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 29072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 27784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 35696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 43240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 43884 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__S
timestamp 1676037725
transform -1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 41216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 46276 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 31096 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 42596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 29716 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 43056 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 43424 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 33856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 34040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 42228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 34224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1
timestamp 1676037725
transform -1 0 34592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 36892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 41308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 31740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 41216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 39192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41584 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 41952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 36892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 41400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 36432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 38824 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 39008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 28336 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 28612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21804 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 19136 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23000 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 10488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20148 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18216 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18952 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16192 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 16100 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 15456 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9476 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 12788 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 15180 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 12604 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 11040 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform -1 0 16376 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform -1 0 16008 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform -1 0 16376 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform -1 0 17480 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform -1 0 18676 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform -1 0 11224 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform -1 0 13524 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 17940 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform -1 0 13800 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform -1 0 13524 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255
timestamp 1676037725
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform -1 0 14720 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform -1 0 16008 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform -1 0 8556 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform -1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 16744 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform -1 0 10212 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256
timestamp 1676037725
transform -1 0 11224 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform -1 0 12512 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform -1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform -1 0 12972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform -1 0 13800 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15640 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257
timestamp 1676037725
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform -1 0 11868 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29072 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform -1 0 27048 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 23828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20976 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform -1 0 26128 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 23000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 24104 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24196 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform -1 0 26496 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28888 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28980 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 22540 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform -1 0 18768 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform -1 0 23000 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 28796 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform -1 0 29256 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 34040 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 29900 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform -1 0 35604 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform -1 0 35880 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_247
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1676037725
transform 1 0 26036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1676037725
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1676037725
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_311
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1676037725
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1676037725
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_372
timestamp 1676037725
transform 1 0 35328 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_376
timestamp 1676037725
transform 1 0 35696 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_388
timestamp 1676037725
transform 1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1676037725
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_459
timestamp 1676037725
transform 1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1676037725
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1676037725
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1676037725
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_130
timestamp 1676037725
transform 1 0 13064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1676037725
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_171
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1676037725
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_235
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1676037725
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1676037725
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1676037725
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_301
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_323
timestamp 1676037725
transform 1 0 30820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp 1676037725
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1676037725
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1676037725
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1676037725
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_101
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_113
timestamp 1676037725
transform 1 0 11500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_125
timestamp 1676037725
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1676037725
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_170
timestamp 1676037725
transform 1 0 16744 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_182
timestamp 1676037725
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_236
timestamp 1676037725
transform 1 0 22816 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_242
timestamp 1676037725
transform 1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1676037725
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1676037725
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_387
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_391
timestamp 1676037725
transform 1 0 37076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1676037725
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_479
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_485
timestamp 1676037725
transform 1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1676037725
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1676037725
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_233
timestamp 1676037725
transform 1 0 22540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_240
timestamp 1676037725
transform 1 0 23184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1676037725
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1676037725
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1676037725
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1676037725
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1676037725
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_507
timestamp 1676037725
transform 1 0 47748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_218
timestamp 1676037725
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_234
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1676037725
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_282
timestamp 1676037725
transform 1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_294
timestamp 1676037725
transform 1 0 28152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1676037725
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_385
timestamp 1676037725
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_390
timestamp 1676037725
transform 1 0 36984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1676037725
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_404
timestamp 1676037725
transform 1 0 38272 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_408
timestamp 1676037725
transform 1 0 38640 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_491
timestamp 1676037725
transform 1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_497
timestamp 1676037725
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1676037725
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_201
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1676037725
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1676037725
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_395
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_401
timestamp 1676037725
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_409
timestamp 1676037725
transform 1 0 38732 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_413
timestamp 1676037725
transform 1 0 39100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_425
timestamp 1676037725
transform 1 0 40204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_437
timestamp 1676037725
transform 1 0 41308 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1676037725
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1676037725
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_461
timestamp 1676037725
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1676037725
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1676037725
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_192
timestamp 1676037725
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1676037725
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1676037725
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_399
timestamp 1676037725
transform 1 0 37812 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_403
timestamp 1676037725
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1676037725
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1676037725
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1676037725
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_469
timestamp 1676037725
transform 1 0 44252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_481
timestamp 1676037725
transform 1 0 45356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_493
timestamp 1676037725
transform 1 0 46460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1676037725
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1676037725
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1676037725
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_204
timestamp 1676037725
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_216
timestamp 1676037725
transform 1 0 20976 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_224
timestamp 1676037725
transform 1 0 21712 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_227
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_239
timestamp 1676037725
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1676037725
transform 1 0 47564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1676037725
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1676037725
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1676037725
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_196
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_208
timestamp 1676037725
transform 1 0 20240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_216
timestamp 1676037725
transform 1 0 20976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1676037725
transform 1 0 22816 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1676037725
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_252
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1676037725
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1676037725
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_327
timestamp 1676037725
transform 1 0 31188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_342
timestamp 1676037725
transform 1 0 32568 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1676037725
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_358
timestamp 1676037725
transform 1 0 34040 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_370
timestamp 1676037725
transform 1 0 35144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1676037725
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_396
timestamp 1676037725
transform 1 0 37536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1676037725
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_410
timestamp 1676037725
transform 1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_414
timestamp 1676037725
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_426
timestamp 1676037725
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1676037725
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1676037725
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_479
timestamp 1676037725
transform 1 0 45172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_491
timestamp 1676037725
transform 1 0 46276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_9
timestamp 1676037725
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_160
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1676037725
transform 1 0 16560 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_191
timestamp 1676037725
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1676037725
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_225
timestamp 1676037725
transform 1 0 21804 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1676037725
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_314
timestamp 1676037725
transform 1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_323
timestamp 1676037725
transform 1 0 30820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_334
timestamp 1676037725
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_338
timestamp 1676037725
transform 1 0 32200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_348
timestamp 1676037725
transform 1 0 33120 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_352
timestamp 1676037725
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_395
timestamp 1676037725
transform 1 0 37444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_398
timestamp 1676037725
transform 1 0 37720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_404
timestamp 1676037725
transform 1 0 38272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_412
timestamp 1676037725
transform 1 0 39008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1676037725
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1676037725
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_160
timestamp 1676037725
transform 1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1676037725
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_247
timestamp 1676037725
transform 1 0 23828 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_251
timestamp 1676037725
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1676037725
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1676037725
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1676037725
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_359
timestamp 1676037725
transform 1 0 34132 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_367
timestamp 1676037725
transform 1 0 34868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_379
timestamp 1676037725
transform 1 0 35972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1676037725
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_410
timestamp 1676037725
transform 1 0 38824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_414
timestamp 1676037725
transform 1 0 39192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_422
timestamp 1676037725
transform 1 0 39928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1676037725
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1676037725
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_471
timestamp 1676037725
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_483
timestamp 1676037725
transform 1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1676037725
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_146
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1676037725
transform 1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_162
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_269
timestamp 1676037725
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_281
timestamp 1676037725
transform 1 0 26956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_292
timestamp 1676037725
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1676037725
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_314
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1676037725
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_342
timestamp 1676037725
transform 1 0 32568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_348
timestamp 1676037725
transform 1 0 33120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_359
timestamp 1676037725
transform 1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_376
timestamp 1676037725
transform 1 0 35696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_384
timestamp 1676037725
transform 1 0 36432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_388
timestamp 1676037725
transform 1 0 36800 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_396
timestamp 1676037725
transform 1 0 37536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_400
timestamp 1676037725
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_412
timestamp 1676037725
transform 1 0 39008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1676037725
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_423
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_435
timestamp 1676037725
transform 1 0 41124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_447
timestamp 1676037725
transform 1 0 42228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_459
timestamp 1676037725
transform 1 0 43332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_471
timestamp 1676037725
transform 1 0 44436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_227
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1676037725
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_263
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1676037725
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_331
timestamp 1676037725
transform 1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_339
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1676037725
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp 1676037725
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_376
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1676037725
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1676037725
transform 1 0 12512 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 1676037725
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1676037725
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_243
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_275
timestamp 1676037725
transform 1 0 26404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_279
timestamp 1676037725
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_305
timestamp 1676037725
transform 1 0 29164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1676037725
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1676037725
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_351
timestamp 1676037725
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1676037725
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_387
timestamp 1676037725
transform 1 0 36708 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_391
timestamp 1676037725
transform 1 0 37076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_407
timestamp 1676037725
transform 1 0 38548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_411
timestamp 1676037725
transform 1 0 38916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_427
timestamp 1676037725
transform 1 0 40388 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_431
timestamp 1676037725
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_443
timestamp 1676037725
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_455
timestamp 1676037725
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_467
timestamp 1676037725
transform 1 0 44068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1676037725
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1676037725
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_17
timestamp 1676037725
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1676037725
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1676037725
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1676037725
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_183
timestamp 1676037725
transform 1 0 17940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1676037725
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_267
timestamp 1676037725
transform 1 0 25668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_296
timestamp 1676037725
transform 1 0 28336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_299
timestamp 1676037725
transform 1 0 28612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_312
timestamp 1676037725
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_348
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_352
timestamp 1676037725
transform 1 0 33488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1676037725
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1676037725
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_397
timestamp 1676037725
transform 1 0 37628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_409
timestamp 1676037725
transform 1 0 38732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_423
timestamp 1676037725
transform 1 0 40020 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_427
timestamp 1676037725
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_439
timestamp 1676037725
transform 1 0 41492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1676037725
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_192
timestamp 1676037725
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_279
timestamp 1676037725
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_300
timestamp 1676037725
transform 1 0 28704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_320
timestamp 1676037725
transform 1 0 30544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_324
timestamp 1676037725
transform 1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1676037725
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_367
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_375
timestamp 1676037725
transform 1 0 35604 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_406
timestamp 1676037725
transform 1 0 38456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_410
timestamp 1676037725
transform 1 0 38824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_427
timestamp 1676037725
transform 1 0 40388 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_434
timestamp 1676037725
transform 1 0 41032 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_446
timestamp 1676037725
transform 1 0 42136 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_458
timestamp 1676037725
transform 1 0 43240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 1676037725
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_487
timestamp 1676037725
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_499
timestamp 1676037725
transform 1 0 47012 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_507
timestamp 1676037725
transform 1 0 47748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1676037725
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1676037725
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1676037725
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_115
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1676037725
transform 1 0 12144 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_191
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_268
timestamp 1676037725
transform 1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1676037725
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_296
timestamp 1676037725
transform 1 0 28336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_318
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_331
timestamp 1676037725
transform 1 0 31556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1676037725
transform 1 0 33120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_367
timestamp 1676037725
transform 1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_425
timestamp 1676037725
transform 1 0 40204 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1676037725
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1676037725
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_481
timestamp 1676037725
transform 1 0 45356 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1676037725
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1676037725
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1676037725
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1676037725
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_275
timestamp 1676037725
transform 1 0 26404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_279
timestamp 1676037725
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1676037725
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_294
timestamp 1676037725
transform 1 0 28152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_331
timestamp 1676037725
transform 1 0 31556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_335
timestamp 1676037725
transform 1 0 31924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1676037725
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_400
timestamp 1676037725
transform 1 0 37904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_427
timestamp 1676037725
transform 1 0 40388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1676037725
transform 1 0 41032 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_441
timestamp 1676037725
transform 1 0 41676 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_453
timestamp 1676037725
transform 1 0 42780 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_465
timestamp 1676037725
transform 1 0 43884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1676037725
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_485
timestamp 1676037725
transform 1 0 45724 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_490
timestamp 1676037725
transform 1 0 46184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_502
timestamp 1676037725
transform 1 0 47288 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_508
timestamp 1676037725
transform 1 0 47840 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_9
timestamp 1676037725
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1676037725
transform 1 0 2300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1676037725
transform 1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 1676037725
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1676037725
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1676037725
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_150
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1676037725
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1676037725
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_206
timestamp 1676037725
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1676037725
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1676037725
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_277
timestamp 1676037725
transform 1 0 26588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_306
timestamp 1676037725
transform 1 0 29256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_311
timestamp 1676037725
transform 1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_348
timestamp 1676037725
transform 1 0 33120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_356
timestamp 1676037725
transform 1 0 33856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_369
timestamp 1676037725
transform 1 0 35052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_382
timestamp 1676037725
transform 1 0 36248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1676037725
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_426
timestamp 1676037725
transform 1 0 40296 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_430
timestamp 1676037725
transform 1 0 40664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_442
timestamp 1676037725
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_490
timestamp 1676037725
transform 1 0 46184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1676037725
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1676037725
transform 1 0 10580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1676037725
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1676037725
transform 1 0 19504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1676037725
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_256
timestamp 1676037725
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1676037725
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_274
timestamp 1676037725
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_280
timestamp 1676037725
transform 1 0 26864 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_292
timestamp 1676037725
transform 1 0 27968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_295
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1676037725
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1676037725
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_324
timestamp 1676037725
transform 1 0 30912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1676037725
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_359
timestamp 1676037725
transform 1 0 34132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_376
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_382
timestamp 1676037725
transform 1 0 36248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_404
timestamp 1676037725
transform 1 0 38272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_408
timestamp 1676037725
transform 1 0 38640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_416
timestamp 1676037725
transform 1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_440
timestamp 1676037725
transform 1 0 41584 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_452
timestamp 1676037725
transform 1 0 42688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_464
timestamp 1676037725
transform 1 0 43792 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1676037725
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_128
timestamp 1676037725
transform 1 0 12880 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1676037725
transform 1 0 15364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1676037725
transform 1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_183
timestamp 1676037725
transform 1 0 17940 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1676037725
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1676037725
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1676037725
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_359
timestamp 1676037725
transform 1 0 34132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_372
timestamp 1676037725
transform 1 0 35328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_404
timestamp 1676037725
transform 1 0 38272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_408
timestamp 1676037725
transform 1 0 38640 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_413
timestamp 1676037725
transform 1 0 39100 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_425
timestamp 1676037725
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1676037725
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1676037725
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_480
timestamp 1676037725
transform 1 0 45264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1676037725
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1676037725
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_509
timestamp 1676037725
transform 1 0 47932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_512
timestamp 1676037725
transform 1 0 48208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1676037725
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1676037725
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1676037725
transform 1 0 15640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1676037725
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_242
timestamp 1676037725
transform 1 0 23368 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_257
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1676037725
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1676037725
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1676037725
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_346
timestamp 1676037725
transform 1 0 32936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_359
timestamp 1676037725
transform 1 0 34132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_411
timestamp 1676037725
transform 1 0 38916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_425
timestamp 1676037725
transform 1 0 40204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_437
timestamp 1676037725
transform 1 0 41308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_449
timestamp 1676037725
transform 1 0 42412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_461
timestamp 1676037725
transform 1 0 43516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1676037725
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_519
timestamp 1676037725
transform 1 0 48852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1676037725
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_99
timestamp 1676037725
transform 1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_126
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_130
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1676037725
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_229
timestamp 1676037725
transform 1 0 22172 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1676037725
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1676037725
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1676037725
transform 1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_312
timestamp 1676037725
transform 1 0 29808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_325
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_332
timestamp 1676037725
transform 1 0 31648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1676037725
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_387
timestamp 1676037725
transform 1 0 36708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1676037725
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_428
timestamp 1676037725
transform 1 0 40480 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_435
timestamp 1676037725
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_519
timestamp 1676037725
transform 1 0 48852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_61
timestamp 1676037725
transform 1 0 6716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_87
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_99
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_179
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_185
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_191
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_201
timestamp 1676037725
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_217
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1676037725
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_278
timestamp 1676037725
transform 1 0 26680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_284
timestamp 1676037725
transform 1 0 27232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_295
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_315
timestamp 1676037725
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_339
timestamp 1676037725
transform 1 0 32292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_359
timestamp 1676037725
transform 1 0 34132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_387
timestamp 1676037725
transform 1 0 36708 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1676037725
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1676037725
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_443
timestamp 1676037725
transform 1 0 41860 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_447
timestamp 1676037725
transform 1 0 42228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_459
timestamp 1676037725
transform 1 0 43332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1676037725
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_517
timestamp 1676037725
transform 1 0 48668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_520
timestamp 1676037725
transform 1 0 48944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_91
timestamp 1676037725
transform 1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_99
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1676037725
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1676037725
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1676037725
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1676037725
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1676037725
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_248
timestamp 1676037725
transform 1 0 23920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1676037725
transform 1 0 26404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1676037725
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_367
timestamp 1676037725
transform 1 0 34868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_398
timestamp 1676037725
transform 1 0 37720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_402
timestamp 1676037725
transform 1 0 38088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_423
timestamp 1676037725
transform 1 0 40020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_427
timestamp 1676037725
transform 1 0 40388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_437
timestamp 1676037725
transform 1 0 41308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_519
timestamp 1676037725
transform 1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1676037725
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_87
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_95
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1676037725
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_171
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1676037725
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_213
timestamp 1676037725
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_240
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_302
timestamp 1676037725
transform 1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_320
timestamp 1676037725
transform 1 0 30544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1676037725
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_358
timestamp 1676037725
transform 1 0 34040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_378
timestamp 1676037725
transform 1 0 35880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_391
timestamp 1676037725
transform 1 0 37076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_395
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1676037725
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_432
timestamp 1676037725
transform 1 0 40848 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_440
timestamp 1676037725
transform 1 0 41584 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_452
timestamp 1676037725
transform 1 0 42688 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_464
timestamp 1676037725
transform 1 0 43792 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_519
timestamp 1676037725
transform 1 0 48852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1676037725
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1676037725
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1676037725
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1676037725
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1676037725
transform 1 0 18768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1676037725
transform 1 0 20976 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1676037725
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_230
timestamp 1676037725
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_267
timestamp 1676037725
transform 1 0 25668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1676037725
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1676037725
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_308
timestamp 1676037725
transform 1 0 29440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_321
timestamp 1676037725
transform 1 0 30636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1676037725
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1676037725
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_388
timestamp 1676037725
transform 1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_404
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_408
timestamp 1676037725
transform 1 0 38640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_431
timestamp 1676037725
transform 1 0 40756 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_435
timestamp 1676037725
transform 1 0 41124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_513
timestamp 1676037725
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1676037725
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1676037725
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_127
timestamp 1676037725
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1676037725
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_163
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1676037725
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1676037725
transform 1 0 19688 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_232
timestamp 1676037725
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_281
timestamp 1676037725
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_311
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1676037725
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1676037725
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_353
timestamp 1676037725
transform 1 0 33580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_359
timestamp 1676037725
transform 1 0 34132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_370
timestamp 1676037725
transform 1 0 35144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_374
timestamp 1676037725
transform 1 0 35512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_397
timestamp 1676037725
transform 1 0 37628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_410
timestamp 1676037725
transform 1 0 38824 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1676037725
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_427
timestamp 1676037725
transform 1 0 40388 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_437
timestamp 1676037725
transform 1 0 41308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_449
timestamp 1676037725
transform 1 0 42412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_461
timestamp 1676037725
transform 1 0 43516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1676037725
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_519
timestamp 1676037725
transform 1 0 48852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1676037725
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_32
timestamp 1676037725
transform 1 0 4048 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_87
timestamp 1676037725
transform 1 0 9108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1676037725
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1676037725
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1676037725
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_324
timestamp 1676037725
transform 1 0 30912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1676037725
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1676037725
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1676037725
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_377
timestamp 1676037725
transform 1 0 35788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_387
timestamp 1676037725
transform 1 0 36708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_399
timestamp 1676037725
transform 1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_421
timestamp 1676037725
transform 1 0 39836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_425
timestamp 1676037725
transform 1 0 40204 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_436
timestamp 1676037725
transform 1 0 41216 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_513
timestamp 1676037725
transform 1 0 48300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_519
timestamp 1676037725
transform 1 0 48852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1676037725
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 1676037725
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1676037725
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1676037725
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_167
timestamp 1676037725
transform 1 0 16468 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_199
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1676037725
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_288
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_300
timestamp 1676037725
transform 1 0 28704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_328
timestamp 1676037725
transform 1 0 31280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_352
timestamp 1676037725
transform 1 0 33488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_371
timestamp 1676037725
transform 1 0 35236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_395
timestamp 1676037725
transform 1 0 37444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_399
timestamp 1676037725
transform 1 0 37812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_410
timestamp 1676037725
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_443
timestamp 1676037725
transform 1 0 41860 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_447
timestamp 1676037725
transform 1 0 42228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_459
timestamp 1676037725
transform 1 0 43332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1676037725
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_517
timestamp 1676037725
transform 1 0 48668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1676037725
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1676037725
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_116
timestamp 1676037725
transform 1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1676037725
transform 1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1676037725
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1676037725
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1676037725
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_242
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_263
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_267
timestamp 1676037725
transform 1 0 25668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1676037725
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1676037725
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_310
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_314
timestamp 1676037725
transform 1 0 29992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_320
timestamp 1676037725
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1676037725
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1676037725
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1676037725
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_397
timestamp 1676037725
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1676037725
transform 1 0 39744 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_433
timestamp 1676037725
transform 1 0 40940 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_439
timestamp 1676037725
transform 1 0 41492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_513
timestamp 1676037725
transform 1 0 48300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_519
timestamp 1676037725
transform 1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1676037725
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1676037725
transform 1 0 7268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1676037725
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1676037725
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1676037725
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1676037725
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_231
timestamp 1676037725
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_239
timestamp 1676037725
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1676037725
transform 1 0 24840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1676037725
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_288
timestamp 1676037725
transform 1 0 27600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_305
timestamp 1676037725
transform 1 0 29164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_346
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_350
timestamp 1676037725
transform 1 0 33304 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_360
timestamp 1676037725
transform 1 0 34224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1676037725
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_397
timestamp 1676037725
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_408
timestamp 1676037725
transform 1 0 38640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_414
timestamp 1676037725
transform 1 0 39192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_432
timestamp 1676037725
transform 1 0 40848 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_438
timestamp 1676037725
transform 1 0 41400 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_450
timestamp 1676037725
transform 1 0 42504 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_462
timestamp 1676037725
transform 1 0 43608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1676037725
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_519
timestamp 1676037725
transform 1 0 48852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1676037725
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_83
timestamp 1676037725
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1676037725
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1676037725
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1676037725
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1676037725
transform 1 0 12788 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_199
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1676037725
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_274
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1676037725
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_330
timestamp 1676037725
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_359
timestamp 1676037725
transform 1 0 34132 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_372
timestamp 1676037725
transform 1 0 35328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_378
timestamp 1676037725
transform 1 0 35880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1676037725
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_395
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_418
timestamp 1676037725
transform 1 0 39560 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_431
timestamp 1676037725
transform 1 0 40756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_438
timestamp 1676037725
transform 1 0 41400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1676037725
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_512
timestamp 1676037725
transform 1 0 48208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 1676037725
transform 1 0 8096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1676037725
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_91
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1676037725
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_112
timestamp 1676037725
transform 1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_120
timestamp 1676037725
transform 1 0 12144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_130
timestamp 1676037725
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_203
timestamp 1676037725
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1676037725
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_238
timestamp 1676037725
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_246
timestamp 1676037725
transform 1 0 23736 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_258
timestamp 1676037725
transform 1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_276
timestamp 1676037725
transform 1 0 26496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_282
timestamp 1676037725
transform 1 0 27048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_287
timestamp 1676037725
transform 1 0 27508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1676037725
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_314
timestamp 1676037725
transform 1 0 29992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_320
timestamp 1676037725
transform 1 0 30544 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_332
timestamp 1676037725
transform 1 0 31648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_336
timestamp 1676037725
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_340
timestamp 1676037725
transform 1 0 32384 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_387
timestamp 1676037725
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_395
timestamp 1676037725
transform 1 0 37444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1676037725
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1676037725
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_455
timestamp 1676037725
transform 1 0 42964 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_467
timestamp 1676037725
transform 1 0 44068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_505
timestamp 1676037725
transform 1 0 47564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_510
timestamp 1676037725
transform 1 0 48024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_517
timestamp 1676037725
transform 1 0 48668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1676037725
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1676037725
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_101
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1676037725
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1676037725
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1676037725
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_138
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1676037725
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1676037725
transform 1 0 17204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1676037725
transform 1 0 22264 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_266
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_272
timestamp 1676037725
transform 1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1676037725
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1676037725
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_331
timestamp 1676037725
transform 1 0 31556 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_345
timestamp 1676037725
transform 1 0 32844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_358
timestamp 1676037725
transform 1 0 34040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_371
timestamp 1676037725
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_375
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_399
timestamp 1676037725
transform 1 0 37812 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_421
timestamp 1676037725
transform 1 0 39836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_431
timestamp 1676037725
transform 1 0 40756 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_434
timestamp 1676037725
transform 1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_455
timestamp 1676037725
transform 1 0 42964 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_493
timestamp 1676037725
transform 1 0 46460 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1676037725
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_510
timestamp 1676037725
transform 1 0 48024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1676037725
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1676037725
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_103
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_107
timestamp 1676037725
transform 1 0 10948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1676037725
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_243
timestamp 1676037725
transform 1 0 23460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_268
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_279
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1676037725
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_314
timestamp 1676037725
transform 1 0 29992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_320
timestamp 1676037725
transform 1 0 30544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1676037725
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_356
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_376
timestamp 1676037725
transform 1 0 35696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_414
timestamp 1676037725
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_423
timestamp 1676037725
transform 1 0 40020 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_434
timestamp 1676037725
transform 1 0 41032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_447
timestamp 1676037725
transform 1 0 42228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_454
timestamp 1676037725
transform 1 0 42872 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_462
timestamp 1676037725
transform 1 0 43608 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_474
timestamp 1676037725
transform 1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_485
timestamp 1676037725
transform 1 0 45724 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_490
timestamp 1676037725
transform 1 0 46184 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_495
timestamp 1676037725
transform 1 0 46644 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_502
timestamp 1676037725
transform 1 0 47288 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_508
timestamp 1676037725
transform 1 0 47840 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_514
timestamp 1676037725
transform 1 0 48392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_519
timestamp 1676037725
transform 1 0 48852 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_29
timestamp 1676037725
transform 1 0 3772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_67
timestamp 1676037725
transform 1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_85
timestamp 1676037725
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1676037725
transform 1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_141
timestamp 1676037725
transform 1 0 14076 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1676037725
transform 1 0 19228 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_256
timestamp 1676037725
transform 1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_286
timestamp 1676037725
transform 1 0 27416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_290
timestamp 1676037725
transform 1 0 27784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1676037725
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1676037725
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_348
timestamp 1676037725
transform 1 0 33120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_352
timestamp 1676037725
transform 1 0 33488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_378
timestamp 1676037725
transform 1 0 35880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1676037725
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_415
timestamp 1676037725
transform 1 0 39284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_421
timestamp 1676037725
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_432
timestamp 1676037725
transform 1 0 40848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_439
timestamp 1676037725
transform 1 0 41492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1676037725
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_465
timestamp 1676037725
transform 1 0 43884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_472
timestamp 1676037725
transform 1 0 44528 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_479
timestamp 1676037725
transform 1 0 45172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_486
timestamp 1676037725
transform 1 0 45816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_493
timestamp 1676037725
transform 1 0 46460 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1676037725
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1676037725
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_98
timestamp 1676037725
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1676037725
transform 1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_199
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1676037725
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1676037725
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1676037725
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_259
timestamp 1676037725
transform 1 0 24932 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1676037725
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_300
timestamp 1676037725
transform 1 0 28704 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_320
timestamp 1676037725
transform 1 0 30544 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_324
timestamp 1676037725
transform 1 0 30912 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_327
timestamp 1676037725
transform 1 0 31188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_350
timestamp 1676037725
transform 1 0 33304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_367
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_432
timestamp 1676037725
transform 1 0 40848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_436
timestamp 1676037725
transform 1 0 41216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_462
timestamp 1676037725
transform 1 0 43608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1676037725
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_483
timestamp 1676037725
transform 1 0 45540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_487
timestamp 1676037725
transform 1 0 45908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_492
timestamp 1676037725
transform 1 0 46368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_500
timestamp 1676037725
transform 1 0 47104 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_508
timestamp 1676037725
transform 1 0 47840 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_520
timestamp 1676037725
transform 1 0 48944 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_524
timestamp 1676037725
transform 1 0 49312 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_63
timestamp 1676037725
transform 1 0 6900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_256
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1676037725
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_300
timestamp 1676037725
transform 1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_307
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_311
timestamp 1676037725
transform 1 0 29716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_348
timestamp 1676037725
transform 1 0 33120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_352
timestamp 1676037725
transform 1 0 33488 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_377
timestamp 1676037725
transform 1 0 35788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_387
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_404
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_408
timestamp 1676037725
transform 1 0 38640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_419
timestamp 1676037725
transform 1 0 39652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_426
timestamp 1676037725
transform 1 0 40296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_453
timestamp 1676037725
transform 1 0 42780 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_476
timestamp 1676037725
transform 1 0 44896 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_488
timestamp 1676037725
transform 1 0 46000 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_496
timestamp 1676037725
transform 1 0 46736 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_509
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_519
timestamp 1676037725
transform 1 0 48852 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1676037725
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_272
timestamp 1676037725
transform 1 0 26128 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_287
timestamp 1676037725
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1676037725
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1676037725
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_349
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1676037725
transform 1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1676037725
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_411
timestamp 1676037725
transform 1 0 38916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1676037725
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_432
timestamp 1676037725
transform 1 0 40848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_436
timestamp 1676037725
transform 1 0 41216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_446
timestamp 1676037725
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_459
timestamp 1676037725
transform 1 0 43332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_466
timestamp 1676037725
transform 1 0 43976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_473
timestamp 1676037725
transform 1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_487
timestamp 1676037725
transform 1 0 45908 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_502
timestamp 1676037725
transform 1 0 47288 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_518
timestamp 1676037725
transform 1 0 48760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 42136 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold2
timestamp 1676037725
transform -1 0 44896 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform -1 0 43332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 44712 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 48208 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform -1 0 46000 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1676037725
transform 1 0 12328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1676037725
transform -1 0 47288 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1676037725
transform -1 0 48852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1676037725
transform -1 0 10764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform -1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 47012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform -1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1676037725
transform -1 0 2484 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform -1 0 2484 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform -1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform -1 0 2484 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform -1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform -1 0 2484 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform -1 0 2484 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1676037725
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 48392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1676037725
transform -1 0 49404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform -1 0 49404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 48392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform -1 0 49404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform -1 0 49404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform -1 0 49404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 48392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform -1 0 49404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform -1 0 49404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform -1 0 49404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform -1 0 49404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 48392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform -1 0 49404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform -1 0 48668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform -1 0 47840 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 46368 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 46184 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform -1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 47748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 47012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 49128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform -1 0 49404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform -1 0 49404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 49128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform -1 0 49404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform -1 0 49404 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform -1 0 49404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 48392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform -1 0 49404 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform -1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform -1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform -1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 38640 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1676037725
transform 1 0 33672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 39284 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1676037725
transform 1 0 43700 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1676037725
transform 1 0 40020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1676037725
transform 1 0 44344 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1676037725
transform -1 0 11960 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1676037725
transform 1 0 41216 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1676037725
transform 1 0 40664 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1676037725
transform 1 0 42596 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1676037725
transform 1 0 43792 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 42596 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 41216 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1676037725
transform 1 0 43240 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 41860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 45540 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 44896 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1676037725
transform -1 0 12696 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1676037725
transform -1 0 22908 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform -1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1676037725
transform -1 0 30636 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1676037725
transform -1 0 24104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1676037725
transform -1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform -1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1676037725
transform -1 0 28796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1676037725
transform -1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform -1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1676037725
transform -1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform -1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1676037725
transform -1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1676037725
transform -1 0 47104 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform -1 0 47288 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1676037725
transform -1 0 48392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1676037725
transform -1 0 46368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1676037725
transform -1 0 44528 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform -1 0 45540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform -1 0 4876 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform -1 0 3036 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform -1 0 3036 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform -1 0 3036 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform -1 0 3036 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform -1 0 3036 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform -1 0 3036 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform -1 0 3036 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform -1 0 4876 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform -1 0 3036 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform -1 0 3036 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform -1 0 3036 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform -1 0 3036 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform -1 0 5428 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform -1 0 5428 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform -1 0 7268 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform -1 0 7268 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform -1 0 5428 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform -1 0 7268 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform -1 0 3036 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform -1 0 3036 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform -1 0 3036 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform -1 0 3036 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform -1 0 3036 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform -1 0 3036 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform -1 0 3036 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform -1 0 3036 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 45816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 43976 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 45816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 45816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 45816 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform -1 0 5428 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform -1 0 9384 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform -1 0 11224 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform -1 0 11224 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform -1 0 11960 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform -1 0 11224 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform -1 0 14076 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform -1 0 13800 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform -1 0 13800 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform -1 0 4876 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform -1 0 16376 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform -1 0 16744 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform -1 0 16376 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform -1 0 18860 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform -1 0 16376 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform -1 0 18400 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform -1 0 18952 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform -1 0 21528 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform -1 0 3496 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform -1 0 4232 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform -1 0 6072 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform -1 0 13248 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform -1 0 15732 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform -1 0 18308 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform -1 0 19596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 22356 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 29256 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 26404 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 24472 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 24104 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22356 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 18952 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 23828 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22816 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 20976 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21528 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 18952 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22172 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 20608 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23828 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 25300 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 28888 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 27416 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 29900 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 26680 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25668 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 26680 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 23000 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 30452 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32200 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 36984 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 35144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 37812 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33856 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 35696 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32108 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 32936 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27968 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 30360 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 28796 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 32200 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31096 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 32568 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 29348 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26864 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 43608 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30820 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 31832 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31372 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33672 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 35420 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35052 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 36708 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 34132 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32476 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 39284 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39100 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 39192 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37996 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39468 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 39560 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 37628 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33580 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35604 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 39744 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 41860 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 40756 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39560 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 38180 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39560 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 38916 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 34132 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 31188 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 27416 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 26680 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 25668 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 26404 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 25300 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 24104 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23828 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21528 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 21252 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21252 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22080 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22264 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18676 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 14904 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16100 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 14536 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 13524 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 12420 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16100 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 17020 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 18952 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27232 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1676037725
transform -1 0 23460 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__258
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1676037725
transform -1 0 21712 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1676037725
transform -1 0 23920 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__211
timestamp 1676037725
transform -1 0 15732 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1676037725
transform -1 0 17572 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__214
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1676037725
transform -1 0 20332 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1676037725
transform -1 0 20516 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__216
timestamp 1676037725
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19872 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27968 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__259
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__260
timestamp 1676037725
transform -1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27876 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__261
timestamp 1676037725
transform -1 0 17112 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__262
timestamp 1676037725
transform -1 0 22908 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__212
timestamp 1676037725
transform 1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1676037725
transform -1 0 24104 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__213
timestamp 1676037725
transform -1 0 27968 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__215
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19964 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform -1 0 30268 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 33304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1676037725
transform -1 0 28612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform -1 0 31832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__217
timestamp 1676037725
transform -1 0 30084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31740 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform -1 0 34316 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 39560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform -1 0 34040 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33120 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform -1 0 30544 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform -1 0 36708 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform -1 0 34316 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform -1 0 38824 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1676037725
transform -1 0 30544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform -1 0 36800 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform -1 0 36524 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__224
timestamp 1676037725
transform -1 0 31832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform -1 0 38272 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform -1 0 36248 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__227
timestamp 1676037725
transform 1 0 33764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1676037725
transform -1 0 33120 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform -1 0 36708 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38640 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform -1 0 39100 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform -1 0 34224 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1676037725
transform -1 0 34132 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1676037725
transform -1 0 31832 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__218
timestamp 1676037725
transform -1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform -1 0 35328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform -1 0 36892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform -1 0 38272 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform -1 0 33120 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1676037725
transform -1 0 27968 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform -1 0 34132 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform -1 0 33120 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__219
timestamp 1676037725
transform -1 0 29992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform -1 0 37904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1676037725
transform -1 0 30636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1676037725
transform -1 0 27968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform -1 0 31372 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform -1 0 29256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform -1 0 34316 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 38456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform -1 0 30544 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 30176 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1676037725
transform -1 0 26496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform -1 0 30544 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31004 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__222
timestamp 1676037725
transform -1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1676037725
transform -1 0 33396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 37904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform -1 0 32108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1676037725
transform -1 0 32936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform -1 0 33120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__223
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 39192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform -1 0 30544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__225
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform -1 0 28980 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform -1 0 33396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 37720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform -1 0 29440 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1676037725
transform -1 0 27784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__226
timestamp 1676037725
transform -1 0 26680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform -1 0 33120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 36800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38824 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform -1 0 24104 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__228
timestamp 1676037725
transform 1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 28428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 29164 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform -1 0 31740 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33028 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__234
timestamp 1676037725
transform -1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35696 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__244
timestamp 1676037725
transform 1 0 31280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform -1 0 30912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40204 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41400 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform -1 0 33488 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__252
timestamp 1676037725
transform -1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform -1 0 38272 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41216 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1676037725
transform -1 0 34316 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform -1 0 36892 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__253
timestamp 1676037725
transform 1 0 41124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36064 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35512 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40112 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31740 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 31464 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform -1 0 40848 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__230
timestamp 1676037725
transform -1 0 35144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform -1 0 40756 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1676037725
transform -1 0 35512 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform -1 0 40848 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 37076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1676037725
transform -1 0 35696 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform -1 0 38640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31556 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 25760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27324 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__235
timestamp 1676037725
transform -1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform -1 0 25668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__236
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1676037725
transform -1 0 22908 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__237
timestamp 1676037725
transform -1 0 20056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__238
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24196 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__239
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__240
timestamp 1676037725
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 12604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__242
timestamp 1676037725
transform -1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__243
timestamp 1676037725
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__245
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__246
timestamp 1676037725
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__247
timestamp 1676037725
transform -1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__248
timestamp 1676037725
transform -1 0 9936 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__249
timestamp 1676037725
transform -1 0 10764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__250
timestamp 1676037725
transform -1 0 10120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__251
timestamp 1676037725
transform -1 0 10120 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 26200 49294 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 26200 1638 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 13608 51000 13728 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 17688 51000 17808 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 18096 51000 18216 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 18912 51000 19032 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 19320 51000 19440 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 19728 51000 19848 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 20136 51000 20256 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 21360 51000 21480 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 14016 51000 14136 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 21768 51000 21888 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 22176 51000 22296 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 22992 51000 23112 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 23400 51000 23520 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 24216 51000 24336 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 25032 51000 25152 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 25440 51000 25560 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 14832 51000 14952 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 15240 51000 15360 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 15648 51000 15768 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 16056 51000 16176 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 16872 51000 16992 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 17280 51000 17400 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 1368 51000 1488 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 5448 51000 5568 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 5856 51000 5976 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 6672 51000 6792 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 7080 51000 7200 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 7488 51000 7608 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 7896 51000 8016 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 8712 51000 8832 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 9120 51000 9240 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 1776 51000 1896 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 9528 51000 9648 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 9936 51000 10056 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 10752 51000 10872 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 11160 51000 11280 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 11568 51000 11688 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 11976 51000 12096 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 12792 51000 12912 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 13200 51000 13320 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 2184 51000 2304 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 2592 51000 2712 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 3000 51000 3120 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 3408 51000 3528 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 3816 51000 3936 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 4632 51000 4752 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 5040 51000 5160 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 test_enable
port 206 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal1 21850 4658 21850 4658 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 19872 4658 19872 4658 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 18906 6596 18906 6596 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 16284 6222 16284 6222 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20424 20978 20424 20978 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal2 18630 9044 18630 9044 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 16284 15538 16284 15538 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 16790 13498 16790 13498 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 16100 9146 16100 9146 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 15226 9010 15226 9010 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 12650 12954 12650 12954 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 15640 13838 15640 13838 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 14122 9894 14122 9894 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 11040 11186 11040 11186 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 18124 14450 18124 14450 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 14950 13056 14950 13056 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 12926 11696 12926 11696 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 14674 14926 14674 14926 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 16146 14892 16146 14892 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 13018 16014 13018 16014 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal2 15502 14892 15502 14892 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17848 7786 17848 7786 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 19642 7276 19642 7276 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 15594 14314 15594 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17618 14994 17618 14994 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17526 14450 17526 14450 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16882 10098 16882 10098 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15916 11186 15916 11186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16882 14042 16882 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 16974 8908 16974 8908 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 17066 9146 17066 9146 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 17710 7854 17710 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 12972 15470 12972 15470 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15594 9690 15594 9690 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 16836 6766 16836 6766 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13432 15470 13432 15470 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17802 13974 17802 13974 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15962 13974 15962 13974 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14536 10098 14536 10098 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 13616 12852 13616 12852 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15410 14042 15410 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 14260 10234 14260 10234 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 16560 10778 16560 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 15502 10302 15502 10302 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 9706 15810 9706 15810 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12374 10540 12374 10540 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15272 7854 15272 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 9798 15538 9798 15538 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 14586 18308 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14582 14586 14582 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15824 10710 15824 10710 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12006 13906 12006 13906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12144 12954 12144 12954 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 14398 11186 14398 11186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 12742 12274 12742 12274 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 12512 12614 12512 12614 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13570 16014 13570 16014 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 14586 12926 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 12466 14586 12466 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14214 15878 14214 15878 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 14926 15870 14926 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17158 15130 17158 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14858 11356 14858 11356 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12834 16218 12834 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15088 15130 15088 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 13708 14246 13708 14246 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 14214 14314 14214 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11684 16218 11684 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 20332 3434 20332 3434 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 20194 3060 20194 3060 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 26312 3026 26312 3026 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 28842 4012 28842 4012 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 23506 2856 23506 2856 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 19113 2414 19113 2414 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 21298 3740 21298 3740 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 23161 4114 23161 4114 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 27600 2958 27600 2958 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 19090 4080 19090 4080 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 20654 4012 20654 4012 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 25898 4318 25898 4318 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 16606 3740 16606 3740 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 19090 6086 19090 6086 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 24564 3570 24564 3570 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9568 3026 9568 3026 0 ccff_head
rlabel metal2 49358 24259 49358 24259 0 ccff_head_1
rlabel metal2 41354 1622 41354 1622 0 ccff_tail
rlabel metal2 1610 24524 1610 24524 0 ccff_tail_0
rlabel metal1 2990 2414 2990 2414 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6290 1472 6290 0 chanx_left_in[11]
rlabel metal1 1840 6766 1840 6766 0 chanx_left_in[12]
rlabel metal1 1472 6698 1472 6698 0 chanx_left_in[13]
rlabel metal1 1472 7378 1472 7378 0 chanx_left_in[14]
rlabel metal1 1472 7854 1472 7854 0 chanx_left_in[15]
rlabel metal1 1748 8058 1748 8058 0 chanx_left_in[16]
rlabel metal1 1794 8942 1794 8942 0 chanx_left_in[17]
rlabel metal1 1518 8874 1518 8874 0 chanx_left_in[18]
rlabel metal1 1472 9554 1472 9554 0 chanx_left_in[19]
rlabel metal1 1840 2346 1840 2346 0 chanx_left_in[1]
rlabel metal1 1748 9690 1748 9690 0 chanx_left_in[20]
rlabel metal1 2346 10676 2346 10676 0 chanx_left_in[21]
rlabel metal1 1472 10642 1472 10642 0 chanx_left_in[22]
rlabel metal2 1610 11033 1610 11033 0 chanx_left_in[23]
rlabel metal1 2346 11696 2346 11696 0 chanx_left_in[24]
rlabel metal1 1886 12274 1886 12274 0 chanx_left_in[25]
rlabel metal1 1426 11730 1426 11730 0 chanx_left_in[26]
rlabel metal2 1242 12699 1242 12699 0 chanx_left_in[27]
rlabel metal1 1518 12886 1518 12886 0 chanx_left_in[28]
rlabel metal2 3542 13651 3542 13651 0 chanx_left_in[29]
rlabel metal1 2208 2414 2208 2414 0 chanx_left_in[2]
rlabel metal1 1472 3026 1472 3026 0 chanx_left_in[3]
rlabel metal1 1748 3162 1748 3162 0 chanx_left_in[4]
rlabel metal1 1840 4114 1840 4114 0 chanx_left_in[5]
rlabel metal1 1564 4182 1564 4182 0 chanx_left_in[6]
rlabel metal1 1472 4590 1472 4590 0 chanx_left_in[7]
rlabel metal1 1748 4794 1748 4794 0 chanx_left_in[8]
rlabel metal2 2806 5457 2806 5457 0 chanx_left_in[9]
rlabel metal3 1234 13804 1234 13804 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal3 1234 18292 1234 18292 0 chanx_left_out[11]
rlabel metal3 1096 18700 1096 18700 0 chanx_left_out[12]
rlabel metal1 2645 20366 2645 20366 0 chanx_left_out[13]
rlabel metal2 2898 20247 2898 20247 0 chanx_left_out[14]
rlabel metal3 1234 19924 1234 19924 0 chanx_left_out[15]
rlabel metal3 1004 20332 1004 20332 0 chanx_left_out[16]
rlabel metal3 866 20740 866 20740 0 chanx_left_out[17]
rlabel metal3 1740 21148 1740 21148 0 chanx_left_out[18]
rlabel metal3 1234 21556 1234 21556 0 chanx_left_out[19]
rlabel metal3 866 14212 866 14212 0 chanx_left_out[1]
rlabel via2 3266 21947 3266 21947 0 chanx_left_out[20]
rlabel metal3 1395 22372 1395 22372 0 chanx_left_out[21]
rlabel metal2 4002 22457 4002 22457 0 chanx_left_out[22]
rlabel metal2 2990 22797 2990 22797 0 chanx_left_out[23]
rlabel metal1 6440 21454 6440 21454 0 chanx_left_out[24]
rlabel metal1 3864 18802 3864 18802 0 chanx_left_out[25]
rlabel metal1 5888 19890 5888 19890 0 chanx_left_out[26]
rlabel metal1 6486 20366 6486 20366 0 chanx_left_out[27]
rlabel metal1 6348 21318 6348 21318 0 chanx_left_out[28]
rlabel metal2 3174 25551 3174 25551 0 chanx_left_out[29]
rlabel metal3 820 14620 820 14620 0 chanx_left_out[2]
rlabel metal3 820 15028 820 15028 0 chanx_left_out[3]
rlabel metal3 820 15436 820 15436 0 chanx_left_out[4]
rlabel metal3 866 15844 866 15844 0 chanx_left_out[5]
rlabel metal3 866 16252 866 16252 0 chanx_left_out[6]
rlabel metal3 820 16660 820 16660 0 chanx_left_out[7]
rlabel metal3 866 17068 866 17068 0 chanx_left_out[8]
rlabel metal3 1234 17476 1234 17476 0 chanx_left_out[9]
rlabel metal1 48438 13906 48438 13906 0 chanx_right_in_0[0]
rlabel metal2 49358 18003 49358 18003 0 chanx_right_in_0[10]
rlabel metal1 49404 18734 49404 18734 0 chanx_right_in_0[11]
rlabel metal2 48806 18479 48806 18479 0 chanx_right_in_0[12]
rlabel metal2 49266 19159 49266 19159 0 chanx_right_in_0[13]
rlabel metal1 49312 19754 49312 19754 0 chanx_right_in_0[14]
rlabel metal1 49404 20434 49404 20434 0 chanx_right_in_0[15]
rlabel metal2 48806 20111 48806 20111 0 chanx_right_in_0[16]
rlabel metal2 49358 20757 49358 20757 0 chanx_right_in_0[17]
rlabel metal1 49404 22950 49404 22950 0 chanx_right_in_0[18]
rlabel metal2 49266 21675 49266 21675 0 chanx_right_in_0[19]
rlabel metal2 49266 14025 49266 14025 0 chanx_right_in_0[1]
rlabel via2 48806 21845 48806 21845 0 chanx_right_in_0[20]
rlabel metal1 49358 22576 49358 22576 0 chanx_right_in_0[21]
rlabel metal3 49274 22644 49274 22644 0 chanx_right_in_0[22]
rlabel metal1 47794 23052 47794 23052 0 chanx_right_in_0[23]
rlabel metal2 47610 22831 47610 22831 0 chanx_right_in_0[24]
rlabel metal1 47748 22746 47748 22746 0 chanx_right_in_0[25]
rlabel metal2 49266 23783 49266 23783 0 chanx_right_in_0[26]
rlabel metal3 47380 23596 47380 23596 0 chanx_right_in_0[27]
rlabel metal3 48906 25092 48906 25092 0 chanx_right_in_0[28]
rlabel metal1 49220 24174 49220 24174 0 chanx_right_in_0[29]
rlabel metal2 49266 14433 49266 14433 0 chanx_right_in_0[2]
rlabel metal2 49358 14943 49358 14943 0 chanx_right_in_0[3]
rlabel metal2 49358 15385 49358 15385 0 chanx_right_in_0[4]
rlabel metal2 49358 15895 49358 15895 0 chanx_right_in_0[5]
rlabel metal1 49404 16558 49404 16558 0 chanx_right_in_0[6]
rlabel metal1 49312 17170 49312 17170 0 chanx_right_in_0[7]
rlabel metal2 48806 16847 48806 16847 0 chanx_right_in_0[8]
rlabel metal2 49358 17493 49358 17493 0 chanx_right_in_0[9]
rlabel metal2 46690 2737 46690 2737 0 chanx_right_out_0[0]
rlabel metal1 49312 4658 49312 4658 0 chanx_right_out_0[10]
rlabel metal2 49174 5593 49174 5593 0 chanx_right_out_0[11]
rlabel metal3 49504 6324 49504 6324 0 chanx_right_out_0[12]
rlabel metal1 49220 5746 49220 5746 0 chanx_right_out_0[13]
rlabel metal1 49312 6358 49312 6358 0 chanx_right_out_0[14]
rlabel metal3 49734 7548 49734 7548 0 chanx_right_out_0[15]
rlabel metal2 46874 8177 46874 8177 0 chanx_right_out_0[16]
rlabel metal1 49266 7446 49266 7446 0 chanx_right_out_0[17]
rlabel metal1 49220 7922 49220 7922 0 chanx_right_out_0[18]
rlabel metal2 49174 8857 49174 8857 0 chanx_right_out_0[19]
rlabel metal2 46782 2397 46782 2397 0 chanx_right_out_0[1]
rlabel metal3 48814 9588 48814 9588 0 chanx_right_out_0[20]
rlabel metal1 49266 9010 49266 9010 0 chanx_right_out_0[21]
rlabel metal1 49220 9622 49220 9622 0 chanx_right_out_0[22]
rlabel metal2 49174 10455 49174 10455 0 chanx_right_out_0[23]
rlabel metal1 49220 10710 49220 10710 0 chanx_right_out_0[24]
rlabel metal2 49174 11407 49174 11407 0 chanx_right_out_0[25]
rlabel metal2 49174 11917 49174 11917 0 chanx_right_out_0[26]
rlabel metal3 49734 12444 49734 12444 0 chanx_right_out_0[27]
rlabel via2 49174 12835 49174 12835 0 chanx_right_out_0[28]
rlabel metal3 49734 13260 49734 13260 0 chanx_right_out_0[29]
rlabel metal3 49412 2244 49412 2244 0 chanx_right_out_0[2]
rlabel metal2 46874 2805 46874 2805 0 chanx_right_out_0[3]
rlabel metal3 49504 3060 49504 3060 0 chanx_right_out_0[4]
rlabel metal2 49174 2975 49174 2975 0 chanx_right_out_0[5]
rlabel metal1 49220 3094 49220 3094 0 chanx_right_out_0[6]
rlabel metal2 49174 3927 49174 3927 0 chanx_right_out_0[7]
rlabel metal1 47610 5134 47610 5134 0 chanx_right_out_0[8]
rlabel metal1 49266 4114 49266 4114 0 chanx_right_out_0[9]
rlabel metal2 26082 21471 26082 21471 0 chany_top_in[0]
rlabel metal1 29118 23664 29118 23664 0 chany_top_in[10]
rlabel metal2 28658 25306 28658 25306 0 chany_top_in[11]
rlabel metal2 32522 24378 32522 24378 0 chany_top_in[12]
rlabel metal1 33028 24174 33028 24174 0 chany_top_in[13]
rlabel metal2 33258 23239 33258 23239 0 chany_top_in[14]
rlabel metal1 33488 23086 33488 23086 0 chany_top_in[15]
rlabel metal1 39468 24174 39468 24174 0 chany_top_in[16]
rlabel metal1 43930 24140 43930 24140 0 chany_top_in[17]
rlabel metal2 33166 25442 33166 25442 0 chany_top_in[18]
rlabel metal2 44574 24378 44574 24378 0 chany_top_in[19]
rlabel metal1 16974 22440 16974 22440 0 chany_top_in[1]
rlabel metal1 40940 21590 40940 21590 0 chany_top_in[20]
rlabel metal2 40710 21563 40710 21563 0 chany_top_in[21]
rlabel via2 42642 22627 42642 22627 0 chany_top_in[22]
rlabel metal1 37398 21930 37398 21930 0 chany_top_in[23]
rlabel metal3 42205 22100 42205 22100 0 chany_top_in[24]
rlabel metal2 37858 24633 37858 24633 0 chany_top_in[25]
rlabel metal1 39008 21658 39008 21658 0 chany_top_in[26]
rlabel metal1 42090 22542 42090 22542 0 chany_top_in[27]
rlabel metal2 45770 23800 45770 23800 0 chany_top_in[28]
rlabel metal1 44344 22610 44344 22610 0 chany_top_in[29]
rlabel metal1 16698 23290 16698 23290 0 chany_top_in[2]
rlabel metal1 22862 23562 22862 23562 0 chany_top_in[3]
rlabel metal1 24104 21114 24104 21114 0 chany_top_in[4]
rlabel metal2 30406 24378 30406 24378 0 chany_top_in[5]
rlabel metal2 25254 24769 25254 24769 0 chany_top_in[6]
rlabel metal1 27094 24174 27094 24174 0 chany_top_in[7]
rlabel metal2 27830 23868 27830 23868 0 chany_top_in[8]
rlabel metal1 28566 24208 28566 24208 0 chany_top_in[9]
rlabel metal2 2254 24252 2254 24252 0 chany_top_out[0]
rlabel metal1 8464 24242 8464 24242 0 chany_top_out[10]
rlabel metal1 9062 23630 9062 23630 0 chany_top_out[11]
rlabel metal2 9982 24490 9982 24490 0 chany_top_out[12]
rlabel metal2 10626 24966 10626 24966 0 chany_top_out[13]
rlabel metal2 11270 24728 11270 24728 0 chany_top_out[14]
rlabel metal1 11270 24242 11270 24242 0 chany_top_out[15]
rlabel metal2 12703 26316 12703 26316 0 chany_top_out[16]
rlabel metal1 13340 23154 13340 23154 0 chany_top_out[17]
rlabel metal1 13570 24242 13570 24242 0 chany_top_out[18]
rlabel metal1 14352 23766 14352 23766 0 chany_top_out[19]
rlabel metal1 3496 21590 3496 21590 0 chany_top_out[1]
rlabel metal2 15134 24490 15134 24490 0 chany_top_out[20]
rlabel metal2 15778 24728 15778 24728 0 chany_top_out[21]
rlabel metal1 16146 23630 16146 23630 0 chany_top_out[22]
rlabel metal1 17342 22134 17342 22134 0 chany_top_out[23]
rlabel metal1 16790 24242 16790 24242 0 chany_top_out[24]
rlabel metal1 18124 23630 18124 23630 0 chany_top_out[25]
rlabel metal1 19688 21930 19688 21930 0 chany_top_out[26]
rlabel metal1 18998 24242 18998 24242 0 chany_top_out[27]
rlabel metal2 20286 24796 20286 24796 0 chany_top_out[28]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[29]
rlabel metal1 3266 24242 3266 24242 0 chany_top_out[2]
rlabel metal1 3956 23630 3956 23630 0 chany_top_out[3]
rlabel metal2 4830 24490 4830 24490 0 chany_top_out[4]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[5]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[6]
rlabel metal1 6302 24242 6302 24242 0 chany_top_out[7]
rlabel metal1 7682 22542 7682 22542 0 chany_top_out[8]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[9]
rlabel metal1 18400 12818 18400 12818 0 clknet_0_prog_clk
rlabel metal1 13662 8534 13662 8534 0 clknet_4_0_0_prog_clk
rlabel metal2 32154 11152 32154 11152 0 clknet_4_10_0_prog_clk
rlabel metal1 37628 11186 37628 11186 0 clknet_4_11_0_prog_clk
rlabel metal1 32338 17238 32338 17238 0 clknet_4_12_0_prog_clk
rlabel metal2 34086 19584 34086 19584 0 clknet_4_13_0_prog_clk
rlabel metal1 34868 15538 34868 15538 0 clknet_4_14_0_prog_clk
rlabel metal1 39330 22066 39330 22066 0 clknet_4_15_0_prog_clk
rlabel metal1 18860 12886 18860 12886 0 clknet_4_1_0_prog_clk
rlabel metal2 21022 3230 21022 3230 0 clknet_4_2_0_prog_clk
rlabel metal1 25622 12886 25622 12886 0 clknet_4_3_0_prog_clk
rlabel metal1 14490 19380 14490 19380 0 clknet_4_4_0_prog_clk
rlabel metal2 21114 14654 21114 14654 0 clknet_4_5_0_prog_clk
rlabel metal2 22770 16898 22770 16898 0 clknet_4_6_0_prog_clk
rlabel metal1 25484 19346 25484 19346 0 clknet_4_7_0_prog_clk
rlabel metal2 28842 5712 28842 5712 0 clknet_4_8_0_prog_clk
rlabel metal2 31142 14722 31142 14722 0 clknet_4_9_0_prog_clk
rlabel metal2 11730 1554 11730 1554 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 13846 1554 13846 1554 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 15962 1554 15962 1554 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 18078 823 18078 823 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 29118 2414 29118 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[1]
rlabel metal2 33166 1989 33166 1989 0 gfpga_pad_io_soc_in[2]
rlabel metal1 35144 2414 35144 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal2 20194 1622 20194 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 22310 1622 22310 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 24426 1622 24426 1622 0 gfpga_pad_io_soc_out[2]
rlabel metal2 26542 1622 26542 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 37122 1520 37122 1520 0 isol_n
rlabel metal1 9706 2550 9706 2550 0 net1
rlabel metal2 2162 8772 2162 8772 0 net10
rlabel metal1 39422 3638 39422 3638 0 net100
rlabel metal1 42136 4658 42136 4658 0 net101
rlabel metal2 38962 6528 38962 6528 0 net102
rlabel via3 46115 23460 46115 23460 0 net103
rlabel metal1 45218 24378 45218 24378 0 net104
rlabel metal2 46782 23528 46782 23528 0 net105
rlabel metal2 47058 23511 47058 23511 0 net106
rlabel metal1 47288 22134 47288 22134 0 net107
rlabel metal1 46092 24038 46092 24038 0 net108
rlabel metal1 34546 21930 34546 21930 0 net109
rlabel metal1 2530 8840 2530 8840 0 net11
rlabel via2 42458 23477 42458 23477 0 net110
rlabel metal2 38318 2652 38318 2652 0 net111
rlabel metal1 8050 18938 8050 18938 0 net112
rlabel metal1 2990 13396 2990 13396 0 net113
rlabel metal1 9844 17306 9844 17306 0 net114
rlabel metal2 9246 17816 9246 17816 0 net115
rlabel metal1 3174 19822 3174 19822 0 net116
rlabel via2 15594 19261 15594 19261 0 net117
rlabel metal1 11546 19278 11546 19278 0 net118
rlabel metal1 6670 18326 6670 18326 0 net119
rlabel metal1 38318 10064 38318 10064 0 net12
rlabel metal1 8096 20026 8096 20026 0 net120
rlabel metal1 12512 20434 12512 20434 0 net121
rlabel metal1 3450 22610 3450 22610 0 net122
rlabel metal1 6670 21930 6670 21930 0 net123
rlabel metal1 2990 13940 2990 13940 0 net124
rlabel metal1 11592 20434 11592 20434 0 net125
rlabel metal1 5382 20978 5382 20978 0 net126
rlabel metal1 11914 20808 11914 20808 0 net127
rlabel metal1 7544 20910 7544 20910 0 net128
rlabel metal1 6072 20570 6072 20570 0 net129
rlabel via2 1794 9435 1794 9435 0 net13
rlabel metal2 5382 18785 5382 18785 0 net130
rlabel metal1 7314 19822 7314 19822 0 net131
rlabel metal1 6486 20434 6486 20434 0 net132
rlabel metal1 7222 21386 7222 21386 0 net133
rlabel metal1 8004 22474 8004 22474 0 net134
rlabel metal1 6256 14382 6256 14382 0 net135
rlabel metal1 3864 14994 3864 14994 0 net136
rlabel metal2 10258 14994 10258 14994 0 net137
rlabel metal2 10902 15606 10902 15606 0 net138
rlabel metal1 13018 17136 13018 17136 0 net139
rlabel metal2 36478 4794 36478 4794 0 net14
rlabel metal1 3680 17170 3680 17170 0 net140
rlabel metal2 10442 17204 10442 17204 0 net141
rlabel metal1 10810 15878 10810 15878 0 net142
rlabel metal1 41906 3536 41906 3536 0 net143
rlabel metal2 38686 7616 38686 7616 0 net144
rlabel metal1 47886 5202 47886 5202 0 net145
rlabel metal1 40158 7786 40158 7786 0 net146
rlabel metal1 47840 5678 47840 5678 0 net147
rlabel metal1 47794 6290 47794 6290 0 net148
rlabel metal1 47932 6766 47932 6766 0 net149
rlabel metal2 2162 10948 2162 10948 0 net15
rlabel metal2 45862 9248 45862 9248 0 net150
rlabel metal2 38410 9792 38410 9792 0 net151
rlabel metal2 47150 9180 47150 9180 0 net152
rlabel metal2 46782 9214 46782 9214 0 net153
rlabel metal1 41998 3026 41998 3026 0 net154
rlabel metal1 42941 11050 42941 11050 0 net155
rlabel metal1 42826 11560 42826 11560 0 net156
rlabel metal2 47242 10948 47242 10948 0 net157
rlabel metal2 46598 10812 46598 10812 0 net158
rlabel metal1 47472 10642 47472 10642 0 net159
rlabel metal1 39560 11254 39560 11254 0 net16
rlabel metal1 47380 11118 47380 11118 0 net160
rlabel metal1 47058 11730 47058 11730 0 net161
rlabel metal1 47058 12614 47058 12614 0 net162
rlabel metal1 47932 12818 47932 12818 0 net163
rlabel metal1 47288 13294 47288 13294 0 net164
rlabel metal2 37398 4352 37398 4352 0 net165
rlabel metal2 45770 4318 45770 4318 0 net166
rlabel metal2 41354 4386 41354 4386 0 net167
rlabel metal2 37858 4896 37858 4896 0 net168
rlabel metal2 37674 5984 37674 5984 0 net169
rlabel metal1 38686 11798 38686 11798 0 net17
rlabel metal2 47058 4828 47058 4828 0 net170
rlabel metal1 42090 7208 42090 7208 0 net171
rlabel metal2 37950 7038 37950 7038 0 net172
rlabel metal1 7314 22950 7314 22950 0 net173
rlabel metal1 7452 24174 7452 24174 0 net174
rlabel metal1 9338 23732 9338 23732 0 net175
rlabel metal2 11178 23324 11178 23324 0 net176
rlabel metal1 12558 23664 12558 23664 0 net177
rlabel metal1 12144 22202 12144 22202 0 net178
rlabel metal1 12880 21590 12880 21590 0 net179
rlabel via2 40434 11747 40434 11747 0 net18
rlabel metal1 14352 22610 14352 22610 0 net180
rlabel metal1 13846 21658 13846 21658 0 net181
rlabel metal1 14398 22066 14398 22066 0 net182
rlabel metal1 13110 23630 13110 23630 0 net183
rlabel metal1 4370 22950 4370 22950 0 net184
rlabel metal1 17618 21590 17618 21590 0 net185
rlabel metal1 19458 19958 19458 19958 0 net186
rlabel metal2 19642 23528 19642 23528 0 net187
rlabel metal1 19067 21998 19067 21998 0 net188
rlabel metal1 20976 21590 20976 21590 0 net189
rlabel metal1 4232 18190 4232 18190 0 net19
rlabel metal1 18676 23698 18676 23698 0 net190
rlabel metal2 19458 23018 19458 23018 0 net191
rlabel metal2 18906 24446 18906 24446 0 net192
rlabel metal2 21482 23834 21482 23834 0 net193
rlabel metal1 21390 24140 21390 24140 0 net194
rlabel metal1 4600 19278 4600 19278 0 net195
rlabel metal1 4278 18258 4278 18258 0 net196
rlabel metal2 6026 23052 6026 23052 0 net197
rlabel metal2 4738 23494 4738 23494 0 net198
rlabel metal1 4508 23018 4508 23018 0 net199
rlabel metal1 46506 21658 46506 21658 0 net2
rlabel metal1 5658 19346 5658 19346 0 net20
rlabel metal2 4646 24004 4646 24004 0 net200
rlabel metal2 7498 23324 7498 23324 0 net201
rlabel metal1 6946 23086 6946 23086 0 net202
rlabel metal1 13662 2414 13662 2414 0 net203
rlabel metal1 16560 2414 16560 2414 0 net204
rlabel metal1 18492 2414 18492 2414 0 net205
rlabel metal1 19550 3094 19550 3094 0 net206
rlabel metal1 19872 2414 19872 2414 0 net207
rlabel metal1 22264 2414 22264 2414 0 net208
rlabel metal1 23046 3162 23046 3162 0 net209
rlabel metal1 16192 15334 16192 15334 0 net21
rlabel metal1 26910 2822 26910 2822 0 net210
rlabel metal1 16836 17646 16836 17646 0 net211
rlabel metal2 23690 13311 23690 13311 0 net212
rlabel metal2 27922 21250 27922 21250 0 net213
rlabel metal1 18906 14042 18906 14042 0 net214
rlabel metal2 24610 20910 24610 20910 0 net215
rlabel metal1 19504 13226 19504 13226 0 net216
rlabel metal1 31096 14382 31096 14382 0 net217
rlabel metal2 31142 8058 31142 8058 0 net218
rlabel metal1 30314 10098 30314 10098 0 net219
rlabel metal1 7866 16490 7866 16490 0 net22
rlabel metal2 33902 15232 33902 15232 0 net220
rlabel metal1 28934 13294 28934 13294 0 net221
rlabel metal2 29946 9282 29946 9282 0 net222
rlabel metal2 31418 7616 31418 7616 0 net223
rlabel metal1 32844 14042 32844 14042 0 net224
rlabel metal1 29164 8874 29164 8874 0 net225
rlabel metal1 27002 11866 27002 11866 0 net226
rlabel metal1 32752 7854 32752 7854 0 net227
rlabel metal1 29302 19346 29302 19346 0 net228
rlabel metal1 31372 15130 31372 15130 0 net229
rlabel metal2 9522 14858 9522 14858 0 net23
rlabel metal1 36478 17306 36478 17306 0 net230
rlabel metal1 35374 15130 35374 15130 0 net231
rlabel metal1 35834 13226 35834 13226 0 net232
rlabel metal1 31280 10778 31280 10778 0 net233
rlabel metal1 33120 21658 33120 21658 0 net234
rlabel metal1 25208 13294 25208 13294 0 net235
rlabel metal1 24104 13838 24104 13838 0 net236
rlabel metal2 20010 11611 20010 11611 0 net237
rlabel metal1 25024 10642 25024 10642 0 net238
rlabel metal2 22678 10880 22678 10880 0 net239
rlabel metal1 20332 19822 20332 19822 0 net24
rlabel metal1 18492 12750 18492 12750 0 net240
rlabel metal1 18446 8398 18446 8398 0 net241
rlabel metal1 19688 10098 19688 10098 0 net242
rlabel metal1 22310 7854 22310 7854 0 net243
rlabel metal1 30912 18258 30912 18258 0 net244
rlabel metal1 12972 13362 12972 13362 0 net245
rlabel metal1 13064 18394 13064 18394 0 net246
rlabel metal1 12880 18666 12880 18666 0 net247
rlabel metal1 10350 18394 10350 18394 0 net248
rlabel metal1 13984 20570 13984 20570 0 net249
rlabel metal1 4370 2414 4370 2414 0 net25
rlabel metal1 12650 21080 12650 21080 0 net250
rlabel metal1 15824 20570 15824 20570 0 net251
rlabel metal1 35742 18598 35742 18598 0 net252
rlabel metal1 39330 20570 39330 20570 0 net253
rlabel metal2 18722 9792 18722 9792 0 net254
rlabel metal1 17296 10710 17296 10710 0 net255
rlabel metal1 11638 13906 11638 13906 0 net256
rlabel metal1 16376 14314 16376 14314 0 net257
rlabel metal1 21528 12206 21528 12206 0 net258
rlabel metal1 21574 11730 21574 11730 0 net259
rlabel metal2 1794 3570 1794 3570 0 net26
rlabel metal1 18492 18598 18492 18598 0 net260
rlabel metal1 18584 19822 18584 19822 0 net261
rlabel metal1 23276 17578 23276 17578 0 net262
rlabel metal1 45218 24242 45218 24242 0 net263
rlabel metal2 42734 23171 42734 23171 0 net264
rlabel metal1 42366 24174 42366 24174 0 net265
rlabel metal1 48714 24208 48714 24208 0 net266
rlabel metal2 44022 23494 44022 23494 0 net267
rlabel metal1 48852 23290 48852 23290 0 net268
rlabel metal1 43424 23018 43424 23018 0 net269
rlabel metal1 2438 3570 2438 3570 0 net27
rlabel metal1 10534 3366 10534 3366 0 net270
rlabel metal1 13938 2958 13938 2958 0 net271
rlabel metal1 48254 23120 48254 23120 0 net272
rlabel metal1 47794 23562 47794 23562 0 net273
rlabel metal2 10350 3332 10350 3332 0 net274
rlabel metal1 9752 2414 9752 2414 0 net275
rlabel metal1 38732 5270 38732 5270 0 net28
rlabel metal1 37766 5304 37766 5304 0 net29
rlabel metal1 5083 2550 5083 2550 0 net3
rlabel metal1 37812 6290 37812 6290 0 net30
rlabel metal1 15870 17238 15870 17238 0 net31
rlabel metal1 2576 5882 2576 5882 0 net32
rlabel metal2 48438 14552 48438 14552 0 net33
rlabel metal2 35466 16167 35466 16167 0 net34
rlabel metal4 14260 14892 14260 14892 0 net35
rlabel metal2 48438 18462 48438 18462 0 net36
rlabel metal1 15318 19822 15318 19822 0 net37
rlabel via2 16238 19363 16238 19363 0 net38
rlabel metal1 19458 15674 19458 15674 0 net39
rlabel metal1 1794 5576 1794 5576 0 net4
rlabel metal2 48438 19822 48438 19822 0 net40
rlabel metal1 18446 15674 18446 15674 0 net41
rlabel metal1 12742 20502 12742 20502 0 net42
rlabel metal1 15088 19142 15088 19142 0 net43
rlabel metal2 14490 13532 14490 13532 0 net44
rlabel metal1 48438 21012 48438 21012 0 net45
rlabel metal1 48852 22406 48852 22406 0 net46
rlabel metal2 18998 16235 18998 16235 0 net47
rlabel metal1 47288 22950 47288 22950 0 net48
rlabel metal1 45816 21862 45816 21862 0 net49
rlabel metal1 37812 7786 37812 7786 0 net5
rlabel metal1 40572 22610 40572 22610 0 net50
rlabel metal1 13248 17306 13248 17306 0 net51
rlabel metal1 41170 24072 41170 24072 0 net52
rlabel metal1 46966 22202 46966 22202 0 net53
rlabel metal2 49174 24089 49174 24089 0 net54
rlabel metal3 17457 13668 17457 13668 0 net55
rlabel metal1 16744 14246 16744 14246 0 net56
rlabel metal1 48944 15674 48944 15674 0 net57
rlabel metal1 21298 13226 21298 13226 0 net58
rlabel metal1 21344 9622 21344 9622 0 net59
rlabel metal1 2530 6664 2530 6664 0 net6
rlabel metal2 13938 18445 13938 18445 0 net60
rlabel metal2 48438 17442 48438 17442 0 net61
rlabel metal3 16928 13804 16928 13804 0 net62
rlabel metal1 26404 19414 26404 19414 0 net63
rlabel metal2 27554 18530 27554 18530 0 net64
rlabel metal2 31786 18173 31786 18173 0 net65
rlabel metal2 32062 23800 32062 23800 0 net66
rlabel metal2 30038 23341 30038 23341 0 net67
rlabel metal1 38732 24038 38732 24038 0 net68
rlabel metal1 33166 19822 33166 19822 0 net69
rlabel metal2 1794 6460 1794 6460 0 net7
rlabel metal1 35236 19822 35236 19822 0 net70
rlabel metal2 43746 23885 43746 23885 0 net71
rlabel metal1 34132 21658 34132 21658 0 net72
rlabel metal2 44390 24412 44390 24412 0 net73
rlabel metal2 21114 21981 21114 21981 0 net74
rlabel metal2 36662 19788 36662 19788 0 net75
rlabel metal2 41170 20111 41170 20111 0 net76
rlabel metal1 43332 22542 43332 22542 0 net77
rlabel metal3 36524 18632 36524 18632 0 net78
rlabel metal1 33166 20774 33166 20774 0 net79
rlabel metal1 40572 8466 40572 8466 0 net8
rlabel via2 31786 20859 31786 20859 0 net80
rlabel metal1 34316 19890 34316 19890 0 net81
rlabel via2 41906 22389 41906 22389 0 net82
rlabel via2 45586 22491 45586 22491 0 net83
rlabel metal1 44206 22474 44206 22474 0 net84
rlabel metal2 16238 24242 16238 24242 0 net85
rlabel metal2 27278 19516 27278 19516 0 net86
rlabel metal1 32982 15606 32982 15606 0 net87
rlabel metal1 32706 21522 32706 21522 0 net88
rlabel metal1 35972 16626 35972 16626 0 net89
rlabel metal1 1794 7752 1794 7752 0 net9
rlabel metal1 32614 18156 32614 18156 0 net90
rlabel metal1 28060 21930 28060 21930 0 net91
rlabel metal1 26910 19754 26910 19754 0 net92
rlabel metal1 27738 3502 27738 3502 0 net93
rlabel metal1 29256 2550 29256 2550 0 net94
rlabel metal1 32890 2550 32890 2550 0 net95
rlabel metal1 33994 2618 33994 2618 0 net96
rlabel metal2 37766 2822 37766 2822 0 net97
rlabel metal2 46506 23698 46506 23698 0 net98
rlabel metal1 43838 2516 43838 2516 0 net99
rlabel metal2 39238 2132 39238 2132 0 prog_clk
rlabel metal1 43056 24174 43056 24174 0 prog_reset
rlabel metal1 43378 2278 43378 2278 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 45586 2098 45586 2098 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 47702 2336 47702 2336 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 46690 4488 46690 4488 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 30682 12750 30682 12750 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal1 23644 18666 23644 18666 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal1 31418 21386 31418 21386 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 24380 17102 24380 17102 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal2 21390 14994 21390 14994 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal1 18630 18258 18630 18258 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel metal1 21436 13362 21436 13362 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 21068 17238 21068 17238 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 18446 21114 18446 21114 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal2 21390 17578 21390 17578 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 19826 20570 19826 20570 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal1 18262 21454 18262 21454 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 21436 18802 21436 18802 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal1 18998 19890 18998 19890 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal1 21735 19278 21735 19278 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal1 24426 20366 24426 20366 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 24932 19278 24932 19278 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal1 18860 20570 18860 20570 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal1 25254 18836 25254 18836 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 17112 20366 17112 20366 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal1 26864 20366 26864 20366 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal1 32706 19924 32706 19924 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal1 26404 16626 26404 16626 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal2 24886 23324 24886 23324 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal1 32890 22508 32890 22508 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 28520 22066 28520 22066 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal1 17986 16082 17986 16082 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel metal2 21482 20638 21482 20638 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 18630 15164 18630 15164 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal1 27462 22984 27462 22984 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel metal1 22954 22066 22954 22066 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal1 25254 15572 25254 15572 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 21988 13838 21988 13838 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal1 18032 21930 18032 21930 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal2 32614 16354 32614 16354 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel metal2 33902 13056 33902 13056 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 30774 16252 30774 16252 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal1 37950 11050 37950 11050 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal2 36662 10948 36662 10948 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal2 36110 10268 36110 10268 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 36202 10608 36202 10608 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal1 37214 12342 37214 12342 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal1 33120 10778 33120 10778 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 32430 11424 32430 11424 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal1 36984 16014 36984 16014 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal1 32476 16490 32476 16490 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 35558 15538 35558 15538 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal1 33626 11696 33626 11696 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal2 29946 17408 29946 17408 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal1 29808 15130 29808 15130 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal2 31878 9146 31878 9146 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal1 30774 14960 30774 14960 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 30130 10574 30130 10574 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal2 34086 8738 34086 8738 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal1 32384 14450 32384 14450 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal1 32430 8398 32430 8398 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal2 38226 13634 38226 13634 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel metal1 33948 11050 33948 11050 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 36524 14586 36524 14586 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal1 32660 10098 32660 10098 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal1 29670 16626 29670 16626 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 27830 17034 27830 17034 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 34132 7922 34132 7922 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 36708 12070 36708 12070 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal2 30314 23324 30314 23324 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel metal1 41538 22984 41538 22984 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 32338 21862 32338 21862 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal2 37674 20570 37674 20570 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal1 35788 18666 35788 18666 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal2 37766 19720 37766 19720 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 34224 18190 34224 18190 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal2 38042 18224 38042 18224 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel metal2 39422 19108 39422 19108 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 37950 17102 37950 17102 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 38548 16150 38548 16150 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal1 40112 18598 40112 18598 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 38548 16626 38548 16626 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal2 37766 16932 37766 16932 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 40158 15878 40158 15878 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 39238 14416 39238 14416 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal2 32338 14450 32338 14450 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal1 38456 14314 38456 14314 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 38272 14246 38272 14246 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal1 34086 23630 34086 23630 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal1 32430 19788 32430 19788 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 35190 23630 35190 23630 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 25576 14586 25576 14586 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel via1 27094 13838 27094 13838 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 23736 12750 23736 12750 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal1 25116 14042 25116 14042 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal2 24886 11730 24886 11730 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 26864 12342 26864 12342 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 22908 13362 22908 13362 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 27324 15538 27324 15538 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 21390 10506 21390 10506 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 23644 9350 23644 9350 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 19826 8602 19826 8602 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal1 21620 8602 21620 8602 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 19596 9622 19596 9622 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal2 19458 9078 19458 9078 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 20056 12750 20056 12750 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal2 21114 10132 21114 10132 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20884 12750 20884 12750 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal1 25622 15130 25622 15130 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal2 32338 20672 32338 20672 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal1 36432 20842 36432 20842 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 33764 20502 33764 20502 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal2 13294 14212 13294 14212 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal1 14214 10574 14214 10574 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal2 14582 18428 14582 18428 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 17342 15572 17342 15572 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 13110 18836 13110 18836 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal1 16008 18938 16008 18938 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 11362 18190 11362 18190 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal1 12466 14892 12466 14892 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14306 21352 14306 21352 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal1 15962 20842 15962 20842 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 15364 22202 15364 22202 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal1 16468 21318 16468 21318 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 18676 23018 18676 23018 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel metal1 36846 23154 36846 23154 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal1 40848 22066 40848 22066 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal2 37490 23018 37490 23018 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal2 37398 21505 37398 21505 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 36248 22066 36248 22066 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 14720 18258 14720 18258 0 sb_1__0_.mux_left_track_1.out
rlabel metal1 26910 18258 26910 18258 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26772 18394 26772 18394 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23414 14348 23414 14348 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22402 12376 22402 12376 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 25070 17884 25070 17884 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24380 15946 24380 15946 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 22034 18190 22034 18190 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 8326 18088 8326 18088 0 sb_1__0_.mux_left_track_11.out
rlabel metal1 22908 18258 22908 18258 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23276 18326 23276 18326 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 14246 20930 14246 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20378 15062 20378 15062 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20930 18088 20930 18088 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19504 15130 19504 15130 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16606 18394 16606 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 15548 16218 15548 16218 0 sb_1__0_.mux_left_track_13.out
rlabel metal1 27186 21624 27186 21624 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21850 21896 21850 21896 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 15674 21022 15674 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21482 21896 21482 21896 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 18938 18262 18938 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13662 19788 13662 19788 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9706 21318 9706 21318 0 sb_1__0_.mux_left_track_21.out
rlabel metal1 26496 23290 26496 23290 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24610 22168 24610 22168 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21068 18938 21068 18938 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19780 24582 19780 24582 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 20026 18262 20026 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel via2 9890 20451 9890 20451 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 13570 16813 13570 16813 0 sb_1__0_.mux_left_track_29.out
rlabel metal2 29578 21182 29578 21182 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 26818 20434 26818 20434 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23966 15130 23966 15130 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23966 20264 23966 20264 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22954 17850 22954 17850 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14122 17646 14122 17646 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9982 20740 9982 20740 0 sb_1__0_.mux_left_track_3.out
rlabel metal2 20378 18394 20378 18394 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22494 18632 22494 18632 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19918 19210 19918 19210 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17388 17850 17388 17850 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13570 19924 13570 19924 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9338 16048 9338 16048 0 sb_1__0_.mux_left_track_37.out
rlabel metal2 32154 19006 32154 19006 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29256 18394 29256 18394 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 16660 23782 16660 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23874 13498 23874 13498 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21850 15504 21850 15504 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8326 18768 8326 18768 0 sb_1__0_.mux_left_track_45.out
rlabel metal1 29670 21930 29670 21930 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28336 22134 28336 22134 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28106 21658 28106 21658 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 11362 21981 11362 21981 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9154 19482 9154 19482 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 24058 20026 24058 20026 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24242 18122 24242 18122 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17894 15980 17894 15980 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18354 15130 18354 15130 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16928 16218 16928 16218 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13570 20978 13570 20978 0 sb_1__0_.mux_left_track_53.out
rlabel metal1 26956 21998 26956 21998 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22080 20774 22080 20774 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20792 20910 20792 20910 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13754 20944 13754 20944 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14766 16048 14766 16048 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 25392 15470 25392 15470 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 15402 24104 15402 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20148 13158 20148 13158 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21942 15504 21942 15504 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20378 13498 20378 13498 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19918 16388 19918 16388 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39514 14110 39514 14110 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 31142 17306 31142 17306 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33350 13396 33350 13396 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29900 14314 29900 14314 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32798 16218 32798 16218 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33350 15300 33350 15300 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 39330 14909 39330 14909 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43263 11254 43263 11254 0 sb_1__0_.mux_right_track_10.out
rlabel metal1 34776 13906 34776 13906 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34684 14042 34684 14042 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 36386 9860 36386 9860 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 36478 9520 36478 9520 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel via1 35834 11883 35834 11883 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 36846 11254 36846 11254 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 40526 11118 40526 11118 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 43056 11798 43056 11798 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 33258 14382 33258 14382 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 33718 15130 33718 15130 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32614 10540 32614 10540 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 37398 12347 37398 12347 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36754 10472 36754 10472 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39330 12206 39330 12206 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45678 14348 45678 14348 0 sb_1__0_.mux_right_track_2.out
rlabel metal1 35098 19414 35098 19414 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34132 18394 34132 18394 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33810 14756 33810 14756 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37490 17510 37490 17510 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 34270 14688 34270 14688 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 40894 16388 40894 16388 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44390 10642 44390 10642 0 sb_1__0_.mux_right_track_20.out
rlabel metal2 30866 18156 30866 18156 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30820 16218 30820 16218 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28336 11866 28336 11866 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33764 11730 33764 11730 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33856 11730 33856 11730 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38226 11220 38226 11220 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 41998 8534 41998 8534 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 30268 13362 30268 13362 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30176 13294 30176 13294 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27232 9418 27232 9418 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32476 9690 32476 9690 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32384 9554 32384 9554 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37674 8976 37674 8976 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44942 7888 44942 7888 0 sb_1__0_.mux_right_track_36.out
rlabel metal1 32292 11866 32292 11866 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32752 11866 32752 11866 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34914 8806 34914 8806 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32982 8058 32982 8058 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38962 8500 38962 8500 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 45954 12988 45954 12988 0 sb_1__0_.mux_right_track_4.out
rlabel metal1 35972 17170 35972 17170 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36340 16762 36340 16762 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33994 11696 33994 11696 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37260 13974 37260 13974 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37168 14042 37168 14042 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 41354 13668 41354 13668 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 42734 6358 42734 6358 0 sb_1__0_.mux_right_track_44.out
rlabel metal1 32568 10166 32568 10166 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 31970 9384 31970 9384 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36570 9928 36570 9928 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 41860 5678 41860 5678 0 sb_1__0_.mux_right_track_52.out
rlabel metal1 32384 12818 32384 12818 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29762 12954 29762 12954 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35558 8942 35558 8942 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43585 12070 43585 12070 0 sb_1__0_.mux_right_track_6.out
rlabel metal1 36018 15062 36018 15062 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36202 15130 36202 15130 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38364 12614 38364 12614 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 39054 9860 39054 9860 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38686 12274 38686 12274 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 38686 11968 38686 11968 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 41446 12240 41446 12240 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 23828 23290 23828 23290 0 sb_1__0_.mux_top_track_0.out
rlabel metal1 35834 21862 35834 21862 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38502 23562 38502 23562 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24932 19958 24932 19958 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 19482 28612 19482 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32246 23528 32246 23528 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29624 20774 29624 20774 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 29762 23426 29762 23426 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 21390 21471 21390 21471 0 sb_1__0_.mux_top_track_10.out
rlabel metal1 36018 19482 36018 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40112 19482 40112 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36018 19686 36018 19686 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 31694 17510 31694 17510 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 31096 18938 31096 18938 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal3 27462 22372 27462 22372 0 sb_1__0_.mux_top_track_12.out
rlabel metal2 40894 19040 40894 19040 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39100 18394 39100 18394 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36984 17034 36984 17034 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36064 20298 36064 20298 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 22831 19826 22831 0 sb_1__0_.mux_top_track_14.out
rlabel metal1 40848 17714 40848 17714 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40250 17850 40250 17850 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35926 14790 35926 14790 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 38042 19057 38042 19057 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20746 19295 20746 19295 0 sb_1__0_.mux_top_track_16.out
rlabel metal2 40986 16320 40986 16320 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38870 16218 38870 16218 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35604 13498 35604 13498 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35742 18394 35742 18394 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24702 17850 24702 17850 0 sb_1__0_.mux_top_track_18.out
rlabel metal1 39422 15130 39422 15130 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39238 14858 39238 14858 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32246 14994 32246 14994 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32039 14858 32039 14858 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21390 23722 21390 23722 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 36800 23766 36800 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38962 23834 38962 23834 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32798 20978 32798 20978 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35144 23834 35144 23834 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32890 21862 32890 21862 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 28658 23766 28658 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel via2 8418 20893 8418 20893 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 26358 17306 26358 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 25622 15334 25622 15334 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24932 17306 24932 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20102 16456 20102 16456 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 24656 15062 24656 15062 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 13158 23322 13158 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21206 16456 21206 16456 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15962 18122 15962 18122 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 26956 15878 26956 15878 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23276 12138 23276 12138 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 18538 15470 18538 15470 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19412 17850 19412 17850 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 23184 13158 23184 13158 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22678 13226 22678 13226 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20470 17578 20470 17578 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14490 17306 14490 17306 0 sb_1__0_.mux_top_track_28.out
rlabel metal2 22310 10200 22310 10200 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15594 12682 15594 12682 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13248 17850 13248 17850 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 21344 7514 21344 7514 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15732 17850 15732 17850 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12650 16422 12650 16422 0 sb_1__0_.mux_top_track_32.out
rlabel metal1 18262 10234 18262 10234 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14766 11254 14766 11254 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13662 24140 13662 24140 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 19642 10778 19642 10778 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18538 12682 18538 12682 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14490 22100 14490 22100 0 sb_1__0_.mux_top_track_36.out
rlabel metal2 22678 13872 22678 13872 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 12818 21528 12818 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20746 12903 20746 12903 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27370 23290 27370 23290 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 35742 20570 35742 20570 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37214 21590 37214 21590 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35742 21216 35742 21216 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31050 18394 31050 18394 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30866 20808 30866 20808 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9798 18360 9798 18360 0 sb_1__0_.mux_top_track_40.out
rlabel metal1 13018 10778 13018 10778 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11546 14586 11546 14586 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9522 22882 9522 22882 0 sb_1__0_.mux_top_track_42.out
rlabel metal1 16698 15674 16698 15674 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13938 18156 13938 18156 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2162 23732 2162 23732 0 sb_1__0_.mux_top_track_44.out
rlabel metal2 15594 17952 15594 17952 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12558 19941 12558 19941 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3450 18292 3450 18292 0 sb_1__0_.mux_top_track_46.out
rlabel metal1 11868 15130 11868 15130 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10120 18054 10120 18054 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7084 23222 7084 23222 0 sb_1__0_.mux_top_track_48.out
rlabel metal1 16422 19482 16422 19482 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11086 20740 11086 20740 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7636 23630 7636 23630 0 sb_1__0_.mux_top_track_50.out
rlabel metal1 16882 18938 16882 18938 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8602 21930 8602 21930 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9246 23086 9246 23086 0 sb_1__0_.mux_top_track_58.out
rlabel metal1 18906 24786 18906 24786 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15594 22440 15594 22440 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19642 24242 19642 24242 0 sb_1__0_.mux_top_track_6.out
rlabel metal1 40388 22202 40388 22202 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 41446 22491 41446 22491 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 36202 21964 36202 21964 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40112 22950 40112 22950 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35834 22746 35834 22746 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 29946 24021 29946 24021 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 31510 22457 31510 22457 0 sb_1__0_.mux_top_track_8.out
rlabel metal1 40112 20978 40112 20978 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40848 20842 40848 20842 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 34270 19482 34270 19482 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40204 21114 40204 21114 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36662 24106 36662 24106 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 36110 23817 36110 23817 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45402 25493 45402 25493 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 47886 24106 47886 24106 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46828 23086 46828 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal2 47242 24463 47242 24463 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal2 47932 24140 47932 24140 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48162 23834 48162 23834 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44252 22678 44252 22678 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 45080 23018 45080 23018 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 1150 2115 1150 2115 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 3266 1299 3266 1299 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 19136 13906 19136 13906 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 19872 12614 19872 12614 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
