* NGSPICE file created from right_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

.subckt right_tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ ccff_head_0_0 ccff_head_1 ccff_head_2 ccff_tail ccff_tail_0 ccff_tail_1 chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23]
+ chanx_left_in[24] chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28]
+ chanx_left_in[29] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23]
+ chanx_left_out[24] chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28]
+ chanx_left_out[29] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21]
+ chany_bottom_in[22] chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25]
+ chany_bottom_in[26] chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29]
+ chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6]
+ chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10]
+ chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14]
+ chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18]
+ chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21]
+ chany_bottom_out[22] chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25]
+ chany_bottom_out[26] chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in_0[0] chany_top_in_0[10] chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13]
+ chany_top_in_0[14] chany_top_in_0[15] chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18]
+ chany_top_in_0[19] chany_top_in_0[1] chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22]
+ chany_top_in_0[23] chany_top_in_0[24] chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27]
+ chany_top_in_0[28] chany_top_in_0[29] chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4]
+ chany_top_in_0[5] chany_top_in_0[6] chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9]
+ chany_top_out_0[0] chany_top_out_0[10] chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13]
+ chany_top_out_0[14] chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17]
+ chany_top_out_0[18] chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21]
+ chany_top_out_0[22] chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25]
+ chany_top_out_0[26] chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29]
+ chany_top_out_0[2] chany_top_out_0[3] chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6]
+ chany_top_out_0[7] chany_top_out_0[8] chany_top_out_0[9] clk0 gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n left_width_0_height_0_subtile_0__pin_inpad_0_
+ left_width_0_height_0_subtile_1__pin_inpad_0_ left_width_0_height_0_subtile_2__pin_inpad_0_
+ left_width_0_height_0_subtile_3__pin_inpad_0_ prog_clk prog_reset_bottom_in prog_reset_bottom_out
+ prog_reset_left_in prog_reset_top_in prog_reset_top_out reset_bottom_in reset_bottom_out
+ reset_left_out reset_right_in reset_top_in reset_top_out right_width_0_height_0_subtile_0__pin_O_10_
+ right_width_0_height_0_subtile_0__pin_O_11_ right_width_0_height_0_subtile_0__pin_O_12_
+ right_width_0_height_0_subtile_0__pin_O_13_ right_width_0_height_0_subtile_0__pin_O_14_
+ right_width_0_height_0_subtile_0__pin_O_15_ right_width_0_height_0_subtile_0__pin_O_8_
+ right_width_0_height_0_subtile_0__pin_O_9_ sc_in sc_out test_enable_bottom_in test_enable_bottom_out
+ test_enable_left_out test_enable_right_in test_enable_top_in test_enable_top_out
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ top_width_0_height_0_subtile_0__pin_O_0_ top_width_0_height_0_subtile_0__pin_O_1_
+ top_width_0_height_0_subtile_0__pin_O_2_ top_width_0_height_0_subtile_0__pin_O_3_
+ top_width_0_height_0_subtile_0__pin_O_4_ top_width_0_height_0_subtile_0__pin_O_5_
+ top_width_0_height_0_subtile_0__pin_O_6_ top_width_0_height_0_subtile_0__pin_O_7_
+ top_width_0_height_0_subtile_0__pin_cin_0_ top_width_0_height_0_subtile_0__pin_reg_in_0_
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_36.mux_l2_in_1__374 VGND VGND VPWR VPWR net374 sb_8__1_.mux_top_track_36.mux_l2_in_1__374/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_2__A0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_53_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_2__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net307 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_2.mux_l2_in_3_ net371 net32 sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_2.mem_out\[2\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_363_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input92_A chany_top_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_294_ sb_8__1_.mux_left_track_3.out VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_29.mux_l2_in_1__334 VGND VGND VPWR VPWR net334 sb_8__1_.mux_bottom_track_29.mux_l2_in_1__334/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__304__A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_2_ net7 net19 sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_17.mux_l1_in_0__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net311 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk sb_8__1_.mem_left_track_21.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_23.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_346_ net47 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_277_ sb_8__1_.mux_left_track_37.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_36.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput242 net242 VGND VGND VPWR VPWR test_enable_top_out sky130_fd_sc_hd__buf_12
Xoutput231 net231 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
Xoutput220 net220 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_87_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_44_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_3__330 VGND VGND VPWR VPWR net330 sb_8__1_.mux_bottom_track_1.mux_l2_in_3__330/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input55_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ sb_8__1_.mux_top_track_52.out VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_2.mux_l4_in_0_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X
+ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sb_8__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_3__259 VGND VGND VPWR VPWR net259 cbx_8__1_.mux_top_ipin_7.mux_l2_in_3__259/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mux_top_ipin_5.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_2_ sb_8__1_.mux_left_track_21.out net14 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_0__A0 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk sb_8__1_.mem_left_track_29.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_15.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_45_prog_clk sb_8__1_.mem_bottom_track_7.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__312__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_45.mux_l1_in_0_ net243 net92 sb_8__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__291
+ VGND VGND VPWR VPWR net291 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__291/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_57.mux_l2_in_0_ net365 sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X
+ cbx_8__1_.ccff_head VGND VGND VPWR VPWR sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input18_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_0__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_2.mux_l3_in_1_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_28.mux_l1_in_3__373 VGND VGND VPWR VPWR net373 sb_8__1_.mux_top_track_28.mux_l1_in_3__373/LO
+ sky130_fd_sc_hd__conb_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_0__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2__A0 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l2_in_1__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l2_in_0_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_1_ net9 cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput120 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND VPWR
+ VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_13.mux_l2_in_1__343 VGND VGND VPWR VPWR net343 sb_8__1_.mux_left_track_13.mux_l2_in_1__343/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_sb_8__1_.mux_left_track_25.mux_l1_in_0__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_2__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net97 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_2.mux_l2_in_2_ net14 net63 sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_60_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_2.mem_out\[1\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
X_362_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_293_ sb_8__1_.mux_left_track_5.out VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input85_A chany_top_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_52_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_1_ net231 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_33.mux_l1_in_1__354 VGND VGND VPWR VPWR net354 sb_8__1_.mux_left_track_33.mux_l1_in_1__354/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mux_top_ipin_15.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_17.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_1.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_12_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_2__A0 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__321
+ VGND VGND VPWR VPWR net321 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__321/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
X_345_ sb_8__1_.mux_top_track_20.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
X_276_ net248 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_2__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_36.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__315__A sb_8__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_2
Xoutput210 net210 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xoutput243 net243 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
Xoutput232 net232 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
Xoutput221 net221 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_44_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_3__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_328_ net57 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input102_A reset_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk sb_8__1_.mem_left_track_27.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_0__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_45_prog_clk sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_66_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_15.mux_l2_in_1__A1 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_45_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_80_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_33.mux_l1_in_0__A0 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_2.mux_l3_in_0_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net291 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__mux2_8
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__A1 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2__A1 net68 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_14_prog_clk sb_8__1_.mem_left_track_41.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_41.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_15_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_29_prog_clk cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ net99 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfrtp_2
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput110 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput121 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input30_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_42_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3_ net276 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_25.mux_l1_in_0__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__284
+ VGND VGND VPWR VPWR net284 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__284/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_0__A0 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_1.ccff_tail net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__318__A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_15.mux_l3_in_0_ sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_15.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_57.mux_l1_in_0_ net249 net83 sb_8__1_.mem_left_track_57.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_2.mux_l2_in_1_ net49 net119 sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_45_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk sb_8__1_.mem_top_track_2.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net325 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_361_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_292_ sb_8__1_.mux_left_track_7.out VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input78_A chany_top_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output234_A net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_0_ net87 net73 sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_86_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_2__A0 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_20.mux_l1_in_3_ net372 net26 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_8__1_.mem_bottom_track_1.ccff_head
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_2__A1 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4_ net65 net63 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_344_ net44 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_275_ sb_8__1_.mux_left_track_41.out VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_41.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_41.out sky130_fd_sc_hd__clkbuf_2
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_37.mux_l3_in_0_ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__265 VGND VGND VPWR VPWR net265 cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__265/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_15.mux_l2_in_1_ net344 net244 sb_8__1_.mem_left_track_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_91_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2__A0 net74 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_28.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_9_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput200 net200 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput211 net211 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput244 net244 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
Xoutput233 net233 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
XANTENNA__331__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_44_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_23.mux_l2_in_1__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_327_ net56 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__314
+ VGND VGND VPWR VPWR net314 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__314/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__326__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_41.mux_l1_in_0__A0 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.out sky130_fd_sc_hd__clkbuf_1
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net292 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_37.mux_l2_in_1_ net336 net33 sb_8__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3_ net281 net86 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input60_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_1__A0 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_43_prog_clk sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_66_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.mux_l3_in_0_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_44_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_32_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_33.mux_l1_in_0__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__298
+ VGND VGND VPWR VPWR net298 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__298/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_14_prog_clk sb_8__1_.mem_left_track_37.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_41.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_20.mux_l2_in_1_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput111 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net111 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput100 prog_reset_left_in VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
Xinput122 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net122
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__buf_2
XANTENNA_input23_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net320 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__mux2_4
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_3_ net380 sb_8__1_.mux_left_track_51.out cbx_8__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_2_ net57 cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_0__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__334__A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_2.mux_l2_in_0_ net114 sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk sb_8__1_.mem_top_track_0.ccff_tail
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_360_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ sb_8__1_.mux_left_track_9.out VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_31_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_15.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_left_track_19.mux_l2_in_0__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_5.mux_l3_in_0_ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_8__1_.mem_left_track_3.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_15.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_2__A1 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.mux_l1_in_2_ net8 net20 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk cbx_8__1_.mem_top_ipin_1.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3_ sb_8__1_.mux_bottom_track_29.out
+ net40 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_343_ net43 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input90_A chany_top_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_274_ net88 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_47.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_37_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_15.mux_l2_in_0_ net40 sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_15.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2__A1 net43 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput201 net201 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput234 net234 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
Xoutput245 net245 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_1.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_5.mux_l2_in_1_ net361 net248 sb_8__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_326_ net45 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l2_in_2__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__342__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_3_ net258 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.out sky130_fd_sc_hd__buf_4
Xsb_8__1_.mux_bottom_track_37.mux_l2_in_0_ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2_ net45 net66 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input53_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk sb_8__1_.mem_bottom_track_5.ccff_tail
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net127 net98 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_44_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_309_ net69 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mux_top_ipin_1.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_3__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_3__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_2__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_57.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_57.out sky130_fd_sc_hd__clkbuf_2
XFILLER_8_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_4_ sb_8__1_.mux_left_track_37.out net6 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_37.mux_l1_in_1_ net16 net234 sb_8__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_20.mux_l2_in_0_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cbx_8__1_.mem_top_ipin_4.mem_out\[2\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 prog_reset_top_in VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput112 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input16_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_2_ net28 sb_8__1_.mux_left_track_33.out cbx_8__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_8__1_.mux_top_ipin_6.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_35_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_290_ sb_8__1_.mux_left_track_11.out VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__272 VGND VGND VPWR VPWR net272
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__272/LO sky130_fd_sc_hd__conb_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk sb_8__1_.mem_left_track_15.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__282
+ VGND VGND VPWR VPWR net282 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__282/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_76_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_8__1_.mem_left_track_3.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_20.mux_l1_in_1_ net56 net42 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk cbx_8__1_.mem_top_ipin_1.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input118_A top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_342_ net42 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
X_273_ sb_8__1_.mux_left_track_45.out VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input83_A chany_top_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_45.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
Xcbx_8__1_.mux_top_ipin_6.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_37_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_top_track_2.mux_l1_in_0_ net111 net116 sb_8__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3_ net269 net93 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xoutput202 net202 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput213 net213 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput235 net235 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput224 net224 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
Xoutput246 net246 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_5.mux_l2_in_0_ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_51_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_325_ sb_8__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__279 VGND VGND VPWR VPWR net279
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__279/LO sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__A1 net89 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk sb_8__1_.mem_left_track_9.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__303
+ VGND VGND VPWR VPWR net303 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__303/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_2_ net29 cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__269 VGND VGND VPWR VPWR net269
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__269/LO sky130_fd_sc_hd__conb_1
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1_ net35 cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_15.mux_l1_in_0_ net41 net70 sb_8__1_.mem_left_track_15.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_7.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input46_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_43_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_27.mux_l1_in_1__A1 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_1__A0 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ net68 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mux_top_ipin_1.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_27.mux_l2_in_0_ sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_27.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_5.mux_l1_in_1_ net245 net48 sb_8__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_92_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input100_A prog_reset_left_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net106 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_3_ net338 net28 sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_9 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net328 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_3_ sb_8__1_.mux_left_track_25.out net12 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_2__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_37.mux_l1_in_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ net69 sb_8__1_.mem_bottom_track_37.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2_ net72 net41 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail net98 VGND
+ VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XANTENNA__348__A net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__294
+ VGND VGND VPWR VPWR net294 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__294/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput102 reset_bottom_in VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_12
Xinput113 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net113 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_1_ net8 cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_27.mux_l1_in_1_ net350 net250 sb_8__1_.mem_left_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_3__260 VGND VGND VPWR VPWR net260 cbx_8__1_.mux_top_ipin_8.mux_l2_in_3__260/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\] net254 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net302 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__mux2_4
Xsb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_12.mux_l1_in_3__370 VGND VGND VPWR VPWR net370 sb_8__1_.mux_top_track_12.mux_l1_in_3__370/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_2_prog_clk sb_8__1_.mem_left_track_13.ccff_tail
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_40_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_8__1_.mem_left_track_1.ccff_tail
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_20.mux_l1_in_0_ net114 net116 sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_5.mux_l4_in_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk cbx_8__1_.mem_top_ipin_1.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_1.mux_l1_in_2_ sb_8__1_.mux_left_track_15.out net18 cbx_8__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_41_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_28.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_341_ sb_8__1_.mux_top_track_28.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2__A0 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_272_ sb_8__1_.mux_left_track_47.out VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l2_in_2__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input76_A chany_top_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_6.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output232_A net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_44.mux_l3_in_0_ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2_ net62 net70 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xoutput203 net203 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput214 net214 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput225 net225 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
Xoutput247 net247 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
Xoutput236 net236 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_3__385 VGND VGND VPWR VPWR net385 cbx_8__1_.mux_top_ipin_14.mux_l2_in_3__385/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_8_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__322
+ VGND VGND VPWR VPWR net322 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__322/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_left_track_35.mux_l1_in_1__A1 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_27.mux_l1_in_1__350 VGND VGND VPWR VPWR net350 sb_8__1_.mux_left_track_27.mux_l1_in_1__350/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_0.mux_l2_in_3__368 VGND VGND VPWR VPWR net368 sb_8__1_.mux_top_track_0.mux_l2_in_3__368/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__266__A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_324_ sb_8__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_5.mux_l3_in_1_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3_ net265 net87 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_3__257 VGND VGND VPWR VPWR net257 cbx_8__1_.mux_top_ipin_5.mux_l2_in_3__257/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__1_.mem_left_track_9.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_3_ net382 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_59_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_top_track_44.mux_l2_in_1_ net376 sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input39_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_44_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_1__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_307_ sb_8__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_5.mux_l1_in_0_ net54 net78 sb_8__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_25_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_2_ net10 net22 sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4_ net93 net62 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_44.mux_l1_in_2_ net29 net11 sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA__364__A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xinput114 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xinput103 reset_right_in VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_27.mux_l1_in_0_ net61 net91 sb_8__1_.mem_left_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__274__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4__A1 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_3__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_11.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_4__A0 sb_8__1_.mux_left_track_45.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_41.mux_l2_in_0_ net357 sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_41.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__269__A sb_8__1_.mux_left_track_53.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__317
+ VGND VGND VPWR VPWR net317 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__317/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk cbx_8__1_.mem_top_ipin_0.ccff_tail
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_1.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_28.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_340_ net40 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2__A1 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_271_ sb_8__1_.mux_left_track_49.out VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input69_A chany_top_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1_ net39 cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput204 net204 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput226 net226 VGND VGND VPWR VPWR prog_reset_bottom_out sky130_fd_sc_hd__buf_12
Xoutput248 net248 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput237 net237 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_0.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_11_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__372__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_2__S sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_323_ sb_8__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_5.mux_l3_in_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_0__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net288 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_2_ net56 cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_8__1_.mem_left_track_7.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__367__A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_70_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net317 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_2_ net27 sb_8__1_.mux_left_track_35.out cbx_8__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_8__1_.mem_top_ipin_7.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mux_top_track_44.mux_l2_in_0_ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_306_ net66 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_2.mux_l1_in_0__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_1_ net236 net233 sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_12_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__1_.mem_left_track_33.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_29_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3_ net70 net39 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_21_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_top_track_44.mux_l1_in_1_ net23 net38 sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_0__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk cbx_8__1_.mem_top_ipin_3.ccff_tail
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput115 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR
+ VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xinput104 reset_top_in VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_11.mux_l2_in_1__342 VGND VGND VPWR VPWR net342 sb_8__1_.mux_left_track_11.mux_l2_in_1__342/LO
+ sky130_fd_sc_hd__conb_1
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input99_A prog_reset_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_left_track_51.mux_l1_in_1__A1 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__375__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_0__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_4__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input14_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_1__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net284 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__mux2_8
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_31.mux_l1_in_1__353 VGND VGND VPWR VPWR net353 sb_8__1_.mux_left_track_31.mux_l1_in_1__353/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_3__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_1.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_3_ net333 net4 sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_1__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input6_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_20.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_270_ sb_8__1_.mux_left_track_51.out VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_2__A0 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__263 VGND VGND VPWR VPWR net263 cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__263/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xoutput205 net205 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput216 net216 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_10.mem_out\[2\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput227 net227 VGND VGND VPWR VPWR prog_reset_top_out sky130_fd_sc_hd__buf_12
Xoutput249 net249 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
Xoutput238 net238 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
XFILLER_87_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l2_in_3__A1 sb_8__1_.mux_left_track_57.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_41.mux_l1_in_0_ net249 net64 sb_8__1_.mem_left_track_41.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input116_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2__A0 net74 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_322_ sb_8__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_53.mux_l2_in_0_ net363 sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_53.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input81_A chany_top_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__S
+ net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_1_ net7 cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk cbx_8__1_.mem_top_ipin_6.ccff_tail
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_305_ net65 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_bottom_track_21.mux_l3_in_0_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_47.mux_l1_in_0__A0 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_0__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__378__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l1_in_0__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_0_ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk sb_8__1_.mem_left_track_31.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input44_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_29_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2_ net77 net46 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_6.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l1_in_2_ sb_8__1_.mux_left_track_23.out net13 cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_44.mux_l1_in_0_ net119 net111 sb_8__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput116 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR
+ VPWR net116 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput105 sc_in VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_bottom_track_21.mux_l2_in_1_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output248_A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_14.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cbx_8__1_.mem_top_ipin_13.mem_out\[2\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew251 net252 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mux_bottom_track_5.mux_l1_in_1_ net238 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_1__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_2_ net6 net18 sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_1__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_left_track_47.mux_l2_in_0__359 VGND VGND VPWR VPWR net359 sb_8__1_.mux_left_track_47.mux_l2_in_0__359/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_2__A1 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__296__A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_72_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput206 net206 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput217 net217 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xoutput228 net228 VGND VGND VPWR VPWR reset_bottom_out sky130_fd_sc_hd__buf_12
Xoutput239 net239 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_1__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2__A1 net43 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input109_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_321_ net82 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input74_A chany_top_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_55.mux_l1_in_0__A0 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_0__A0 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_top_track_52.mux_l2_in_1__377 VGND VGND VPWR VPWR net377 sb_8__1_.mux_top_track_52.mux_l2_in_1__377/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net306 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_21_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_45.mux_l2_in_1__337 VGND VGND VPWR VPWR net337 sb_8__1_.mux_bottom_track_45.mux_l2_in_1__337/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_74_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_304_ net93 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_4__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_7_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3_ net266 net86 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_1__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_11.mux_l3_in_0_ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_53.mux_l1_in_0_ net247 net80 sb_8__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_13.mux_l1_in_0__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input37_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_43_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_11.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput117 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput106 test_enable_bottom_in VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_21.mux_l2_in_0_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_44_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4_ sb_8__1_.mux_bottom_track_45.out
+ net61 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net298 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__280 VGND VGND VPWR VPWR net280
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__280/LO sky130_fd_sc_hd__conb_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__266 VGND VGND VPWR VPWR net266
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__266/LO sky130_fd_sc_hd__conb_1
XFILLER_90_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_11.mux_l2_in_1_ net342 net248 sb_8__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xload_slew252 net253 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_5.mux_l1_in_0_ net91 net78 sb_8__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.out sky130_fd_sc_hd__clkbuf_2
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__270 VGND VGND VPWR VPWR net270
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__270/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_1__A0 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_1_ net232 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_0__A0 net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3_ net277 net90 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_30_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_25.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.out sky130_fd_sc_hd__clkbuf_2
Xoutput207 net207 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xoutput229 net229 VGND VGND VPWR VPWR reset_left_out sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_1__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_320_ sb_8__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_51.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_51.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input67_A chany_top_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__277 VGND VGND VPWR VPWR net277
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__277/LO sky130_fd_sc_hd__conb_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__292
+ VGND VGND VPWR VPWR net292 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__292/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_21.mux_l1_in_0__A0 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_0__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.out sky130_fd_sc_hd__clkbuf_2
XFILLER_75_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input121_A top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_0__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_303_ sb_8__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2_ net45 cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_0__A0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_13.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_27_prog_clk net389 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_1.mux_l3_in_0_ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2__A0 net77 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_11.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_53_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput118 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND VPWR
+ VPWR net118 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput107 test_enable_right_in VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3_ net69 net38 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_1__A0 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__288
+ VGND VGND VPWR VPWR net288 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__288/LO
+ sky130_fd_sc_hd__conb_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_11.mux_l2_in_0_ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_13.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A0 net66 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_left_track_23.mux_l3_in_0_ sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_23.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_1__A0 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_1.mux_l2_in_1_ net341 sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input97_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_1__S sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_1__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_3__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_0_ net86 net72 sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_11.mux_l2_in_1__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_53.out sky130_fd_sc_hd__buf_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net321 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__mux2_2
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_3_ net387 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_0__A1 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__287
+ VGND VGND VPWR VPWR net287 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__287/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2_ net59 net70 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_11.mux_l1_in_1_ net245 net43 sb_8__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input12_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput208 net208 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_10.ccff_head
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xoutput219 net219 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_bottom_track_45.mux_l3_in_0_ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_3__383 VGND VGND VPWR VPWR net383 cbx_8__1_.mux_top_ipin_12.mux_l2_in_3__383/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_left_track_23.mux_l2_in_1_ net348 net248 sb_8__1_.mem_left_track_23.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2__A0 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.mux_l1_in_2_ net249 net246 sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net106 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_49.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net324 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_47.out sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_3__255 VGND VGND VPWR VPWR net255 cbx_8__1_.mux_top_ipin_3.mux_l2_in_3__255/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_2__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_4_ sb_8__1_.mux_left_track_41.out net33 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_21.mux_l1_in_0__A1 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input114_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_302_ net91 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mux_bottom_track_45.mux_l2_in_1_ net337 net32 sb_8__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net287 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_2.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net295 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_1__A0 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_52_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
XFILLER_10_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_29_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk sb_8__1_.mem_left_track_57.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_2__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_3_ net259 sb_8__1_.mux_left_track_45.out cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_88_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 test_enable_top_in VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput119 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND VPWR
+ VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_10_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input42_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_2.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_12.ccff_tail
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew254 net99 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_16
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_1__A0 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 chany_top_in_0[6] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_4
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_1__A1 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_1.mux_l2_in_0_ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_67_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output246_A net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_9.mux_l2_in_1__367 VGND VGND VPWR VPWR net367 sb_8__1_.mux_left_track_9.mux_l2_in_1__367/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_2_ net27 cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_1_ net39 cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_11.mux_l1_in_0_ net50 net73 sb_8__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_3__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__A1 net89 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net121 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xoutput209 net209 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
XFILLER_67_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_23.mux_l2_in_0_ net34 sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_23.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2__A1 net66 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.mux_l1_in_1_ net243 net52 sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_3__387 VGND VGND VPWR VPWR net387 cbx_8__1_.mux_top_ipin_2.mux_l2_in_3__387/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_3_ net330 net30 sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_378_ net106 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__304
+ VGND VGND VPWR VPWR net304 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__304/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_52_prog_clk
+ sb_8__1_.mem_bottom_track_11.mem_out\[2\] net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_3_ sb_8__1_.mux_left_track_29.out net10 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2_ net77 net46 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_7.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input107_A test_enable_right_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_301_ net90 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_45.mux_l2_in_0_ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_42_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ net99 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input72_A chany_top_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3_ net270 net86 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk sb_8__1_.mem_left_track_25.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_25.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_3.mem_out\[2\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_left_track_15.mux_l2_in_0__A0 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__302__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_1__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_28_prog_clk net388 net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk sb_8__1_.mem_left_track_55.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_57.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_bottom_track_1.mux_l4_in_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_2_ net31 sb_8__1_.mux_left_track_27.out cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput109 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_45.mux_l1_in_1_ net14 net235 sb_8__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4_ sb_8__1_.mux_bottom_track_45.out
+ net61 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input35_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_2.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_2__A0 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_1__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 chany_top_in_0[24] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
Xinput91 chany_top_in_0[7] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
Xcbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_1.mux_l3_in_1_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_sb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__310__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_1__A0 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_1__A0 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.mux_l1_in_0_ net82 net85 sb_8__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net303 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__mux2_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__305__A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_3__A0 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_2_ net12 net24 sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.out sky130_fd_sc_hd__buf_4
X_377_ net106 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_8__1_.mem_bottom_track_11.mem_out\[1\] net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_4.mem_out\[2\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_2_ sb_8__1_.mux_left_track_17.out net17 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_91_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_7.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_300_ net89 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_23.mux_l1_in_0_ net35 net65 sb_8__1_.mem_left_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input65_A chany_top_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_23.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_25.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_2_ net45 cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_35.mux_l2_in_0_ sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_35.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l2_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput1 ccff_head_0_0 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net313 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_2__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_29_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__311
+ VGND VGND VPWR VPWR net311 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__311/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__313__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_1_ net11 cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_45.mux_l1_in_0_ net237 net68 sb_8__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_3_ net383 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net323 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3_ net69 net38 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xoutput190 net190 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_35.mux_l1_in_1_ net355 net246 sb_8__1_.mem_left_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_1__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l2_in_1__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_1__A0 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_2__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__308__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput70 chany_top_in_0[15] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
Xinput81 chany_top_in_0[25] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
Xinput92 chany_top_in_0[8] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__A1 net93 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_1.mux_l3_in_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_7.mux_l1_in_2_ sb_8__1_.mux_left_track_15.out net18 cbx_8__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_90_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_4_ sb_8__1_.mux_left_track_37.out net6 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_1__A0 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_1__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_2.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_1__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input95_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_10.mux_l2_in_3__369 VGND VGND VPWR VPWR net369 sb_8__1_.mux_top_track_10.mux_l2_in_3__369/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_12.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_52.mux_l3_in_0_ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__321__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_3__A1 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_1_ net234 net231 sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_77_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input10_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_376_ net106 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk
+ sb_8__1_.mem_bottom_track_11.mem_out\[0\] net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_3__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_4.mem_out\[1\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__316__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input2_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_10_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_52.mux_l2_in_1_ net377 sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_21.mux_l1_in_3__333 VGND VGND VPWR VPWR net333 sb_8__1_.mux_bottom_track_21.mux_l1_in_3__333/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_3.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_33_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_359_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xinput2 ccff_head_1 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_2__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_0.ccff_tail net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_20_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input112_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_19.mux_l1_in_0__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_2_ net29 cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_52.mux_l1_in_2_ net30 net12 sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_21_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput191 net191 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput180 net180 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_35.mux_l1_in_0_ net56 net86 sb_8__1_.mem_left_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_31.mux_l1_in_1__A1 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_1__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_47.mux_l2_in_0_ net359 sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_47.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__324__A sb_8__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput82 chany_top_in_0[26] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xinput71 chany_top_in_0[16] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
Xinput60 chany_bottom_in[6] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
Xinput93 chany_top_in_0[9] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_0__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input40_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_11.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_7.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_3_ sb_8__1_.mux_left_track_25.out net12 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_10.mux_l2_in_3_ net369 net4 sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l2_in_3__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_1__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_45.mux_l2_in_0__358 VGND VGND VPWR VPWR net358 sb_8__1_.mux_left_track_45.mux_l2_in_0__358/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__D
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input88_A chany_top_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output244_A net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_3__340 VGND VGND VPWR VPWR net340 sb_8__1_.mux_bottom_track_7.mux_l2_in_3__340/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_1.mux_l2_in_0_ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.ccff_tail net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_89_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__275 VGND VGND VPWR VPWR net275
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__275/LO sky130_fd_sc_hd__conb_1
XFILLER_33_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net285 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__mux2_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_375_ net106 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_45_prog_clk
+ sb_8__1_.mem_bottom_track_11.ccff_head net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_4.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net99
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_2.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l2_in_1__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__332__A net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_12.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_10.mux_l4_in_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X sb_8__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_52.mux_l2_in_0_ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_77_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_27.mux_l1_in_0__A0 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_1.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
X_358_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ sb_8__1_.mux_left_track_13.out VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xinput3 ccff_head_2 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_4.mux_l2_in_3_ net375 net33 sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_1.mux_l1_in_1_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__327__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A sc_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input70_A chany_top_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_left_track_19.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_10.mux_l3_in_1_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_52.mux_l1_in_1_ net24 net36 sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_52_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput170 net170 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_14_prog_clk cbx_8__1_.mem_top_ipin_0.mem_out\[2\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire253 net99 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_49_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput72 chany_top_in_0[17] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
Xinput61 chany_bottom_in[7] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_4
Xinput50 chany_bottom_in[24] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
Xinput83 chany_top_in_0[27] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
Xinput94 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__340__A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_top_track_4.mux_l4_in_0_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_8__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.ccff_tail net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input33_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk sb_8__1_.mem_left_track_11.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_7.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_90_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_10.mux_l2_in_2_ net6 net18 sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_1__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__335__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_0__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net304 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_47.mux_l1_in_0_ net244 net67 sb_8__1_.mem_left_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_68_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output237_A net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_17.mux_l2_in_1__A1 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_3__381 VGND VGND VPWR VPWR net381 cbx_8__1_.mux_top_ipin_10.mux_l2_in_3__381/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__296
+ VGND VGND VPWR VPWR net296 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__296/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_4.mux_l3_in_1_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_35.mux_l1_in_0__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_10.mux_l1_in_3_ net59 net44 sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_374_ net106 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A1 net66 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_2.ccff_tail
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk sb_8__1_.mem_left_track_17.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk sb_8__1_.mem_left_track_5.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net314 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__mux2_2
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__301
+ VGND VGND VPWR VPWR net301 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__301/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_27.mux_l1_in_0__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk cbx_8__1_.mem_top_ipin_3.mem_out\[2\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
X_357_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_0__A0 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_4__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_288_ sb_8__1_.mux_left_track_15.out VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_4.mux_l2_in_2_ net16 net61 sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xinput4 chanx_left_in[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_1.mux_l1_in_0_ net65 net82 sb_8__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_49.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__343__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l2_in_3__A1 sb_8__1_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input63_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.out sky130_fd_sc_hd__clkbuf_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\] net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_2__A0 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA__338__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_10.mux_l3_in_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_52.mux_l1_in_0_ net120 net112 sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_3__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__326
+ VGND VGND VPWR VPWR net326 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__326/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput160 net160 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput193 net193 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_14_prog_clk cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3_ net267 net75 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net106 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2__A0 net79 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput40 chany_bottom_in[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
Xinput73 chany_top_in_0[18] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_4
Xinput51 chany_bottom_in[25] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
Xinput62 chany_bottom_in[8] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
Xinput84 chany_top_in_0[28] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
Xinput95 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_15.out sky130_fd_sc_hd__clkbuf_2
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input26_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk sb_8__1_.mem_left_track_11.ccff_head
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_10.mux_l2_in_1_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__351__A net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1__A0 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_6.mem_out\[2\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_0__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_3__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__346__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_4.mux_l3_in_0_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__313
+ VGND VGND VPWR VPWR net313 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__313/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_35.mux_l1_in_0__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_10.mux_l1_in_2_ net120 net118 sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_373_ net124 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input93_A chany_top_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk sb_8__1_.mem_left_track_17.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_17.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_8__1_.mem_left_track_5.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3_ net278 net86 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_8__1_.mem_top_ipin_3.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__buf_2
Xsb_8__1_.mux_left_track_17.mux_l3_in_0_ sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_17.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_356_ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_5.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_287_ sb_8__1_.mux_left_track_17.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_4.mux_l2_in_1_ net48 net120 sb_8__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput5 chanx_left_in[10] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_47.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_43_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input56_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
X_339_ net39 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_2__A1 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4_ sb_8__1_.mux_bottom_track_45.out
+ net61 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_10 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput161 net161 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_left_track_17.mux_l2_in_1_ net345 net245 sb_8__1_.mem_left_track_17.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_14_prog_clk cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input110_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2_ net34 net65 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_57.mux_l2_in_0__365 VGND VGND VPWR VPWR net365 sb_8__1_.mux_left_track_57.mux_l2_in_0__365/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_2__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_51.mux_l1_in_0__A0 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput30 chanx_left_in[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_9.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xinput63 chany_bottom_in[9] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
Xinput52 chany_bottom_in[26] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
Xinput41 chany_bottom_in[16] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput85 chany_top_in_0[29] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
Xinput74 chany_top_in_0[19] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net293 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xinput96 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_3__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_43_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_12.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_10.mux_l2_in_0_ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__325
+ VGND VGND VPWR VPWR net325 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__325/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_7.mux_l2_in_1__366 VGND VGND VPWR VPWR net366 sb_8__1_.mux_left_track_7.mux_l2_in_1__366/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_2
XFILLER_9_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output125_A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_6.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l2_in_2__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__285
+ VGND VGND VPWR VPWR net285 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__285/LO
+ sky130_fd_sc_hd__conb_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_372_ net102 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_10.mux_l1_in_1_ net114 net112 sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input86_A chany_top_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__A1 net75 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_15.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_3_ net255 sb_8__1_.mux_left_track_55.out cbx_8__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_94_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_8__1_.mem_left_track_3.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_2_ net45 cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__D cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__267__A sb_8__1_.mux_left_track_57.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
X_355_ sb_8__1_.mux_top_track_0.out VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_286_ sb_8__1_.mux_left_track_19.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_4.mux_l2_in_0_ net117 sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 chanx_left_in[11] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__329
+ VGND VGND VPWR VPWR net329 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__329/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net296 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__mux2_8
Xsb_8__1_.mux_left_track_7.mux_l3_in_0_ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input49_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ net38 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
X_269_ sb_8__1_.mux_left_track_53.out VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__A1 net63 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3_ net69 net38 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__370__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput140 net140 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput151 net151 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
XFILLER_87_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput173 net173 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_17.mux_l2_in_0_ net37 sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_17.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_14_prog_clk cbx_8__1_.ccff_head
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_1_ net63 cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input103_A reset_right_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_1__A0 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_0__S sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__315
+ VGND VGND VPWR VPWR net315 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__315/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_3.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_7.mux_l2_in_1_ net366 sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_21.out sky130_fd_sc_hd__buf_4
Xinput31 chanx_left_in[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xinput20 chanx_left_in[24] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
Xinput64 chany_top_in_0[0] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xinput42 chany_bottom_in[17] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xinput53 chany_bottom_in[27] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
Xinput86 chany_top_in_0[2] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xinput75 chany_top_in_0[1] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xinput97 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__365__A net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_3__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_41_prog_clk
+ net1 net99 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_0__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_3_ net260 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2_ net74 net43 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_48_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_3.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_29.mux_l1_in_1__A1 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_7.mux_l1_in_2_ net249 net246 sb_8__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input31_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_1__A0 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk cbx_8__1_.mem_top_ipin_6.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_53.mux_l3_in_0_ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_bottom_track_53.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_4_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_371_ net102 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_top_track_10.mux_l1_in_0_ net110 net116 sb_8__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input79_A chany_top_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_4_ sb_8__1_.mux_left_track_41.out net33 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_79_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output235_A net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_2_ net26 sb_8__1_.mux_left_track_37.out cbx_8__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net253 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_8.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4__A0 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk cbx_8__1_.mem_top_ipin_2.ccff_tail
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_53.mux_l2_in_1_ net339 sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_bottom_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_354_ sb_8__1_.mux_top_track_2.out VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_285_ sb_8__1_.mux_left_track_21.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 chanx_left_in[12] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_1__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__368__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_44_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_8__1_.mem_top_track_10.mem_out\[2\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_8__1_.mux_top_track_36.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_268_ sb_8__1_.mux_left_track_55.out VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_19.mux_l2_in_1__346 VGND VGND VPWR VPWR net346 sb_8__1_.mux_left_track_19.mux_l2_in_1__346/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_64_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_12 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_8.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xoutput141 net141 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
XFILLER_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_53.mux_l1_in_2_ net31 net13 sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_87_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_1__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_4.mux_l1_in_0_ net112 net109 sb_8__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3_ net271 net91 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input61_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.out sky130_fd_sc_hd__buf_4
XFILLER_19_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_7.mux_l2_in_0_ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_load_slew251_A net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput10 chanx_left_in[15] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput21 chanx_left_in[25] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xinput43 chany_bottom_in[18] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput54 chany_bottom_in[28] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xinput32 chanx_left_in[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput76 chany_top_in_0[20] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xinput65 chany_top_in_0[10] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
Xinput87 chany_top_in_0[3] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput98 isol_n VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_38_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_37.mux_l1_in_1__A1 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net294 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA__291__A sb_8__1_.mux_left_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_2_ net27 cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk sb_8__1_.mem_left_track_35.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_3_ net331 net26 sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_17.mux_l1_in_0_ net39 net69 sb_8__1_.mem_left_track_17.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__308
+ VGND VGND VPWR VPWR net308 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__308/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk sb_8__1_.mem_bottom_track_53.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_53.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_5.mux_l2_in_1__361 VGND VGND VPWR VPWR net361 sb_8__1_.mux_left_track_5.mux_l2_in_1__361/LO
+ sky130_fd_sc_hd__conb_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__376__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_3.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net329 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net125 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_29.mux_l2_in_0_ sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_7.mux_l1_in_1_ net243 net47 sb_8__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input24_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_14_prog_clk cbx_8__1_.mem_top_ipin_5.ccff_tail
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_12_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_31.mux_l2_in_0_ sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_31.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_81_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_0__A0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_6.mux_l2_in_3__378 VGND VGND VPWR VPWR net378 sb_8__1_.mux_top_track_6.mux_l2_in_3__378/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_3_ net340 net27 sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_50_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_370_ net102 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_3_ sb_8__1_.mux_left_track_29.out net10 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_3_0__leaf_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_37.out sky130_fd_sc_hd__clkbuf_2
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3_ net262 net90 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__273 VGND VGND VPWR VPWR net273
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__273/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_1_ net6 cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_29.mux_l1_in_1_ net351 net243 sb_8__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_bottom_track_11.mux_l4_in_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X sb_8__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_23.mux_l2_in_1__348 VGND VGND VPWR VPWR net348 sb_8__1_.mux_left_track_23.mux_l2_in_1__348/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_53.mux_l2_in_0_ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_353_ sb_8__1_.mux_top_track_4.out VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input91_A chany_top_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_284_ sb_8__1_.mux_left_track_23.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_left_track_31.mux_l1_in_1_ net353 net244 sb_8__1_.mem_left_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_3__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput8 chanx_left_in[13] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_12.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_8__1_.mem_top_track_10.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l4_in_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X sb_8__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__294__A sb_8__1_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ net36 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
X_267_ sb_8__1_.mux_left_track_57.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_3.mux_l1_in_2_ sb_8__1_.mux_left_track_19.out net16 cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_28_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_8.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xoutput142 net142 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_11.mux_l3_in_1_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xoutput153 net153 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_53.mux_l1_in_1_ net25 net236 sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_87_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2__A1 net70 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2_ net60 net68 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input54_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_11.mux_l1_in_1__A0 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_319_ sb_8__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[16] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput22 chanx_left_in[26] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
Xcbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_8__1_.mem_top_ipin_8.ccff_tail
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xinput44 chany_bottom_in[19] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
Xinput55 chany_bottom_in[29] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput33 chanx_left_in[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
Xinput77 chany_top_in_0[21] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
Xinput66 chany_top_in_0[11] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
Xinput88 chany_top_in_0[4] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 prog_reset_bottom_in VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_21.mem_out\[1\] net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_21.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_7.mux_l3_in_1_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_0__A0 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_8__1_.mem_left_track_33.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_2_ net8 net20 sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_3_ net384 sb_8__1_.mux_left_track_57.out cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_7.mux_l1_in_0_ net53 net77 sb_8__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input17_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_2_ net9 net21 sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l1_in_0__A0 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk cbx_8__1_.mem_top_ipin_15.mem_out\[2\]
+ net251 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_2_ sb_8__1_.mux_left_track_17.out net17 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_79_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_3_ net236 net234 sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_3__261 VGND VGND VPWR VPWR net261 cbx_8__1_.mux_top_ipin_9.mux_l2_in_3__261/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__297__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2_ net59 cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_11_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_3.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_39_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_29.mux_l1_in_0_ net60 net90 sb_8__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_54_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input119_A top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_352_ sb_8__1_.mux_top_track_6.out VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_13.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_81_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_283_ sb_8__1_.mux_left_track_25.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input84_A chany_top_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_31.mux_l1_in_0_ net59 net89 sb_8__1_.mem_left_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_3_ net235 net233 sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_68_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2__A0 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 chanx_left_in[14] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_91_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_4__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_12.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_8__1_.mem_top_track_10.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_3__386 VGND VGND VPWR VPWR net386 cbx_8__1_.mux_top_ipin_15.mux_l2_in_3__386/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_335_ net35 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_266_ net84 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_1__A0 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_3.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_2__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_1__A0 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_14 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput143 net143 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_11.mux_l3_in_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xoutput154 net154 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
Xsb_8__1_.mux_bottom_track_53.mux_l1_in_0_ net238 net66 sb_8__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_13.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_1_ net37 cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_2__A0 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_0__A0 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input47_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_6.mux_l2_in_3__258 VGND VGND VPWR VPWR net258 cbx_8__1_.mux_top_ipin_6.mux_l2_in_3__258/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_11.mux_l1_in_1__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_318_ net79 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[17] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput45 chany_bottom_in[1] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_4
Xinput34 chany_bottom_in[0] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput23 chanx_left_in[27] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
Xinput78 chany_top_in_0[22] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
Xinput67 chany_top_in_0[12] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xinput89 chany_top_in_0[5] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XFILLER_6_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput56 chany_bottom_in[2] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__A0 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l3_in_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2__A0 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input101_A prog_reset_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net312 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__290
+ VGND VGND VPWR VPWR net290 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__290/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_8.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_62_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_1_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_2_ net15 net248 cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk sb_8__1_.mem_bottom_track_45.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_2__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_49.mux_l1_in_0__A0 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ net253 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net283 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_1_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1__A0 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_0.mux_l2_in_3_ net368 net31 sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_4.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_3__379 VGND VGND VPWR VPWR net379 cbx_8__1_.mux_top_ipin_0.mux_l2_in_3__379/LO
+ sky130_fd_sc_hd__conb_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_14_prog_clk cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_2_ net232 net238 sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__307
+ VGND VGND VPWR VPWR net307 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__307/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_47_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_351_ net52 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net106 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_282_ sb_8__1_.mux_left_track_27.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input77_A chany_top_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_2_ net231 net237 sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net310 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__320
+ VGND VGND VPWR VPWR net320 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__320/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk sb_8__1_.mem_left_track_21.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_3_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_0__A0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk cbx_8__1_.mem_top_ipin_12.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_10.ccff_head
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_0.mux_l4_in_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ net63 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_1__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
Xcbx_8__1_.mux_top_ipin_3.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__299
+ VGND VGND VPWR VPWR net299 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__299/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_53.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_53.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_1__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xoutput133 net133 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput177 net177 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xoutput188 net188 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
Xcbx_8__1_.mux_top_ipin_13.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk cby_8__1_.cby_8__8_.ccff_tail net254 VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_2__A1 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_0__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_317_ net78 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
Xinput13 chanx_left_in[18] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput46 chany_bottom_in[20] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput35 chany_bottom_in[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput24 chanx_left_in[28] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xinput68 chany_top_in_0[13] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
Xinput79 chany_top_in_0[23] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput57 chany_bottom_in[3] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_13.ccff_tail net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_21.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_55.mux_l2_in_0_ net364 sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_55.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_0__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_0__A0 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_3__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_0.mux_l3_in_1_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_left_track_57.mux_l1_in_0__A0 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_1_ net5 cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail net98 VGND
+ VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__319
+ VGND VGND VPWR VPWR net319 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__319/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_2__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_4__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_2__S sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_37_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xsb_8__1_.mux_bottom_track_7.mux_l2_in_0_ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_25.mux_l1_in_1__349 VGND VGND VPWR VPWR net349 sb_8__1_.mux_left_track_25.mux_l1_in_1__349/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_top_track_0.mux_l2_in_2_ net13 net25 sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_left_track_15.mux_l1_in_0__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk cbx_8__1_.mem_top_ipin_15.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcbx_8__1_.mux_top_ipin_8.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_1_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_1__pin_inpad_0_ sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_13.mux_l1_in_2_ sb_8__1_.mux_left_track_27.out net11 cbx_8__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_20_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_350_ sb_8__1_.mux_top_track_10.out VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_281_ sb_8__1_.mux_left_track_29.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net121 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_1_ left_width_0_height_0_subtile_2__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_21.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_44.mux_l2_in_1__376 VGND VGND VPWR VPWR net376 sb_8__1_.mux_top_track_44.mux_l2_in_1__376/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_3__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_0__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_8__1_.mem_top_ipin_11.ccff_tail
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__264 VGND VGND VPWR VPWR net264 cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__264/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ sb_8__1_.mux_top_track_44.out VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_bottom_track_37.mux_l2_in_1__336 VGND VGND VPWR VPWR net336 sb_8__1_.mux_bottom_track_37.mux_l2_in_1__336/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l2_in_1__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_51.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput134 net134 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput178 net178 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net315 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__mux2_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_left_track_55.mux_l2_in_0__364 VGND VGND VPWR VPWR net364 sb_8__1_.mux_left_track_55.mux_l2_in_0__364/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_316_ net77 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chany_bottom_in[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
Xinput14 chanx_left_in[19] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 chanx_left_in[29] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xinput69 chany_top_in_0[14] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xinput47 chany_bottom_in[21] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput58 chany_bottom_in[4] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_23_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__316
+ VGND VGND VPWR VPWR net316 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__316/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_1__A0 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_0__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_0.mux_l3_in_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2__A0 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l2_in_1__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input52_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__300__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_23.mux_l1_in_0__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_3__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_0__A0 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3_ net274 net90 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_0__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_13.mux_l3_in_0_ sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_55.mux_l1_in_0_ net248 net81 sb_8__1_.mem_left_track_55.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net301 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_0.mux_l2_in_1_ net35 net52 sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_4.mux_l2_in_3__375 VGND VGND VPWR VPWR net375 sb_8__1_.mux_top_track_4.mux_l2_in_3__375/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net299 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_left_track_15.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_8__1_.mem_top_ipin_14.ccff_tail
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_2__A0 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail net98 VGND
+ VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_11.mux_l1_in_0_ net89 net74 sb_8__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_13.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input15_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk sb_8__1_.mem_top_track_0.mem_out\[2\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input7_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l2_in_1__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_13.mux_l2_in_1_ net343 net243 sb_8__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ sb_8__1_.mux_left_track_31.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_7.mux_l1_in_0_ net90 net77 sb_8__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A0 net93 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk sb_8__1_.mem_left_track_19.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l2_in_1__A0 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.out sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input117_A top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_332_ net61 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A chany_top_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 net105 net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_11.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\] net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput124 net124 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3_ net279 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput146 net146 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
XANTENNA__303__A sb_8__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput168 net168 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput179 net179 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_13.mux_l2_in_1__A1 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_315_ sb_8__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput26 chanx_left_in[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_left_in[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput37 chany_bottom_in[12] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput48 chany_bottom_in[22] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xinput59 chany_bottom_in[5] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
XANTENNA_sb_8__1_.mux_left_track_31.mux_l1_in_0__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_27.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_27.out sky130_fd_sc_hd__clkbuf_2
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_0__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_1__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2__A1 net70 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk sb_8__1_.mem_left_track_27.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_27.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_75_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk sb_8__1_.mem_bottom_track_5.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk sb_8__1_.mem_bottom_track_45.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input45_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_23.mux_l1_in_0__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l2_in_2__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_1.mux_l1_in_0__A0 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2_ net59 cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output249_A net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_12_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_0.mux_l2_in_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_15_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__323
+ VGND VGND VPWR VPWR net323 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__323/LO
+ sky130_fd_sc_hd__conb_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_3.mux_l3_in_0_ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__281 VGND VGND VPWR VPWR net281
+ cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__281/LO sky130_fd_sc_hd__conb_1
XFILLER_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__267 VGND VGND VPWR VPWR net267
+ cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__267/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_2__A1 net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_13.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND
+ VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_2__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__271 VGND VGND VPWR VPWR net271
+ cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__271/LO sky130_fd_sc_hd__conb_1
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_8__1_.mem_top_track_0.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__306__A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_13.mux_l2_in_0_ net42 sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_0.mux_l1_in_1_ net118 net113 sb_8__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_21.mux_l2_in_1__A1 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.mux_l2_in_1_ net352 sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_1__A0 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_28.mux_l1_in_3_ net373 net27 sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ net60 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_46_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input75_A chany_top_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output231_A net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_left_track_17.mux_l2_in_1__345 VGND VGND VPWR VPWR net345 sb_8__1_.mux_left_track_17.mux_l2_in_1__345/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_3_ net256 sb_8__1_.mux_left_track_57.out cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput125 net125 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2_ net57 net68 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xoutput147 net147 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput169 net169 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_3__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__278 VGND VGND VPWR VPWR net278
+ cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__278/LO sky130_fd_sc_hd__conb_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_8__1_.mem_bottom_track_13.mem_out\[1\] net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__A1 net87 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk sb_8__1_.mem_top_track_6.mem_out\[2\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_55.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_55.out sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_3.mux_l1_in_2_ net250 net247 sb_8__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_314_ net74 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__302
+ VGND VGND VPWR VPWR net302 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__302/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput27 chanx_left_in[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
Xinput16 chanx_left_in[20] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_52_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput49 chany_bottom_in[23] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_4
Xinput38 chany_bottom_in[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_31.mux_l1_in_0__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__268 VGND VGND VPWR VPWR net268
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__268/LO sky130_fd_sc_hd__conb_1
XFILLER_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net297 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__mux2_8
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__314__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk sb_8__1_.mem_left_track_25.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_27.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_37.mux_l1_in_1__356 VGND VGND VPWR VPWR net356 sb_8__1_.mux_left_track_37.mux_l1_in_1__356/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk sb_8__1_.mem_bottom_track_5.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_45.mem_out\[0\] net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_45.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_bottom_track_11.mux_l2_in_3__331 VGND VGND VPWR VPWR net331 sb_8__1_.mux_bottom_track_11.mux_l2_in_3__331/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input38_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_4_ sb_8__1_.mux_left_track_45.out net31 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_74_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_2__S sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mux_top_track_28.mux_l3_in_0_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__309__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_49.out sky130_fd_sc_hd__clkbuf_2
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_12_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net319 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_28.mux_l2_in_1_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_28_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
Xcbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_3.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_3_ net261 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_5_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_1__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1__A0 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk sb_8__1_.mem_top_track_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_4.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_36_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_left_track_21.mux_l2_in_1__347 VGND VGND VPWR VPWR net347 sb_8__1_.mux_left_track_21.mux_l2_in_1__347/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_top_track_0.mux_l1_in_0_ net110 net115 sb_8__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_41_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input20_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.mux_l2_in_0_ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_1__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__317__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_28.mux_l1_in_2_ net9 net21 sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l2_in_2__A0 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l2_in_2__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_330_ net59 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_13.mux_l2_in_3__384 VGND VGND VPWR VPWR net384 cbx_8__1_.mux_top_ipin_13.mux_l2_in_3__384/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input68_A chany_top_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_2_ net15 cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_1_ net37 cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xoutput126 net126 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xsb_8__1_.mux_left_track_13.mux_l1_in_0_ net46 net72 sb_8__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_top_track_10.mux_l1_in_3__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_1.mux_l2_in_3__380 VGND VGND VPWR VPWR net380 cbx_8__1_.mux_top_ipin_1.mux_l2_in_3__380/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_9.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_8__1_.mem_top_track_6.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_25.mux_l2_in_0_ sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_25.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input122_A top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_3.mux_l1_in_1_ net244 net49 sb_8__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_14_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_3__256 VGND VGND VPWR VPWR net256 cbx_8__1_.mux_top_ipin_4.mux_l2_in_3__256/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_313_ net73 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 chanx_left_in[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput17 chanx_left_in[21] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput39 chany_bottom_in[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_69_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_3_ net335 net29 sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__330__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_45_prog_clk sb_8__1_.mem_bottom_track_5.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_37.ccff_tail net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_45.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l1_in_3__A0 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__300
+ VGND VGND VPWR VPWR net300 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__300/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_3_ sb_8__1_.mux_left_track_33.out net8 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2_ net74 net43 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_2.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_8_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net326 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__mux2_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_9.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_25.mux_l1_in_1_ net349 net249 sb_8__1_.mem_left_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3_ net272 net90 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input50_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_12_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_2.mux_l2_in_3__371 VGND VGND VPWR VPWR net371 sb_8__1_.mux_top_track_2.mux_l2_in_3__371/LO
+ sky130_fd_sc_hd__conb_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_28.mux_l2_in_0_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input98_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_3.mux_l4_in_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_8__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_2_ net29 sb_8__1_.mux_left_track_31.out cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_8__1_.mem_top_track_52.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk net3
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_45_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] net252 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_4.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk sb_8__1_.mem_left_track_13.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_8__1_.mem_left_track_1.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input13_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l2_in_1__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_0.mux_l1_in_3__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_wire253_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__A1 net91 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_28.mux_l1_in_1_ net45 net40 sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_45.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_13.mux_l2_in_2__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input5_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_3.mux_l3_in_1_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A0 sb_8__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3_ net263 net89 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__S cby_8__1_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_5.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__1_.mux_left_track_25.mux_l1_in_1__A1 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput127 net127 VGND VGND VPWR VPWR ccff_tail_1 sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_1__A0 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__328__A net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__312
+ VGND VGND VPWR VPWR net312 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__312/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk
+ sb_8__1_.mem_bottom_track_11.ccff_tail net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_8__1_.mem_top_track_6.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_86_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input115_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_3.mux_l1_in_0_ net55 net79 sb_8__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_312_ net72 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input80_A chany_top_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[22] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xinput29 chanx_left_in[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_1__A0 sb_8__1_.mux_left_track_9.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_2_ net11 net23 sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_3.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_3__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4_ net66 net35 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__1_.cby_8__8_.mux_left_ipin_0.out cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_78_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_2_ sb_8__1_.mux_left_track_21.out net14 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_47_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1_ sb_8__1_.mux_bottom_track_11.out
+ net50 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__286
+ VGND VGND VPWR VPWR net286 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__286/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l2_in_3__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_49.mux_l2_in_0__360 VGND VGND VPWR VPWR net360 sb_8__1_.mux_left_track_49.mux_l2_in_0__360/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__1_.mux_top_ipin_9.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_41.mux_l2_in_0__357 VGND VGND VPWR VPWR net357 sb_8__1_.mux_left_track_41.mux_l2_in_0__357/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_16_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_25.mux_l1_in_0_ net63 net93 sb_8__1_.mem_left_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net106 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2_ net59 cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_55_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_37.mux_l2_in_0_ sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_20_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_20.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input43_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_12_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_2__S sb_8__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk cbx_8__1_.mem_top_ipin_2.mem_out\[2\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__1_.mux_top_ipin_9.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_7.mux_l2_in_2__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__336__A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mux_bottom_track_13.mux_l1_in_1__S sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_1_ net9 cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_8__1_.mem_top_track_52.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output247_A net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_3_ net385 sb_8__1_.mux_left_track_53.out cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_44_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_8.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk sb_8__1_.mem_left_track_13.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_37.mux_l1_in_1_ net356 net247 sb_8__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk sb_8__1_.mem_left_track_1.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_33.mux_l1_in_1__A1 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__324
+ VGND VGND VPWR VPWR net324 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__324/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_28.mux_l1_in_0_ net117 net109 sb_8__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_14_prog_clk sb_8__1_.mem_left_track_41.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__262 VGND VGND VPWR VPWR net262 cby_8__1_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__262/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_bottom_track_3.mux_l3_in_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_20.mux_l1_in_3__372 VGND VGND VPWR VPWR net372 sb_8__1_.mux_top_track_20.mux_l1_in_3__372/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_9.mux_l1_in_2_ sb_8__1_.mux_left_track_19.out net16 cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_4_ sb_8__1_.mux_left_track_41.out net33 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2_ net58 cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_12_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_4.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_40_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l2_in_3__A1 sb_8__1_.mux_left_track_45.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_3__332 VGND VGND VPWR VPWR net332 sb_8__1_.mux_bottom_track_13.mux_l1_in_3__332/LO
+ sky130_fd_sc_hd__conb_1
Xoutput128 net128 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__1_.mux_left_track_3.mux_l1_in_1__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_21.mux_l1_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__344__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_8__1_.mem_top_track_4.ccff_tail
+ net254 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_14.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_86_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input108_A test_enable_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_311_ sb_8__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk sb_8__1_.mem_left_track_19.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 chanx_left_in[23] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A chany_top_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_8__1_.mem_left_track_7.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net316 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_1_ net235 net232 sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk cbx_8__1_.mem_top_ipin_5.mem_out\[2\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__339__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3_ net72 net41 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_1_ sb_8__1_.mux_left_track_9.out net21 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0_ sb_8__1_.mux_bottom_track_5.out
+ net53 cby_8__1_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_3.mux_l2_in_1__352 VGND VGND VPWR VPWR net352 sb_8__1_.mux_left_track_3.mux_l2_in_1__352/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_14.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_32_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net308 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__mux2_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_20.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_left_track_29.mux_l1_in_0__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input36_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk cbx_8__1_.mem_top_ipin_2.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_9.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_44.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2__A1 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_2_ net27 cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__293
+ VGND VGND VPWR VPWR net293 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__293/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_top_track_10.mux_l2_in_1__S sb_8__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__1_.mem_left_track_11.ccff_tail
+ net252 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_left_track_37.mux_l1_in_0_ net45 net75 sb_8__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__347__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_8__1_.mem_bottom_track_53.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_49.mux_l2_in_0_ net360 sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_49.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_51.mux_l2_in_0_ sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_51.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_9.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_8.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_3_ sb_8__1_.mux_left_track_29.out net10 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_12_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput129 net129 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_35_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_0__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_53.mux_l2_in_0__363 VGND VGND VPWR VPWR net363 sb_8__1_.mux_left_track_53.mux_l2_in_0__363/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ net70 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk sb_8__1_.mem_left_track_19.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_19.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_0__A0 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input66_A chany_top_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_37.mem_out\[1\] net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_37.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_left_track_19.mux_l2_in_1__A1 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk sb_8__1_.mem_left_track_7.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_51.mux_l1_in_1_ net362 net250 sb_8__1_.mem_left_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_0_ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_83_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2_ net79 net48 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_37.mux_l1_in_0__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_4.mux_l1_in_2__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_4.mux_l1_in_0_ sb_8__1_.mux_left_track_3.out net24 cbx_8__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input120_A top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xcbx_8__1_.mux_top_ipin_14.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_12.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__1_.mux_left_track_29.mux_l1_in_0__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_6.mux_l2_in_3_ net378 net5 sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input29_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_0__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_3.mux_l1_in_1_ net237 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l1_in_4__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk cbx_8__1_.mem_top_ipin_2.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_15.mux_l2_in_3__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net106 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__283
+ VGND VGND VPWR VPWR net283 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__283/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_2.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__273__A sb_8__1_.mux_left_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input96_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2__A0 net77 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_6.mux_l4_in_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_8__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__310
+ VGND VGND VPWR VPWR net310 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__310/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net305 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_9.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_8.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net282 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_2_ sb_8__1_.mux_left_track_17.out net17 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_12_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input11_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_4__A0 sb_8__1_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_45.mux_l1_in_0__A0 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__276 VGND VGND VPWR VPWR net276
+ cby_8__1_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__276/LO sky130_fd_sc_hd__conb_1
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l2_in_2__A0 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_49.mux_l1_in_0_ net245 net71 sb_8__1_.mem_left_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input3_A ccff_head_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l2_in_1__A0 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk sb_8__1_.mem_left_track_17.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_42_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_0.mux_l1_in_0__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input59_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_37.mem_out\[0\] net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_37.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_8__1_.mem_left_track_5.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_51.mux_l1_in_0_ net246 net76 sb_8__1_.mem_left_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_6.mux_l3_in_1_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_8__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_369_ net102 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_8__1_.mem_top_ipin_5.mem_out\[0\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_56_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_12.mux_l1_in_3_ net370 net15 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__371__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_37.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input113_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_1__S sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_bottom_track_29.mux_l3_in_0_ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__1_.mem_left_track_31.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__366__A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_bottom_track_5.mux_l2_in_3__338 VGND VGND VPWR VPWR net338 sb_8__1_.mux_bottom_track_5.mux_l2_in_3__338/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__295
+ VGND VGND VPWR VPWR net295 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__295/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_top_track_6.mux_l2_in_2_ net17 net60 sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_59_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_left_track_7.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_3.mux_l1_in_0_ net93 net79 sb_8__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__276__A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk cbx_8__1_.mem_top_ipin_1.ccff_tail
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net290 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__mux2_4
XFILLER_61_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_29.mux_l2_in_1_ net334 sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_bottom_track_29.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__305
+ VGND VGND VPWR VPWR net305 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__305/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input41_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_14.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_12.mux_l3_in_0_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_23.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_23.out sky130_fd_sc_hd__clkbuf_2
XFILLER_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_54_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ cby_8__1_.cby_8__8_.mem_left_ipin_1.ccff_tail net251 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3_ net275 sb_8__1_.mux_bottom_track_45.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input89_A chany_top_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_12.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output245_A net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_left_track_53.mux_l1_in_0__A0 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_29.mux_l1_in_2_ net5 net17 sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_66_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_8.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__374__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_17.out sky130_fd_sc_hd__clkbuf_2
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_12.mux_l2_in_1_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_11.mux_l2_in_3__382 VGND VGND VPWR VPWR net382 cbx_8__1_.mux_top_ipin_11.mux_l2_in_3__382/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__1_.mux_left_track_5.mux_l2_in_1__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_head net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__297
+ VGND VGND VPWR VPWR net297 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__297/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_left_track_15.mux_l2_in_1__344 VGND VGND VPWR VPWR net344 sb_8__1_.mux_left_track_15.mux_l2_in_1__344/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l1_in_4__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_2__S sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__369__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_8__1_.mem_bottom_track_29.ccff_tail net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_37.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_6.mux_l3_in_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_368_ net102 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_51_prog_clk net2 net252 VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_2
X_299_ sb_8__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l2_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_4.ccff_tail
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_56_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_top_track_12.mux_l1_in_2_ net7 net19 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_35.mux_l1_in_1__355 VGND VGND VPWR VPWR net355 sb_8__1_.mux_left_track_35.mux_l1_in_1__355/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_59_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input106_A test_enable_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__A1 sb_8__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_10.mux_l2_in_3__A1 sb_8__1_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input71_A chany_top_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3_ net280 net90 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__S cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk sb_8__1_.mem_left_track_29.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_19.mux_l3_in_0_ sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_19.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mux_bottom_track_53.mux_l2_in_1__339 VGND VGND VPWR VPWR net339 sb_8__1_.mux_bottom_track_53.mux_l2_in_1__339/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__1_.mux_top_track_6.mux_l2_in_1_ net47 sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_21.mux_l3_in_0_ sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sb_8__1_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk sb_8__1_.mem_top_track_44.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__327
+ VGND VGND VPWR VPWR net327 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__327/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2__A0 sb_8__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__377__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__1_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_51.out sky130_fd_sc_hd__clkbuf_2
XFILLER_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_29.mux_l2_in_0_ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4_ sb_8__1_.mux_bottom_track_37.out
+ net36 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_12.ccff_tail net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input34_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_8__1_.mem_top_ipin_11.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__1_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_0_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_3_ net379 sb_8__1_.mux_left_track_49.out cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_19.mux_l2_in_1_ net346 net246 sb_8__1_.mem_left_track_19.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2_ net61 net72 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_top_track_6.mux_l1_in_2_ net119 net117 sb_8__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_28_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_14_prog_clk sb_8__1_.mem_left_track_37.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_left_track_21.mux_l2_in_1_ net347 net247 sb_8__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output238_A net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_bottom_track_29.mux_l1_in_1_ net233 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__1_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk cbx_8__1_.mem_top_ipin_7.ccff_tail
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__1_.mux_top_ipin_6.mux_l1_in_3__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_14.mux_l1_in_0_ sb_8__1_.mux_left_track_5.out net23 cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net300 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_12.mux_l2_in_0_ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_4_ sb_8__1_.mux_left_track_37.out net6 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_13_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_0__A0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_0__A0 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_35_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_42_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_1__A0 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_0.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_left_track_11.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__306
+ VGND VGND VPWR VPWR net306 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__306/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_367_ net254 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ net87 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__A0 net79 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_12.mux_l1_in_1_ net57 net43 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A0 net82 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net286 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_34_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input64_A chany_top_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_3_ net257 net84 cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_77_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_37_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2_ net59 cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_8_prog_clk cbx_8__1_.mem_top_ipin_14.mem_out\[2\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_12.mem_out\[1\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_load_slew254_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_35_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_0.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__D sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_50_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__1_.mux_top_track_6.mux_l2_in_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_1__A0 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__1_.mux_left_track_9.mux_l3_in_0_ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk sb_8__1_.mem_top_track_44.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_0__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2__A1 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3_ net73 net42 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_8__1_.mem_top_ipin_11.mem_out\[1\]
+ net252 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input27_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_2_ net29 cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_19.mux_l2_in_0_ net62 sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_19.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1_ net41 cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_1__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_6.mux_l1_in_1_ net113 net111 sb_8__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_51.mux_l1_in_1__362 VGND VGND VPWR VPWR net362 sb_8__1_.mux_left_track_51.mux_l1_in_1__362/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_5.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk sb_8__1_.mem_left_track_35.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mux_left_track_21.mux_l2_in_0_ net58 sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_9.mux_l2_in_1_ net367 sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_left_track_9.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__298__A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__mux2_1
XFILLER_71_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 cbx_8__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__1_.mux_bottom_track_29.mux_l1_in_0_ net75 net70 sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__1_.mux_bottom_track_29.mux_l1_in_1__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__318
+ VGND VGND VPWR VPWR net318 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__318/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_1.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_3_ sb_8__1_.mux_left_track_25.out net12 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_4__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input94_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2_ net79 net48 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output250_A net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__1_.mux_top_ipin_5.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk0_A clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_9.mux_l1_in_2_ net250 net247 sb_8__1_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_24_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3_ net268 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_left_track_9.mux_l1_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_366_ net254 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_297_ net86 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mux_top_track_12.mux_l1_in_0_ net113 net115 sb_8__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_20.mux_l1_in_3__S sb_8__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_2__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input1_A ccff_head_0_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input57_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_2_ net4 sb_8__1_.mux_left_track_41.out cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_37_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_14.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_12.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_36.mux_l3_in_0_ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_8__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
X_349_ sb_8__1_.mux_top_track_12.out VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4_ net65 net63 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_52_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__A1 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput250 net250 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_3.mux_l1_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input111_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_1.mux_l2_in_1__A1 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_14.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_1__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk sb_8__1_.mem_top_track_36.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net122 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2_ sb_8__1_.mux_bottom_track_13.out
+ net49 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_top_track_36.mux_l2_in_1_ net374 sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_8__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net327 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__mux2_4
XFILLER_87_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_11.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_1_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__A1 net90 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_bottom_track_37.mux_l1_in_1__A1 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_6.mux_l1_in_0_ net109 net115 sb_8__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3_ net273 net89 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_29_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2__A1 net68 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_9.mux_l2_in_0_ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_8__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 cby_8__1_.cby_8__8_.mux_left_ipin_2.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net253
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_top_track_36.mux_l1_in_2_ net28 net10 sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net318 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_2_ sb_8__1_.mux_left_track_13.out net19 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_13_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_19.mux_l1_in_0_ net38 net68 sb_8__1_.mem_left_track_19.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input87_A chany_top_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1_ net82 net51 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_0__S sb_8__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output243_A net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_8__1_.mem_bottom_track_29.mem_out\[1\] net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_29.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__1_.mux_top_ipin_5.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_8__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__1_.mux_left_track_21.mux_l1_in_0_ net36 net66 sb_8__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_9.mux_l1_in_1_ net244 net44 sb_8__1_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_left_track_13.mux_l2_in_0__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_2_ net57 cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_45.out sky130_fd_sc_hd__buf_4
XFILLER_54_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_33.mux_l2_in_0_ sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_left_track_33.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net289 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
X_365_ net252 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
X_296_ net75 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__A0 net73 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_0__A0 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1__A0 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3_ net264 sb_8__1_.mux_bottom_track_53.out
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk sb_8__1_.mem_left_track_23.mem_out\[1\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_23.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_1__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_1_ net33 cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__1_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_37_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l2_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_3_ net381 sb_8__1_.mux_left_track_57.out cbx_8__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_14.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_8__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_8__1_.mem_top_track_10.ccff_tail
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_348_ net49 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_279_ sb_8__1_.mux_left_track_33.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3_ sb_8__1_.mux_bottom_track_29.out
+ net40 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_28.mux_l1_in_2__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_0.mux_l2_in_1__S sb_8__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_33.mux_l1_in_1_ net354 net245 sb_8__1_.mem_left_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xoutput240 net240 VGND VGND VPWR VPWR test_enable_bottom_out sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk sb_8__1_.mem_left_track_55.mem_out\[0\]
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_55.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__1_.mux_bottom_track_3.mux_l2_in_3__335 VGND VGND VPWR VPWR net335 sb_8__1_.mux_bottom_track_3.mux_l2_in_3__335/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input104_A reset_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_30_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net99 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfrtp_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__1_.mux_bottom_track_45.mux_l1_in_1__A1 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net322 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4_ net65 net63 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l1_in_4__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_5.mux_l1_in_2_ sb_8__1_.mux_left_track_23.out net13 cbx_8__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1_ sb_8__1_.mux_bottom_track_7.out
+ net52 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_1__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_4_ sb_8__1_.mux_left_track_45.out net31 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_top_track_36.mux_l2_in_0_ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_8__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk cbx_8__1_.mem_top_ipin_10.ccff_tail
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_1__A0 net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l4_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_8__1_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_1__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2_ net58 net66 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_43_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__328
+ VGND VGND VPWR VPWR net328 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__328/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_8__1_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input32_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__309
+ VGND VGND VPWR VPWR net309 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__309/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net252 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_8.mux_l2_in_3__A1 sb_8__1_.mux_left_track_53.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3__A0 net70 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_3 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mux_left_track_21.mux_l2_in_0__A0 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_0__A0 sb_8__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_36.mux_l1_in_1_ net22 net39 sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net124 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net106 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__sdfrtp_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_13_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__1_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_1_ sb_8__1_.mux_left_track_7.out net22 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_3_ net386 net88 cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_80_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l3_in_1_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_2__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0_ sb_8__1_.mux_bottom_track_3.out
+ net54 cby_8__1_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output236_A net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__D sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_8__1_.mem_bottom_track_29.mem_out\[0\] net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_29.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__1_.mux_top_ipin_10.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_8__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_9.mux_l1_in_0_ net51 net74 sb_8__1_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__274 VGND VGND VPWR VPWR net274
+ cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__274/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_29_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__1_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_34_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_2.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l2_in_1_ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_bottom_track_3.mux_l2_in_2__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_364_ net99 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
X_295_ sb_8__1_.mux_left_track_1.out VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net251 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net254 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__1_.mux_top_track_36.mux_l1_in_2__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__1_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net102 grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net106 VGND
+ VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_6.mux_l1_in_0__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_bottom_track_13.mux_l1_in_3_ net332 net15 sb_8__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_59_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l2_in_2_ net57 cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__1_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk sb_8__1_.mem_left_track_23.mem_out\[0\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_23.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net253 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk sb_8__1_.mem_bottom_track_1.mem_out\[2\]
+ net253 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__1_.mux_bottom_track_53.mux_l1_in_1__A1 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_5.mux_l2_in_0_ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_8__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_37_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk cbx_8__1_.mem_top_ipin_13.ccff_tail
+ net253 VGND VGND VPWR VPWR cbx_8__1_.mem_top_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_35_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_10.mux_l2_in_2_ net15 cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__1_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_347_ net48 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
Xsb_8__1_.mux_left_track_1.mux_l2_in_1__341 VGND VGND VPWR VPWR net341 sb_8__1_.mux_left_track_1.mux_l2_in_1__341/LO
+ sky130_fd_sc_hd__conb_1
X_278_ sb_8__1_.mux_left_track_35.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xcby_8__1_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2_ net78 net47 cby_8__1_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_38_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__1_.mux_top_ipin_5.mux_l2_in_1__A0 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_15.mux_l4_in_0_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X net126 VGND VGND VPWR VPWR
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mux_left_track_33.mux_l1_in_0_ net57 net87 sb_8__1_.mem_left_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput230 net230 VGND VGND VPWR VPWR reset_top_out sky130_fd_sc_hd__buf_12
Xoutput241 net241 VGND VGND VPWR VPWR test_enable_left_out sky130_fd_sc_hd__buf_12
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__1_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk sb_8__1_.mem_left_track_53.ccff_tail
+ net251 VGND VGND VPWR VPWR sb_8__1_.mem_left_track_55.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__1_.mux_left_track_45.mux_l2_in_0_ net358 sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__1_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR sb_8__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_left_track_29.mux_l1_in_1__351 VGND VGND VPWR VPWR net351 sb_8__1_.mux_left_track_29.mux_l1_in_1__351/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input62_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_load_slew252_A net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__289
+ VGND VGND VPWR VPWR net289 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__289/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3_ sb_8__1_.mux_bottom_track_29.out
+ net40 cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net254 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_33_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__301__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_5.mux_l1_in_1_ sb_8__1_.mux_left_track_11.out net20 cbx_8__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0_ sb_8__1_.mux_bottom_track_1.out
+ net55 cby_8__1_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_bottom_track_11.mux_l1_in_1__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__1_.mux_top_ipin_10.mux_l1_in_3_ sb_8__1_.mux_left_track_33.out net8 cbx_8__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__1_.mux_bottom_track_5.mux_l1_in_1__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__1_.mux_bottom_track_13.mux_l3_in_0_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X sb_8__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_8__1_.mux_top_ipin_15.mux_l3_in_1_ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__1_.mux_top_track_4.mux_l2_in_1__A1 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1_ net35 cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net309 grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__mux2_4
Xclkbuf_leaf_38_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ cby_8__1_.cby_8__8_.mem_right_ipin_5.mem_out\[2\] net253 VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mem_right_ipin_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_52.mux_l1_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cby_8__1_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__1_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_4 net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__1_.mux_top_track_12.mux_l1_in_0__A0 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__1_.mux_top_track_2.mux_l2_in_3__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__1_.mux_top_ipin_7.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__1_.mux_top_track_36.mux_l1_in_0_ net118 net110 sb_8__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net251 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_0.mux_l1_in_0_ sb_8__1_.mux_left_track_1.out net25 cbx_8__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mux_bottom_track_13.mux_l2_in_1_ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sb_8__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__1_.mux_top_ipin_15.mux_l2_in_2_ net32 sb_8__1_.mux_left_track_31.out cbx_8__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_8__1_.cby_8__8_.mux_left_ipin_2.mux_l3_in_0_ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__1_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__1_.mux_top_track_44.mux_l1_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__1_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2_ sb_8__1_.mux_bottom_track_21.out
+ net44 cby_8__1_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__1_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ sb_8__1_.mem_bottom_track_21.ccff_tail net252 VGND VGND VPWR VPWR sb_8__1_.mem_bottom_track_29.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__1_.mux_top_ipin_10.mux_l3_in_0_ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_8__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_29_prog_clk grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net99 VGND VGND VPWR VPWR grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
.ends

