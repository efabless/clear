magic
tech sky130A
magscale 1 2
timestamp 1625782874
<< locali >>
rect 8493 17187 8527 17289
rect 9965 16575 9999 16745
rect 9873 5627 9907 5729
rect 9447 5321 9539 5355
rect 9505 5151 9539 5321
<< viali >>
rect 1869 17289 1903 17323
rect 2973 17289 3007 17323
rect 3985 17289 4019 17323
rect 8493 17289 8527 17323
rect 8677 17289 8711 17323
rect 9321 17289 9355 17323
rect 11345 17289 11379 17323
rect 12725 17289 12759 17323
rect 1409 17221 1443 17255
rect 3249 17221 3283 17255
rect 4261 17221 4295 17255
rect 4813 17221 4847 17255
rect 5181 17221 5215 17255
rect 5641 17221 5675 17255
rect 6009 17221 6043 17255
rect 6561 17221 6595 17255
rect 6929 17221 6963 17255
rect 7297 17221 7331 17255
rect 7757 17221 7791 17255
rect 8125 17221 8159 17255
rect 10241 17221 10275 17255
rect 10517 17221 10551 17255
rect 13185 17221 13219 17255
rect 15669 17221 15703 17255
rect 2513 17153 2547 17187
rect 8493 17153 8527 17187
rect 9597 17153 9631 17187
rect 13001 17153 13035 17187
rect 13829 17153 13863 17187
rect 2145 17085 2179 17119
rect 2329 17085 2363 17119
rect 7113 17085 7147 17119
rect 8769 17085 8803 17119
rect 10149 17085 10183 17119
rect 10425 17085 10459 17119
rect 10701 17085 10735 17119
rect 10977 17085 11011 17119
rect 11253 17085 11287 17119
rect 11529 17085 11563 17119
rect 12081 17085 12115 17119
rect 12357 17085 12391 17119
rect 12633 17085 12667 17119
rect 12909 17085 12943 17119
rect 13369 17085 13403 17119
rect 13737 17085 13771 17119
rect 14197 17085 14231 17119
rect 14749 17085 14783 17119
rect 15025 17085 15059 17119
rect 15301 17085 15335 17119
rect 1593 17017 1627 17051
rect 1961 17017 1995 17051
rect 2697 17017 2731 17051
rect 3065 17017 3099 17051
rect 3433 17017 3467 17051
rect 4077 17017 4111 17051
rect 4445 17017 4479 17051
rect 4997 17017 5031 17051
rect 5365 17017 5399 17051
rect 5825 17017 5859 17051
rect 6193 17017 6227 17051
rect 6745 17017 6779 17051
rect 7481 17017 7515 17051
rect 7941 17017 7975 17051
rect 8309 17017 8343 17051
rect 9413 17017 9447 17051
rect 9781 17017 9815 17051
rect 11713 17017 11747 17051
rect 14289 17017 14323 17051
rect 15485 17017 15519 17051
rect 9965 16949 9999 16983
rect 10793 16949 10827 16983
rect 11069 16949 11103 16983
rect 11897 16949 11931 16983
rect 12173 16949 12207 16983
rect 12449 16949 12483 16983
rect 13553 16949 13587 16983
rect 14013 16949 14047 16983
rect 14565 16949 14599 16983
rect 14841 16949 14875 16983
rect 15117 16949 15151 16983
rect 1593 16745 1627 16779
rect 9965 16745 9999 16779
rect 10057 16745 10091 16779
rect 11253 16745 11287 16779
rect 11713 16745 11747 16779
rect 11989 16745 12023 16779
rect 13001 16745 13035 16779
rect 14381 16745 14415 16779
rect 14565 16745 14599 16779
rect 14749 16745 14783 16779
rect 15209 16745 15243 16779
rect 9873 16677 9907 16711
rect 1409 16609 1443 16643
rect 1685 16609 1719 16643
rect 2145 16609 2179 16643
rect 10333 16609 10367 16643
rect 15117 16609 15151 16643
rect 15393 16609 15427 16643
rect 15669 16609 15703 16643
rect 1961 16541 1995 16575
rect 9965 16541 9999 16575
rect 1869 16473 1903 16507
rect 10609 16473 10643 16507
rect 15485 16473 15519 16507
rect 14933 16405 14967 16439
rect 14841 16201 14875 16235
rect 15301 16201 15335 16235
rect 15209 16133 15243 16167
rect 15025 15997 15059 16031
rect 15669 15997 15703 16031
rect 15485 15861 15519 15895
rect 15577 15657 15611 15691
rect 3893 15113 3927 15147
rect 4537 15113 4571 15147
rect 5365 15113 5399 15147
rect 7205 15045 7239 15079
rect 1409 14977 1443 15011
rect 4077 14909 4111 14943
rect 4721 14909 4755 14943
rect 5549 14909 5583 14943
rect 7389 14909 7423 14943
rect 1593 14841 1627 14875
rect 7481 14773 7515 14807
rect 9413 14569 9447 14603
rect 9597 14433 9631 14467
rect 15577 13481 15611 13515
rect 4690 13413 4724 13447
rect 2789 13345 2823 13379
rect 4445 13345 4479 13379
rect 15393 13345 15427 13379
rect 3065 13141 3099 13175
rect 3249 13141 3283 13175
rect 5825 13141 5859 13175
rect 15209 13141 15243 13175
rect 5365 12733 5399 12767
rect 5181 12597 5215 12631
rect 15485 12325 15519 12359
rect 15669 12325 15703 12359
rect 7297 12257 7331 12291
rect 7021 12189 7055 12223
rect 7205 12189 7239 12223
rect 7665 12053 7699 12087
rect 9965 11849 9999 11883
rect 1409 11645 1443 11679
rect 1685 11645 1719 11679
rect 8585 11645 8619 11679
rect 8493 11577 8527 11611
rect 8852 11577 8886 11611
rect 1593 11509 1627 11543
rect 7205 11509 7239 11543
rect 9137 11305 9171 11339
rect 7634 11237 7668 11271
rect 6929 11169 6963 11203
rect 7389 11169 7423 11203
rect 9321 11169 9355 11203
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 10057 11101 10091 11135
rect 7297 11033 7331 11067
rect 8769 10965 8803 10999
rect 7573 10761 7607 10795
rect 10977 10761 11011 10795
rect 3709 10625 3743 10659
rect 7021 10625 7055 10659
rect 7113 10625 7147 10659
rect 9045 10625 9079 10659
rect 9597 10625 9631 10659
rect 9689 10625 9723 10659
rect 10517 10625 10551 10659
rect 2948 10557 2982 10591
rect 10333 10557 10367 10591
rect 10425 10557 10459 10591
rect 3801 10489 3835 10523
rect 4721 10489 4755 10523
rect 7205 10489 7239 10523
rect 8789 10489 8823 10523
rect 3019 10421 3053 10455
rect 7665 10421 7699 10455
rect 9137 10421 9171 10455
rect 9505 10421 9539 10455
rect 9965 10421 9999 10455
rect 10793 10421 10827 10455
rect 6929 10217 6963 10251
rect 9965 10217 9999 10251
rect 1593 10149 1627 10183
rect 8524 10149 8558 10183
rect 8769 10081 8803 10115
rect 1501 10013 1535 10047
rect 1777 10013 1811 10047
rect 6745 10013 6779 10047
rect 6837 10013 6871 10047
rect 10057 10013 10091 10047
rect 10149 10013 10183 10047
rect 7297 9877 7331 9911
rect 7389 9877 7423 9911
rect 9597 9877 9631 9911
rect 7113 9673 7147 9707
rect 7573 9537 7607 9571
rect 7757 9537 7791 9571
rect 8861 9537 8895 9571
rect 7481 9469 7515 9503
rect 8769 9469 8803 9503
rect 8677 9401 8711 9435
rect 8309 9333 8343 9367
rect 7113 9129 7147 9163
rect 7021 9061 7055 9095
rect 12541 9061 12575 9095
rect 13277 8993 13311 9027
rect 7297 8925 7331 8959
rect 6653 8789 6687 8823
rect 13461 8789 13495 8823
rect 1593 8381 1627 8415
rect 1409 8313 1443 8347
rect 3525 7293 3559 7327
rect 3341 7157 3375 7191
rect 7021 5865 7055 5899
rect 9965 5865 9999 5899
rect 4077 5729 4111 5763
rect 6745 5729 6779 5763
rect 7205 5729 7239 5763
rect 7573 5729 7607 5763
rect 7849 5729 7883 5763
rect 9321 5729 9355 5763
rect 9689 5729 9723 5763
rect 9873 5729 9907 5763
rect 10149 5729 10183 5763
rect 10977 5729 11011 5763
rect 11805 5729 11839 5763
rect 7665 5593 7699 5627
rect 9505 5593 9539 5627
rect 9873 5593 9907 5627
rect 3893 5525 3927 5559
rect 6561 5525 6595 5559
rect 7389 5525 7423 5559
rect 9137 5525 9171 5559
rect 10793 5525 10827 5559
rect 11621 5525 11655 5559
rect 6653 5321 6687 5355
rect 8125 5321 8159 5355
rect 8493 5321 8527 5355
rect 8861 5321 8895 5355
rect 9137 5321 9171 5355
rect 9413 5321 9447 5355
rect 10057 5321 10091 5355
rect 10885 5321 10919 5355
rect 11713 5321 11747 5355
rect 12173 5321 12207 5355
rect 12633 5321 12667 5355
rect 12909 5321 12943 5355
rect 5825 5253 5859 5287
rect 7021 5253 7055 5287
rect 8585 5253 8619 5287
rect 10425 5253 10459 5287
rect 11161 5253 11195 5287
rect 1593 5117 1627 5151
rect 4629 5117 4663 5151
rect 4997 5117 5031 5151
rect 5365 5117 5399 5151
rect 5641 5117 5675 5151
rect 6009 5117 6043 5151
rect 6285 5117 6319 5151
rect 6837 5117 6871 5151
rect 7205 5117 7239 5151
rect 7665 5117 7699 5151
rect 7941 5117 7975 5151
rect 8309 5117 8343 5151
rect 8745 5117 8779 5151
rect 9045 5117 9079 5151
rect 9321 5117 9355 5151
rect 9505 5117 9539 5151
rect 9781 5117 9815 5151
rect 10241 5117 10275 5151
rect 10609 5117 10643 5151
rect 11069 5117 11103 5151
rect 11345 5117 11379 5151
rect 11897 5117 11931 5151
rect 12357 5117 12391 5151
rect 12817 5117 12851 5151
rect 13093 5117 13127 5151
rect 13369 5117 13403 5151
rect 1501 4981 1535 5015
rect 4445 4981 4479 5015
rect 4813 4981 4847 5015
rect 5181 4981 5215 5015
rect 5457 4981 5491 5015
rect 6101 4981 6135 5015
rect 7481 4981 7515 5015
rect 9597 4981 9631 5015
rect 13185 4981 13219 5015
rect 9505 4709 9539 4743
rect 9321 4641 9355 4675
rect 9137 4505 9171 4539
rect 15025 3689 15059 3723
rect 15485 3689 15519 3723
rect 15209 3553 15243 3587
rect 15669 3553 15703 3587
rect 15393 3349 15427 3383
rect 1409 3145 1443 3179
rect 15209 3145 15243 3179
rect 14105 3077 14139 3111
rect 14933 3009 14967 3043
rect 1593 2941 1627 2975
rect 15117 2941 15151 2975
rect 15393 2941 15427 2975
rect 15669 2941 15703 2975
rect 3801 2873 3835 2907
rect 4077 2873 4111 2907
rect 4261 2873 4295 2907
rect 14197 2873 14231 2907
rect 1685 2805 1719 2839
rect 3709 2805 3743 2839
rect 9873 2805 9907 2839
rect 11161 2805 11195 2839
rect 11805 2805 11839 2839
rect 12909 2805 12943 2839
rect 13829 2805 13863 2839
rect 14381 2805 14415 2839
rect 14749 2805 14783 2839
rect 15485 2805 15519 2839
rect 8769 2601 8803 2635
rect 9229 2601 9263 2635
rect 9597 2601 9631 2635
rect 10057 2601 10091 2635
rect 10885 2601 10919 2635
rect 11345 2601 11379 2635
rect 11897 2601 11931 2635
rect 13461 2601 13495 2635
rect 13921 2601 13955 2635
rect 14197 2601 14231 2635
rect 14565 2601 14599 2635
rect 14841 2601 14875 2635
rect 15117 2601 15151 2635
rect 2513 2533 2547 2567
rect 4077 2533 4111 2567
rect 4629 2533 4663 2567
rect 5549 2533 5583 2567
rect 6101 2533 6135 2567
rect 6285 2533 6319 2567
rect 7481 2533 7515 2567
rect 10333 2533 10367 2567
rect 11621 2533 11655 2567
rect 12449 2533 12483 2567
rect 15485 2533 15519 2567
rect 1593 2465 1627 2499
rect 1961 2465 1995 2499
rect 2329 2465 2363 2499
rect 2697 2465 2731 2499
rect 3065 2465 3099 2499
rect 3433 2465 3467 2499
rect 5089 2465 5123 2499
rect 5917 2465 5951 2499
rect 6745 2465 6779 2499
rect 7113 2465 7147 2499
rect 7849 2465 7883 2499
rect 8217 2465 8251 2499
rect 8585 2465 8619 2499
rect 8953 2465 8987 2499
rect 9413 2465 9447 2499
rect 9781 2465 9815 2499
rect 10241 2465 10275 2499
rect 10701 2465 10735 2499
rect 11069 2465 11103 2499
rect 11529 2465 11563 2499
rect 12081 2465 12115 2499
rect 12357 2465 12391 2499
rect 12817 2465 12851 2499
rect 13277 2465 13311 2499
rect 13645 2465 13679 2499
rect 14105 2465 14139 2499
rect 14381 2465 14415 2499
rect 14749 2465 14783 2499
rect 15025 2465 15059 2499
rect 15301 2465 15335 2499
rect 15669 2465 15703 2499
rect 2145 2397 2179 2431
rect 3893 2397 3927 2431
rect 6929 2397 6963 2431
rect 7297 2397 7331 2431
rect 9873 2397 9907 2431
rect 11161 2397 11195 2431
rect 12909 2397 12943 2431
rect 13737 2397 13771 2431
rect 1409 2329 1443 2363
rect 3249 2329 3283 2363
rect 4445 2329 4479 2363
rect 4905 2329 4939 2363
rect 5365 2329 5399 2363
rect 5733 2329 5767 2363
rect 6561 2329 6595 2363
rect 7665 2329 7699 2363
rect 8033 2329 8067 2363
rect 8401 2329 8435 2363
rect 12173 2329 12207 2363
rect 12633 2329 12667 2363
rect 1869 2261 1903 2295
rect 2973 2261 3007 2295
rect 10517 2261 10551 2295
rect 13093 2261 13127 2295
<< metal1 >>
rect 8294 17892 8300 17944
rect 8352 17932 8358 17944
rect 11974 17932 11980 17944
rect 8352 17904 11980 17932
rect 8352 17892 8358 17904
rect 11974 17892 11980 17904
rect 12032 17892 12038 17944
rect 6270 17824 6276 17876
rect 6328 17864 6334 17876
rect 10502 17864 10508 17876
rect 6328 17836 10508 17864
rect 6328 17824 6334 17836
rect 10502 17824 10508 17836
rect 10560 17824 10566 17876
rect 7834 17756 7840 17808
rect 7892 17796 7898 17808
rect 11790 17796 11796 17808
rect 7892 17768 11796 17796
rect 7892 17756 7898 17768
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 9214 17688 9220 17740
rect 9272 17728 9278 17740
rect 12250 17728 12256 17740
rect 9272 17700 12256 17728
rect 9272 17688 9278 17700
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 10318 17660 10324 17672
rect 7432 17632 10324 17660
rect 7432 17620 7438 17632
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 8202 17552 8208 17604
rect 8260 17592 8266 17604
rect 11422 17592 11428 17604
rect 8260 17564 11428 17592
rect 8260 17552 8266 17564
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 9306 17524 9312 17536
rect 4212 17496 9312 17524
rect 4212 17484 4218 17496
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 9490 17484 9496 17536
rect 9548 17524 9554 17536
rect 11606 17524 11612 17536
rect 9548 17496 11612 17524
rect 9548 17484 9554 17496
rect 11606 17484 11612 17496
rect 11664 17484 11670 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 16114 17524 16120 17536
rect 15620 17496 16120 17524
rect 15620 17484 15626 17496
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 1104 17434 16008 17456
rect 1104 17382 3480 17434
rect 3532 17382 3544 17434
rect 3596 17382 3608 17434
rect 3660 17382 3672 17434
rect 3724 17382 8478 17434
rect 8530 17382 8542 17434
rect 8594 17382 8606 17434
rect 8658 17382 8670 17434
rect 8722 17382 13475 17434
rect 13527 17382 13539 17434
rect 13591 17382 13603 17434
rect 13655 17382 13667 17434
rect 13719 17382 16008 17434
rect 1104 17360 16008 17382
rect 1026 17280 1032 17332
rect 1084 17320 1090 17332
rect 1857 17323 1915 17329
rect 1857 17320 1869 17323
rect 1084 17292 1869 17320
rect 1084 17280 1090 17292
rect 1857 17289 1869 17292
rect 1903 17289 1915 17323
rect 1857 17283 1915 17289
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2961 17323 3019 17329
rect 2961 17320 2973 17323
rect 2280 17292 2973 17320
rect 2280 17280 2286 17292
rect 2961 17289 2973 17292
rect 3007 17289 3019 17323
rect 2961 17283 3019 17289
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3973 17323 4031 17329
rect 3973 17320 3985 17323
rect 3108 17292 3985 17320
rect 3108 17280 3114 17292
rect 3973 17289 3985 17292
rect 4019 17289 4031 17323
rect 3973 17283 4031 17289
rect 4338 17280 4344 17332
rect 4396 17320 4402 17332
rect 8481 17323 8539 17329
rect 8481 17320 8493 17323
rect 4396 17292 8493 17320
rect 4396 17280 4402 17292
rect 8481 17289 8493 17292
rect 8527 17289 8539 17323
rect 8481 17283 8539 17289
rect 8665 17323 8723 17329
rect 8665 17289 8677 17323
rect 8711 17320 8723 17323
rect 8846 17320 8852 17332
rect 8711 17292 8852 17320
rect 8711 17289 8723 17292
rect 8665 17283 8723 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 9364 17292 9409 17320
rect 9364 17280 9370 17292
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 11333 17323 11391 17329
rect 11333 17320 11345 17323
rect 9640 17292 11345 17320
rect 9640 17280 9646 17292
rect 11333 17289 11345 17292
rect 11379 17289 11391 17323
rect 11333 17283 11391 17289
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 12713 17323 12771 17329
rect 12713 17320 12725 17323
rect 11664 17292 12725 17320
rect 11664 17280 11670 17292
rect 12713 17289 12725 17292
rect 12759 17289 12771 17323
rect 12713 17283 12771 17289
rect 566 17212 572 17264
rect 624 17252 630 17264
rect 1397 17255 1455 17261
rect 1397 17252 1409 17255
rect 624 17224 1409 17252
rect 624 17212 630 17224
rect 1397 17221 1409 17224
rect 1443 17221 1455 17255
rect 1397 17215 1455 17221
rect 2774 17212 2780 17264
rect 2832 17252 2838 17264
rect 3237 17255 3295 17261
rect 3237 17252 3249 17255
rect 2832 17224 3249 17252
rect 2832 17212 2838 17224
rect 3237 17221 3249 17224
rect 3283 17221 3295 17255
rect 3237 17215 3295 17221
rect 3786 17212 3792 17264
rect 3844 17252 3850 17264
rect 4249 17255 4307 17261
rect 4249 17252 4261 17255
rect 3844 17224 4261 17252
rect 3844 17212 3850 17224
rect 4249 17221 4261 17224
rect 4295 17221 4307 17255
rect 4798 17252 4804 17264
rect 4759 17224 4804 17252
rect 4249 17215 4307 17221
rect 4798 17212 4804 17224
rect 4856 17212 4862 17264
rect 5166 17252 5172 17264
rect 5127 17224 5172 17252
rect 5166 17212 5172 17224
rect 5224 17212 5230 17264
rect 5626 17252 5632 17264
rect 5587 17224 5632 17252
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 5994 17252 6000 17264
rect 5955 17224 6000 17252
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 6454 17212 6460 17264
rect 6512 17252 6518 17264
rect 6549 17255 6607 17261
rect 6549 17252 6561 17255
rect 6512 17224 6561 17252
rect 6512 17212 6518 17224
rect 6549 17221 6561 17224
rect 6595 17221 6607 17255
rect 6549 17215 6607 17221
rect 6914 17212 6920 17264
rect 6972 17252 6978 17264
rect 7282 17252 7288 17264
rect 6972 17224 7017 17252
rect 7243 17224 7288 17252
rect 6972 17212 6978 17224
rect 7282 17212 7288 17224
rect 7340 17212 7346 17264
rect 7742 17252 7748 17264
rect 7703 17224 7748 17252
rect 7742 17212 7748 17224
rect 7800 17212 7806 17264
rect 8110 17252 8116 17264
rect 8071 17224 8116 17252
rect 8110 17212 8116 17224
rect 8168 17212 8174 17264
rect 10229 17255 10287 17261
rect 10229 17252 10241 17255
rect 8404 17224 10241 17252
rect 1854 17144 1860 17196
rect 1912 17184 1918 17196
rect 2501 17187 2559 17193
rect 2501 17184 2513 17187
rect 1912 17156 2513 17184
rect 1912 17144 1918 17156
rect 2501 17153 2513 17156
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 5074 17144 5080 17196
rect 5132 17184 5138 17196
rect 8404 17184 8432 17224
rect 10229 17221 10241 17224
rect 10275 17221 10287 17255
rect 10229 17215 10287 17221
rect 10318 17212 10324 17264
rect 10376 17252 10382 17264
rect 10505 17255 10563 17261
rect 10505 17252 10517 17255
rect 10376 17224 10517 17252
rect 10376 17212 10382 17224
rect 10505 17221 10517 17224
rect 10551 17221 10563 17255
rect 10505 17215 10563 17221
rect 10594 17212 10600 17264
rect 10652 17252 10658 17264
rect 13173 17255 13231 17261
rect 13173 17252 13185 17255
rect 10652 17224 13185 17252
rect 10652 17212 10658 17224
rect 13173 17221 13185 17224
rect 13219 17221 13231 17255
rect 15654 17252 15660 17264
rect 15615 17224 15660 17252
rect 13173 17215 13231 17221
rect 15654 17212 15660 17224
rect 15712 17212 15718 17264
rect 5132 17156 8432 17184
rect 8481 17187 8539 17193
rect 5132 17144 5138 17156
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 8527 17156 9597 17184
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 9585 17153 9597 17156
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 9824 17156 10732 17184
rect 9824 17144 9830 17156
rect 1394 17076 1400 17128
rect 1452 17116 1458 17128
rect 2133 17119 2191 17125
rect 2133 17116 2145 17119
rect 1452 17088 2145 17116
rect 1452 17076 1458 17088
rect 2133 17085 2145 17088
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17116 2375 17119
rect 4522 17116 4528 17128
rect 2363 17088 4528 17116
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 4522 17076 4528 17088
rect 4580 17076 4586 17128
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 8662 17116 8668 17128
rect 7147 17088 8668 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 8757 17119 8815 17125
rect 8757 17085 8769 17119
rect 8803 17116 8815 17119
rect 9674 17116 9680 17128
rect 8803 17088 9680 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 10134 17116 10140 17128
rect 10095 17088 10140 17116
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 10410 17116 10416 17128
rect 10371 17088 10416 17116
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 10704 17125 10732 17156
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11330 17184 11336 17196
rect 11112 17156 11336 17184
rect 11112 17144 11118 17156
rect 11330 17144 11336 17156
rect 11388 17184 11394 17196
rect 11388 17156 11560 17184
rect 11388 17144 11394 17156
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 1578 17048 1584 17060
rect 1539 17020 1584 17048
rect 1578 17008 1584 17020
rect 1636 17008 1642 17060
rect 1946 17048 1952 17060
rect 1907 17020 1952 17048
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 2682 17048 2688 17060
rect 2643 17020 2688 17048
rect 2682 17008 2688 17020
rect 2740 17008 2746 17060
rect 3053 17051 3111 17057
rect 3053 17017 3065 17051
rect 3099 17017 3111 17051
rect 3053 17011 3111 17017
rect 3068 16980 3096 17011
rect 3234 17008 3240 17060
rect 3292 17048 3298 17060
rect 3421 17051 3479 17057
rect 3421 17048 3433 17051
rect 3292 17020 3433 17048
rect 3292 17008 3298 17020
rect 3421 17017 3433 17020
rect 3467 17017 3479 17051
rect 4062 17048 4068 17060
rect 4023 17020 4068 17048
rect 3421 17011 3479 17017
rect 4062 17008 4068 17020
rect 4120 17008 4126 17060
rect 4430 17048 4436 17060
rect 4391 17020 4436 17048
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 4982 17048 4988 17060
rect 4943 17020 4988 17048
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 5350 17048 5356 17060
rect 5311 17020 5356 17048
rect 5350 17008 5356 17020
rect 5408 17008 5414 17060
rect 5810 17048 5816 17060
rect 5771 17020 5816 17048
rect 5810 17008 5816 17020
rect 5868 17008 5874 17060
rect 6181 17051 6239 17057
rect 6181 17017 6193 17051
rect 6227 17048 6239 17051
rect 6546 17048 6552 17060
rect 6227 17020 6552 17048
rect 6227 17017 6239 17020
rect 6181 17011 6239 17017
rect 6546 17008 6552 17020
rect 6604 17008 6610 17060
rect 6730 17048 6736 17060
rect 6691 17020 6736 17048
rect 6730 17008 6736 17020
rect 6788 17008 6794 17060
rect 7466 17048 7472 17060
rect 7427 17020 7472 17048
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 7929 17051 7987 17057
rect 7929 17017 7941 17051
rect 7975 17048 7987 17051
rect 8110 17048 8116 17060
rect 7975 17020 8116 17048
rect 7975 17017 7987 17020
rect 7929 17011 7987 17017
rect 8110 17008 8116 17020
rect 8168 17008 8174 17060
rect 8294 17048 8300 17060
rect 8255 17020 8300 17048
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 9401 17051 9459 17057
rect 9401 17048 9413 17051
rect 8772 17020 9413 17048
rect 5258 16980 5264 16992
rect 3068 16952 5264 16980
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 8018 16940 8024 16992
rect 8076 16980 8082 16992
rect 8772 16980 8800 17020
rect 9401 17017 9413 17020
rect 9447 17017 9459 17051
rect 9401 17011 9459 17017
rect 9769 17051 9827 17057
rect 9769 17017 9781 17051
rect 9815 17048 9827 17051
rect 10042 17048 10048 17060
rect 9815 17020 10048 17048
rect 9815 17017 9827 17020
rect 9769 17011 9827 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10226 17008 10232 17060
rect 10284 17048 10290 17060
rect 10980 17048 11008 17079
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11532 17125 11560 17156
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 11940 17156 12388 17184
rect 11940 17144 11946 17156
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 11204 17088 11253 17116
rect 11204 17076 11210 17088
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 11241 17079 11299 17085
rect 11517 17119 11575 17125
rect 11517 17085 11529 17119
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 10284 17020 11008 17048
rect 11256 17048 11284 17079
rect 11606 17076 11612 17128
rect 11664 17116 11670 17128
rect 12360 17125 12388 17156
rect 12636 17156 13001 17184
rect 12069 17119 12127 17125
rect 12069 17116 12081 17119
rect 11664 17088 12081 17116
rect 11664 17076 11670 17088
rect 12069 17085 12081 17088
rect 12115 17085 12127 17119
rect 12069 17079 12127 17085
rect 12345 17119 12403 17125
rect 12345 17085 12357 17119
rect 12391 17085 12403 17119
rect 12345 17079 12403 17085
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12636 17125 12664 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 13817 17187 13875 17193
rect 13817 17184 13829 17187
rect 12989 17147 13047 17153
rect 13372 17156 13829 17184
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12492 17088 12633 17116
rect 12492 17076 12498 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12768 17088 12909 17116
rect 12768 17076 12774 17088
rect 12897 17085 12909 17088
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13372 17125 13400 17156
rect 13817 17153 13829 17156
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 13357 17119 13415 17125
rect 13357 17116 13369 17119
rect 13228 17088 13369 17116
rect 13228 17076 13234 17088
rect 13357 17085 13369 17088
rect 13403 17085 13415 17119
rect 13357 17079 13415 17085
rect 13446 17076 13452 17128
rect 13504 17116 13510 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13504 17088 13737 17116
rect 13504 17076 13510 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 11701 17051 11759 17057
rect 11701 17048 11713 17051
rect 11256 17020 11713 17048
rect 10284 17008 10290 17020
rect 11701 17017 11713 17020
rect 11747 17017 11759 17051
rect 13740 17048 13768 17079
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 14185 17119 14243 17125
rect 14185 17116 14197 17119
rect 14056 17088 14197 17116
rect 14056 17076 14062 17088
rect 14185 17085 14197 17088
rect 14231 17116 14243 17119
rect 14366 17116 14372 17128
rect 14231 17088 14372 17116
rect 14231 17085 14243 17088
rect 14185 17079 14243 17085
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14516 17088 14749 17116
rect 14516 17076 14522 17088
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 14826 17076 14832 17128
rect 14884 17116 14890 17128
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 14884 17088 15025 17116
rect 14884 17076 14890 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15286 17116 15292 17128
rect 15247 17088 15292 17116
rect 15013 17079 15071 17085
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 14277 17051 14335 17057
rect 14277 17048 14289 17051
rect 13740 17020 14289 17048
rect 11701 17011 11759 17017
rect 14277 17017 14289 17020
rect 14323 17017 14335 17051
rect 15470 17048 15476 17060
rect 15431 17020 15476 17048
rect 14277 17011 14335 17017
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 8076 16952 8800 16980
rect 8076 16940 8082 16952
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 8904 16952 9965 16980
rect 8904 16940 8910 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10560 16952 10793 16980
rect 10560 16940 10566 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 11057 16983 11115 16989
rect 11057 16949 11069 16983
rect 11103 16980 11115 16983
rect 11422 16980 11428 16992
rect 11103 16952 11428 16980
rect 11103 16949 11115 16952
rect 11057 16943 11115 16949
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 11848 16952 11897 16980
rect 11848 16940 11854 16952
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 12158 16980 12164 16992
rect 12119 16952 12164 16980
rect 11885 16943 11943 16949
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12250 16940 12256 16992
rect 12308 16980 12314 16992
rect 12437 16983 12495 16989
rect 12437 16980 12449 16983
rect 12308 16952 12449 16980
rect 12308 16940 12314 16952
rect 12437 16949 12449 16952
rect 12483 16949 12495 16983
rect 12437 16943 12495 16949
rect 13354 16940 13360 16992
rect 13412 16980 13418 16992
rect 13541 16983 13599 16989
rect 13541 16980 13553 16983
rect 13412 16952 13553 16980
rect 13412 16940 13418 16952
rect 13541 16949 13553 16952
rect 13587 16949 13599 16983
rect 13998 16980 14004 16992
rect 13959 16952 14004 16980
rect 13541 16943 13599 16949
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14550 16980 14556 16992
rect 14511 16952 14556 16980
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 14826 16980 14832 16992
rect 14787 16952 14832 16980
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 15102 16980 15108 16992
rect 15063 16952 15108 16980
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 1104 16890 16008 16912
rect 1104 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 10976 16890
rect 11028 16838 11040 16890
rect 11092 16838 11104 16890
rect 11156 16838 11168 16890
rect 11220 16838 16008 16890
rect 1104 16816 16008 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 2774 16776 2780 16788
rect 1627 16748 2780 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 9582 16776 9588 16788
rect 6696 16748 9588 16776
rect 6696 16736 6702 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9953 16779 10011 16785
rect 9953 16776 9965 16779
rect 9692 16748 9965 16776
rect 3970 16708 3976 16720
rect 2240 16680 3976 16708
rect 198 16600 204 16652
rect 256 16640 262 16652
rect 1397 16643 1455 16649
rect 1397 16640 1409 16643
rect 256 16612 1409 16640
rect 256 16600 262 16612
rect 1397 16609 1409 16612
rect 1443 16640 1455 16643
rect 1670 16640 1676 16652
rect 1443 16612 1532 16640
rect 1631 16612 1676 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1504 16572 1532 16612
rect 1670 16600 1676 16612
rect 1728 16640 1734 16652
rect 2133 16643 2191 16649
rect 2133 16640 2145 16643
rect 1728 16612 2145 16640
rect 1728 16600 1734 16612
rect 2133 16609 2145 16612
rect 2179 16609 2191 16643
rect 2133 16603 2191 16609
rect 1949 16575 2007 16581
rect 1949 16572 1961 16575
rect 1504 16544 1961 16572
rect 1949 16541 1961 16544
rect 1995 16541 2007 16575
rect 2240 16572 2268 16680
rect 3970 16668 3976 16680
rect 4028 16668 4034 16720
rect 7742 16668 7748 16720
rect 7800 16708 7806 16720
rect 8846 16708 8852 16720
rect 7800 16680 8852 16708
rect 7800 16668 7806 16680
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 9692 16640 9720 16748
rect 9953 16745 9965 16748
rect 9999 16745 10011 16779
rect 9953 16739 10011 16745
rect 10045 16779 10103 16785
rect 10045 16745 10057 16779
rect 10091 16776 10103 16779
rect 10410 16776 10416 16788
rect 10091 16748 10416 16776
rect 10091 16745 10103 16748
rect 10045 16739 10103 16745
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16776 11299 16779
rect 11330 16776 11336 16788
rect 11287 16748 11336 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 11701 16779 11759 16785
rect 11701 16776 11713 16779
rect 11572 16748 11713 16776
rect 11572 16736 11578 16748
rect 11701 16745 11713 16748
rect 11747 16745 11759 16779
rect 11701 16739 11759 16745
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 11977 16779 12035 16785
rect 11977 16776 11989 16779
rect 11940 16748 11989 16776
rect 11940 16736 11946 16748
rect 11977 16745 11989 16748
rect 12023 16745 12035 16779
rect 11977 16739 12035 16745
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 12989 16779 13047 16785
rect 12989 16776 13001 16779
rect 12768 16748 13001 16776
rect 12768 16736 12774 16748
rect 12989 16745 13001 16748
rect 13035 16745 13047 16779
rect 14366 16776 14372 16788
rect 14327 16748 14372 16776
rect 12989 16739 13047 16745
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 14553 16779 14611 16785
rect 14553 16776 14565 16779
rect 14516 16748 14565 16776
rect 14516 16736 14522 16748
rect 14553 16745 14565 16748
rect 14599 16745 14611 16779
rect 14734 16776 14740 16788
rect 14695 16748 14740 16776
rect 14553 16739 14611 16745
rect 14734 16736 14740 16748
rect 14792 16736 14798 16788
rect 15197 16779 15255 16785
rect 15197 16745 15209 16779
rect 15243 16745 15255 16779
rect 15197 16739 15255 16745
rect 9861 16711 9919 16717
rect 9861 16677 9873 16711
rect 9907 16708 9919 16711
rect 10134 16708 10140 16720
rect 9907 16680 10140 16708
rect 9907 16677 9919 16680
rect 9861 16671 9919 16677
rect 10134 16668 10140 16680
rect 10192 16668 10198 16720
rect 11606 16708 11612 16720
rect 10520 16680 11612 16708
rect 8168 16612 9720 16640
rect 8168 16600 8174 16612
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10321 16643 10379 16649
rect 10321 16640 10333 16643
rect 9824 16612 10333 16640
rect 9824 16600 9830 16612
rect 10321 16609 10333 16612
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 1949 16535 2007 16541
rect 2056 16544 2268 16572
rect 9953 16575 10011 16581
rect 1857 16507 1915 16513
rect 1857 16473 1869 16507
rect 1903 16504 1915 16507
rect 2056 16504 2084 16544
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10520 16572 10548 16680
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 11790 16668 11796 16720
rect 11848 16708 11854 16720
rect 15212 16708 15240 16739
rect 11848 16680 15240 16708
rect 11848 16668 11854 16680
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 12158 16640 12164 16652
rect 10836 16612 12164 16640
rect 10836 16600 10842 16612
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 15105 16643 15163 16649
rect 13280 16612 14964 16640
rect 9999 16544 10548 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 13280 16572 13308 16612
rect 10928 16544 13308 16572
rect 10928 16532 10934 16544
rect 1903 16476 2084 16504
rect 1903 16473 1915 16476
rect 1857 16467 1915 16473
rect 8938 16464 8944 16516
rect 8996 16504 9002 16516
rect 10134 16504 10140 16516
rect 8996 16476 10140 16504
rect 8996 16464 9002 16476
rect 10134 16464 10140 16476
rect 10192 16464 10198 16516
rect 10226 16464 10232 16516
rect 10284 16504 10290 16516
rect 10597 16507 10655 16513
rect 10597 16504 10609 16507
rect 10284 16476 10609 16504
rect 10284 16464 10290 16476
rect 10597 16473 10609 16476
rect 10643 16473 10655 16507
rect 14936 16504 14964 16612
rect 15105 16609 15117 16643
rect 15151 16609 15163 16643
rect 15105 16603 15163 16609
rect 15381 16643 15439 16649
rect 15381 16609 15393 16643
rect 15427 16640 15439 16643
rect 15562 16640 15568 16652
rect 15427 16612 15568 16640
rect 15427 16609 15439 16612
rect 15381 16603 15439 16609
rect 15010 16532 15016 16584
rect 15068 16572 15074 16584
rect 15120 16572 15148 16603
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 15746 16640 15752 16652
rect 15703 16612 15752 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 16942 16572 16948 16584
rect 15068 16544 16948 16572
rect 15068 16532 15074 16544
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 15473 16507 15531 16513
rect 15473 16504 15485 16507
rect 14936 16476 15485 16504
rect 10597 16467 10655 16473
rect 15473 16473 15485 16476
rect 15519 16473 15531 16507
rect 15473 16467 15531 16473
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 10410 16436 10416 16448
rect 9456 16408 10416 16436
rect 9456 16396 9462 16408
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 14918 16436 14924 16448
rect 14879 16408 14924 16436
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 1104 16346 16008 16368
rect 1104 16294 3480 16346
rect 3532 16294 3544 16346
rect 3596 16294 3608 16346
rect 3660 16294 3672 16346
rect 3724 16294 8478 16346
rect 8530 16294 8542 16346
rect 8594 16294 8606 16346
rect 8658 16294 8670 16346
rect 8722 16294 13475 16346
rect 13527 16294 13539 16346
rect 13591 16294 13603 16346
rect 13655 16294 13667 16346
rect 13719 16294 16008 16346
rect 1104 16272 16008 16294
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 12618 16232 12624 16244
rect 9732 16204 12624 16232
rect 9732 16192 9738 16204
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 15010 16232 15016 16244
rect 14875 16204 15016 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 15197 16167 15255 16173
rect 15197 16133 15209 16167
rect 15243 16164 15255 16167
rect 15746 16164 15752 16176
rect 15243 16136 15752 16164
rect 15243 16133 15255 16136
rect 15197 16127 15255 16133
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 16028 15071 16031
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 15059 16000 15669 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 15657 15997 15669 16000
rect 15703 16028 15715 16031
rect 16482 16028 16488 16040
rect 15703 16000 16488 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 15473 15895 15531 15901
rect 15473 15892 15485 15895
rect 13136 15864 15485 15892
rect 13136 15852 13142 15864
rect 15473 15861 15485 15864
rect 15519 15861 15531 15895
rect 15473 15855 15531 15861
rect 1104 15802 16008 15824
rect 1104 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 10976 15802
rect 11028 15750 11040 15802
rect 11092 15750 11104 15802
rect 11156 15750 11168 15802
rect 11220 15750 16008 15802
rect 1104 15728 16008 15750
rect 15562 15688 15568 15700
rect 15523 15660 15568 15688
rect 15562 15648 15568 15660
rect 15620 15648 15626 15700
rect 1104 15258 16008 15280
rect 1104 15206 3480 15258
rect 3532 15206 3544 15258
rect 3596 15206 3608 15258
rect 3660 15206 3672 15258
rect 3724 15206 8478 15258
rect 8530 15206 8542 15258
rect 8594 15206 8606 15258
rect 8658 15206 8670 15258
rect 8722 15206 13475 15258
rect 13527 15206 13539 15258
rect 13591 15206 13603 15258
rect 13655 15206 13667 15258
rect 13719 15206 16008 15258
rect 1104 15184 16008 15206
rect 1578 15104 1584 15156
rect 1636 15144 1642 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 1636 15116 3893 15144
rect 1636 15104 1642 15116
rect 3881 15113 3893 15116
rect 3927 15113 3939 15147
rect 4522 15144 4528 15156
rect 4483 15116 4528 15144
rect 3881 15107 3939 15113
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 5258 15104 5264 15156
rect 5316 15144 5322 15156
rect 5353 15147 5411 15153
rect 5353 15144 5365 15147
rect 5316 15116 5365 15144
rect 5316 15104 5322 15116
rect 5353 15113 5365 15116
rect 5399 15113 5411 15147
rect 5353 15107 5411 15113
rect 4982 15036 4988 15088
rect 5040 15076 5046 15088
rect 7193 15079 7251 15085
rect 7193 15076 7205 15079
rect 5040 15048 7205 15076
rect 5040 15036 5046 15048
rect 7193 15045 7205 15048
rect 7239 15045 7251 15079
rect 7193 15039 7251 15045
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 4065 14943 4123 14949
rect 4065 14909 4077 14943
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14909 4767 14943
rect 4709 14903 4767 14909
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14940 5595 14943
rect 7377 14943 7435 14949
rect 5583 14912 7236 14940
rect 5583 14909 5595 14912
rect 5537 14903 5595 14909
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14872 1639 14875
rect 1762 14872 1768 14884
rect 1627 14844 1768 14872
rect 1627 14841 1639 14844
rect 1581 14835 1639 14841
rect 1762 14832 1768 14844
rect 1820 14832 1826 14884
rect 4080 14804 4108 14903
rect 4724 14872 4752 14903
rect 7098 14872 7104 14884
rect 4724 14844 7104 14872
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7208 14872 7236 14912
rect 7377 14909 7389 14943
rect 7423 14940 7435 14943
rect 7423 14912 7696 14940
rect 7423 14909 7435 14912
rect 7377 14903 7435 14909
rect 7558 14872 7564 14884
rect 7208 14844 7564 14872
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 7282 14804 7288 14816
rect 4080 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 7668 14804 7696 14912
rect 9398 14804 9404 14816
rect 7515 14776 9404 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 1104 14714 16008 14736
rect 1104 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 10976 14714
rect 11028 14662 11040 14714
rect 11092 14662 11104 14714
rect 11156 14662 11168 14714
rect 11220 14662 16008 14714
rect 1104 14640 16008 14662
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 7524 14572 9413 14600
rect 7524 14560 7530 14572
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 9950 14464 9956 14476
rect 9631 14436 9956 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 1104 14170 16008 14192
rect 1104 14118 3480 14170
rect 3532 14118 3544 14170
rect 3596 14118 3608 14170
rect 3660 14118 3672 14170
rect 3724 14118 8478 14170
rect 8530 14118 8542 14170
rect 8594 14118 8606 14170
rect 8658 14118 8670 14170
rect 8722 14118 13475 14170
rect 13527 14118 13539 14170
rect 13591 14118 13603 14170
rect 13655 14118 13667 14170
rect 13719 14118 16008 14170
rect 1104 14096 16008 14118
rect 1104 13626 16008 13648
rect 1104 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 10976 13626
rect 11028 13574 11040 13626
rect 11092 13574 11104 13626
rect 11156 13574 11168 13626
rect 11220 13574 16008 13626
rect 1104 13552 16008 13574
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15565 13515 15623 13521
rect 15565 13512 15577 13515
rect 15528 13484 15577 13512
rect 15528 13472 15534 13484
rect 15565 13481 15577 13484
rect 15611 13481 15623 13515
rect 15565 13475 15623 13481
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 4678 13447 4736 13453
rect 4678 13444 4690 13447
rect 4028 13416 4690 13444
rect 4028 13404 4034 13416
rect 4678 13413 4690 13416
rect 4724 13413 4736 13447
rect 4678 13407 4736 13413
rect 2774 13376 2780 13388
rect 2735 13348 2780 13376
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 5534 13376 5540 13388
rect 4479 13348 5540 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15381 13379 15439 13385
rect 15381 13376 15393 13379
rect 15252 13348 15393 13376
rect 15252 13336 15258 13348
rect 15381 13345 15393 13348
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 9582 13240 9588 13252
rect 3068 13212 3372 13240
rect 3068 13181 3096 13212
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13141 3111 13175
rect 3053 13135 3111 13141
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 3237 13175 3295 13181
rect 3237 13172 3249 13175
rect 3200 13144 3249 13172
rect 3200 13132 3206 13144
rect 3237 13141 3249 13144
rect 3283 13141 3295 13175
rect 3344 13172 3372 13212
rect 5368 13212 9588 13240
rect 5368 13172 5396 13212
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 3344 13144 5396 13172
rect 5813 13175 5871 13181
rect 3237 13135 3295 13141
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 7006 13172 7012 13184
rect 5859 13144 7012 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 15194 13172 15200 13184
rect 15155 13144 15200 13172
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 1104 13082 16008 13104
rect 1104 13030 3480 13082
rect 3532 13030 3544 13082
rect 3596 13030 3608 13082
rect 3660 13030 3672 13082
rect 3724 13030 8478 13082
rect 8530 13030 8542 13082
rect 8594 13030 8606 13082
rect 8658 13030 8670 13082
rect 8722 13030 13475 13082
rect 13527 13030 13539 13082
rect 13591 13030 13603 13082
rect 13655 13030 13667 13082
rect 13719 13030 16008 13082
rect 1104 13008 16008 13030
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12764 5411 12767
rect 6362 12764 6368 12776
rect 5399 12736 6368 12764
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5534 12628 5540 12640
rect 5215 12600 5540 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 1104 12538 16008 12560
rect 1104 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 10976 12538
rect 11028 12486 11040 12538
rect 11092 12486 11104 12538
rect 11156 12486 11168 12538
rect 11220 12486 16008 12538
rect 1104 12464 16008 12486
rect 9582 12316 9588 12368
rect 9640 12356 9646 12368
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 9640 12328 15485 12356
rect 9640 12316 9646 12328
rect 15473 12325 15485 12328
rect 15519 12325 15531 12359
rect 15654 12356 15660 12368
rect 15615 12328 15660 12356
rect 15473 12319 15531 12325
rect 15654 12316 15660 12328
rect 15712 12316 15718 12368
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 6972 12260 7297 12288
rect 6972 12248 6978 12260
rect 7285 12257 7297 12260
rect 7331 12288 7343 12291
rect 7374 12288 7380 12300
rect 7331 12260 7380 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7006 12220 7012 12232
rect 6967 12192 7012 12220
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7190 12220 7196 12232
rect 7151 12192 7196 12220
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 7524 12056 7665 12084
rect 7524 12044 7530 12056
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 7653 12047 7711 12053
rect 1104 11994 16008 12016
rect 1104 11942 3480 11994
rect 3532 11942 3544 11994
rect 3596 11942 3608 11994
rect 3660 11942 3672 11994
rect 3724 11942 8478 11994
rect 8530 11942 8542 11994
rect 8594 11942 8606 11994
rect 8658 11942 8670 11994
rect 8722 11942 13475 11994
rect 13527 11942 13539 11994
rect 13591 11942 13603 11994
rect 13655 11942 13667 11994
rect 13719 11942 16008 11994
rect 1104 11920 16008 11942
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9640 11852 9965 11880
rect 9640 11840 9646 11852
rect 9953 11849 9965 11852
rect 9999 11849 10011 11883
rect 9953 11843 10011 11849
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11676 1458 11688
rect 1673 11679 1731 11685
rect 1673 11676 1685 11679
rect 1452 11648 1685 11676
rect 1452 11636 1458 11648
rect 1673 11645 1685 11648
rect 1719 11645 1731 11679
rect 8570 11676 8576 11688
rect 8531 11648 8576 11676
rect 1673 11639 1731 11645
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 12526 11676 12532 11688
rect 8772 11648 12532 11676
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 7742 11608 7748 11620
rect 7156 11580 7748 11608
rect 7156 11568 7162 11580
rect 7742 11568 7748 11580
rect 7800 11568 7806 11620
rect 8481 11611 8539 11617
rect 8481 11577 8493 11611
rect 8527 11608 8539 11611
rect 8772 11608 8800 11648
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 8527 11580 8800 11608
rect 8840 11611 8898 11617
rect 8527 11577 8539 11580
rect 8481 11571 8539 11577
rect 8840 11577 8852 11611
rect 8886 11608 8898 11611
rect 9306 11608 9312 11620
rect 8886 11580 9312 11608
rect 8886 11577 8898 11580
rect 8840 11571 8898 11577
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 3234 11540 3240 11552
rect 1627 11512 3240 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 6420 11512 7205 11540
rect 6420 11500 6426 11512
rect 7193 11509 7205 11512
rect 7239 11540 7251 11543
rect 8110 11540 8116 11552
rect 7239 11512 8116 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 1104 11450 16008 11472
rect 1104 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 10976 11450
rect 11028 11398 11040 11450
rect 11092 11398 11104 11450
rect 11156 11398 11168 11450
rect 11220 11398 16008 11450
rect 1104 11376 16008 11398
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5592 11308 7420 11336
rect 5592 11296 5598 11308
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7098 11200 7104 11212
rect 6963 11172 7104 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7282 11160 7288 11212
rect 7340 11160 7346 11212
rect 7392 11209 7420 11308
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 9030 11336 9036 11348
rect 8628 11308 9036 11336
rect 8628 11296 8634 11308
rect 9030 11296 9036 11308
rect 9088 11336 9094 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 9088 11308 9137 11336
rect 9088 11296 9094 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9125 11299 9183 11305
rect 7558 11228 7564 11280
rect 7616 11277 7622 11280
rect 7616 11271 7680 11277
rect 7616 11237 7634 11271
rect 7668 11237 7680 11271
rect 7616 11231 7680 11237
rect 7616 11228 7622 11231
rect 7742 11228 7748 11280
rect 7800 11228 7806 11280
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11169 7435 11203
rect 7760 11200 7788 11228
rect 7377 11163 7435 11169
rect 7484 11172 7788 11200
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 7300 11132 7328 11160
rect 7484 11132 7512 11172
rect 8110 11160 8116 11212
rect 8168 11200 8174 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 8168 11172 9321 11200
rect 8168 11160 8174 11172
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9309 11163 9367 11169
rect 10042 11132 10048 11144
rect 6871 11104 7512 11132
rect 10003 11104 10048 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 6748 11064 6776 11095
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 7006 11064 7012 11076
rect 6748 11036 7012 11064
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7282 11064 7288 11076
rect 7243 11036 7288 11064
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7024 10996 7052 11024
rect 7558 10996 7564 11008
rect 7024 10968 7564 10996
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8757 10999 8815 11005
rect 8757 10996 8769 10999
rect 8352 10968 8769 10996
rect 8352 10956 8358 10968
rect 8757 10965 8769 10968
rect 8803 10965 8815 10999
rect 8757 10959 8815 10965
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 15194 10996 15200 11008
rect 8996 10968 15200 10996
rect 8996 10956 9002 10968
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 1104 10906 16008 10928
rect 1104 10854 3480 10906
rect 3532 10854 3544 10906
rect 3596 10854 3608 10906
rect 3660 10854 3672 10906
rect 3724 10854 8478 10906
rect 8530 10854 8542 10906
rect 8594 10854 8606 10906
rect 8658 10854 8670 10906
rect 8722 10854 13475 10906
rect 13527 10854 13539 10906
rect 13591 10854 13603 10906
rect 13655 10854 13667 10906
rect 13719 10854 16008 10906
rect 1104 10832 16008 10854
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 7607 10764 9628 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3292 10628 3709 10656
rect 3292 10616 3298 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 7006 10656 7012 10668
rect 6967 10628 7012 10656
rect 3697 10619 3755 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7650 10656 7656 10668
rect 7147 10628 7656 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 9600 10665 9628 10764
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10928 10764 10977 10792
rect 10928 10752 10934 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10656 9735 10659
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 9723 10628 10517 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 2936 10591 2994 10597
rect 2936 10557 2948 10591
rect 2982 10588 2994 10591
rect 3142 10588 3148 10600
rect 2982 10560 3148 10588
rect 2982 10557 2994 10560
rect 2936 10551 2994 10557
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 8938 10588 8944 10600
rect 4724 10560 8944 10588
rect 4724 10529 4752 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 3789 10523 3847 10529
rect 3789 10489 3801 10523
rect 3835 10489 3847 10523
rect 3789 10483 3847 10489
rect 4709 10523 4767 10529
rect 4709 10489 4721 10523
rect 4755 10489 4767 10523
rect 4709 10483 4767 10489
rect 7193 10523 7251 10529
rect 7193 10489 7205 10523
rect 7239 10520 7251 10523
rect 8110 10520 8116 10532
rect 7239 10492 8116 10520
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 3007 10455 3065 10461
rect 3007 10421 3019 10455
rect 3053 10452 3065 10455
rect 3804 10452 3832 10483
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 8386 10480 8392 10532
rect 8444 10520 8450 10532
rect 8777 10523 8835 10529
rect 8777 10520 8789 10523
rect 8444 10492 8789 10520
rect 8444 10480 8450 10492
rect 8772 10489 8789 10492
rect 8823 10489 8835 10523
rect 9582 10520 9588 10532
rect 8772 10483 8835 10489
rect 8956 10492 9588 10520
rect 3053 10424 3832 10452
rect 7653 10455 7711 10461
rect 3053 10421 3065 10424
rect 3007 10415 3065 10421
rect 7653 10421 7665 10455
rect 7699 10452 7711 10455
rect 8294 10452 8300 10464
rect 7699 10424 8300 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8772 10452 8800 10483
rect 8956 10452 8984 10492
rect 9582 10480 9588 10492
rect 9640 10520 9646 10532
rect 9692 10520 9720 10619
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 10100 10560 10333 10588
rect 10100 10548 10106 10560
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10410 10548 10416 10600
rect 10468 10588 10474 10600
rect 10870 10588 10876 10600
rect 10468 10560 10876 10588
rect 10468 10548 10474 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 9640 10492 9720 10520
rect 9784 10492 10548 10520
rect 9640 10480 9646 10492
rect 9122 10452 9128 10464
rect 8772 10424 8984 10452
rect 9083 10424 9128 10452
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 9456 10424 9505 10452
rect 9456 10412 9462 10424
rect 9493 10421 9505 10424
rect 9539 10452 9551 10455
rect 9784 10452 9812 10492
rect 10520 10464 10548 10492
rect 9950 10452 9956 10464
rect 9539 10424 9812 10452
rect 9911 10424 9956 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10560 10424 10793 10452
rect 10560 10412 10566 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 1104 10362 16008 10384
rect 1104 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 10976 10362
rect 11028 10310 11040 10362
rect 11092 10310 11104 10362
rect 11156 10310 11168 10362
rect 11220 10310 16008 10362
rect 1104 10288 16008 10310
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 9122 10248 9128 10260
rect 6963 10220 9128 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10226 10248 10232 10260
rect 9999 10220 10232 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 1578 10180 1584 10192
rect 1491 10152 1584 10180
rect 1578 10140 1584 10152
rect 1636 10180 1642 10192
rect 3142 10180 3148 10192
rect 1636 10152 3148 10180
rect 1636 10140 1642 10152
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 8512 10183 8570 10189
rect 8512 10180 8524 10183
rect 8352 10152 8524 10180
rect 8352 10140 8358 10152
rect 8512 10149 8524 10152
rect 8558 10180 8570 10183
rect 8846 10180 8852 10192
rect 8558 10152 8852 10180
rect 8558 10149 8570 10152
rect 8512 10143 8570 10149
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 8312 10112 8340 10140
rect 6748 10084 8340 10112
rect 8757 10115 8815 10121
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 6748 10053 6776 10084
rect 8757 10081 8769 10115
rect 8803 10112 8815 10115
rect 9030 10112 9036 10124
rect 8803 10084 9036 10112
rect 8803 10081 8815 10084
rect 8757 10075 8815 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 9640 10084 10180 10112
rect 9640 10072 9646 10084
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 7098 10044 7104 10056
rect 6871 10016 7104 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10152 10053 10180 10084
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10060 9976 10088 10004
rect 10594 9976 10600 9988
rect 10060 9948 10600 9976
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 7282 9908 7288 9920
rect 7243 9880 7288 9908
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 7377 9911 7435 9917
rect 7377 9877 7389 9911
rect 7423 9908 7435 9911
rect 7558 9908 7564 9920
rect 7423 9880 7564 9908
rect 7423 9877 7435 9880
rect 7377 9871 7435 9877
rect 7558 9868 7564 9880
rect 7616 9908 7622 9920
rect 9306 9908 9312 9920
rect 7616 9880 9312 9908
rect 7616 9868 7622 9880
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9582 9908 9588 9920
rect 9543 9880 9588 9908
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 1104 9818 16008 9840
rect 1104 9766 3480 9818
rect 3532 9766 3544 9818
rect 3596 9766 3608 9818
rect 3660 9766 3672 9818
rect 3724 9766 8478 9818
rect 8530 9766 8542 9818
rect 8594 9766 8606 9818
rect 8658 9766 8670 9818
rect 8722 9766 13475 9818
rect 13527 9766 13539 9818
rect 13591 9766 13603 9818
rect 13655 9766 13667 9818
rect 13719 9766 16008 9818
rect 1104 9744 16008 9766
rect 7098 9704 7104 9716
rect 7059 9676 7104 9704
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 7432 9540 7573 9568
rect 7432 9528 7438 9540
rect 7561 9537 7573 9540
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 8294 9568 8300 9580
rect 7791 9540 8300 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 8846 9568 8852 9580
rect 8807 9540 8852 9568
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9582 9500 9588 9512
rect 8803 9472 9588 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 8665 9435 8723 9441
rect 8665 9401 8677 9435
rect 8711 9432 8723 9435
rect 9950 9432 9956 9444
rect 8711 9404 9956 9432
rect 8711 9401 8723 9404
rect 8665 9395 8723 9401
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 8294 9364 8300 9376
rect 8255 9336 8300 9364
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 1104 9274 16008 9296
rect 1104 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 10976 9274
rect 11028 9222 11040 9274
rect 11092 9222 11104 9274
rect 11156 9222 11168 9274
rect 11220 9222 16008 9274
rect 1104 9200 16008 9222
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7282 9160 7288 9172
rect 7147 9132 7288 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7009 9095 7067 9101
rect 7009 9061 7021 9095
rect 7055 9092 7067 9095
rect 8294 9092 8300 9104
rect 7055 9064 8300 9092
rect 7055 9061 7067 9064
rect 7009 9055 7067 9061
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 12526 9092 12532 9104
rect 12487 9064 12532 9092
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8956 7343 8959
rect 7558 8956 7564 8968
rect 7331 8928 7564 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 4212 8792 6653 8820
rect 4212 8780 4218 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 6641 8783 6699 8789
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 13449 8823 13507 8829
rect 13449 8820 13461 8823
rect 13320 8792 13461 8820
rect 13320 8780 13326 8792
rect 13449 8789 13461 8792
rect 13495 8789 13507 8823
rect 13449 8783 13507 8789
rect 1104 8730 16008 8752
rect 1104 8678 3480 8730
rect 3532 8678 3544 8730
rect 3596 8678 3608 8730
rect 3660 8678 3672 8730
rect 3724 8678 8478 8730
rect 8530 8678 8542 8730
rect 8594 8678 8606 8730
rect 8658 8678 8670 8730
rect 8722 8678 13475 8730
rect 13527 8678 13539 8730
rect 13591 8678 13603 8730
rect 13655 8678 13667 8730
rect 13719 8678 16008 8730
rect 1104 8656 16008 8678
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 1104 8186 16008 8208
rect 1104 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 10976 8186
rect 11028 8134 11040 8186
rect 11092 8134 11104 8186
rect 11156 8134 11168 8186
rect 11220 8134 16008 8186
rect 1104 8112 16008 8134
rect 1104 7642 16008 7664
rect 1104 7590 3480 7642
rect 3532 7590 3544 7642
rect 3596 7590 3608 7642
rect 3660 7590 3672 7642
rect 3724 7590 8478 7642
rect 8530 7590 8542 7642
rect 8594 7590 8606 7642
rect 8658 7590 8670 7642
rect 8722 7590 13475 7642
rect 13527 7590 13539 7642
rect 13591 7590 13603 7642
rect 13655 7590 13667 7642
rect 13719 7590 16008 7642
rect 1104 7568 16008 7590
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 9030 7392 9036 7404
rect 5500 7364 9036 7392
rect 5500 7352 5506 7364
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7324 3571 7327
rect 4154 7324 4160 7336
rect 3559 7296 4160 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 1104 7098 16008 7120
rect 1104 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 10976 7098
rect 11028 7046 11040 7098
rect 11092 7046 11104 7098
rect 11156 7046 11168 7098
rect 11220 7046 16008 7098
rect 1104 7024 16008 7046
rect 1104 6554 16008 6576
rect 1104 6502 3480 6554
rect 3532 6502 3544 6554
rect 3596 6502 3608 6554
rect 3660 6502 3672 6554
rect 3724 6502 8478 6554
rect 8530 6502 8542 6554
rect 8594 6502 8606 6554
rect 8658 6502 8670 6554
rect 8722 6502 13475 6554
rect 13527 6502 13539 6554
rect 13591 6502 13603 6554
rect 13655 6502 13667 6554
rect 13719 6502 16008 6554
rect 1104 6480 16008 6502
rect 6546 6060 6552 6112
rect 6604 6100 6610 6112
rect 9582 6100 9588 6112
rect 6604 6072 9588 6100
rect 6604 6060 6610 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 1104 6010 16008 6032
rect 1104 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 10976 6010
rect 11028 5958 11040 6010
rect 11092 5958 11104 6010
rect 11156 5958 11168 6010
rect 11220 5958 16008 6010
rect 1104 5936 16008 5958
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 3936 5868 7021 5896
rect 3936 5856 3942 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7834 5896 7840 5908
rect 7009 5859 7067 5865
rect 7208 5868 7840 5896
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 4080 5692 4108 5723
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 7208 5769 7236 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 9953 5899 10011 5905
rect 9953 5896 9965 5899
rect 9180 5868 9965 5896
rect 9180 5856 9186 5868
rect 9953 5865 9965 5868
rect 9999 5865 10011 5899
rect 14550 5896 14556 5908
rect 9953 5859 10011 5865
rect 10152 5868 14556 5896
rect 7926 5828 7932 5840
rect 7576 5800 7932 5828
rect 7576 5769 7604 5800
rect 7926 5788 7932 5800
rect 7984 5788 7990 5840
rect 10042 5828 10048 5840
rect 9232 5800 10048 5828
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6696 5732 6745 5760
rect 6696 5720 6702 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5729 7251 5763
rect 7193 5723 7251 5729
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5729 7619 5763
rect 7561 5723 7619 5729
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 9232 5760 9260 5800
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10152 5769 10180 5868
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15102 5828 15108 5840
rect 10980 5800 15108 5828
rect 10980 5769 11008 5800
rect 15102 5788 15108 5800
rect 15160 5788 15166 5840
rect 7883 5732 9260 5760
rect 9309 5763 9367 5769
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 9309 5729 9321 5763
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 9861 5763 9919 5769
rect 9861 5760 9873 5763
rect 9723 5732 9873 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 9861 5729 9873 5732
rect 9907 5729 9919 5763
rect 9861 5723 9919 5729
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5729 11023 5763
rect 11790 5760 11796 5772
rect 11751 5732 11796 5760
rect 10965 5723 11023 5729
rect 7006 5692 7012 5704
rect 4080 5664 7012 5692
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 9324 5692 9352 5723
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 13262 5692 13268 5704
rect 9324 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 4614 5584 4620 5636
rect 4672 5624 4678 5636
rect 7653 5627 7711 5633
rect 7653 5624 7665 5627
rect 4672 5596 7665 5624
rect 4672 5584 4678 5596
rect 7653 5593 7665 5596
rect 7699 5593 7711 5627
rect 7653 5587 7711 5593
rect 8202 5584 8208 5636
rect 8260 5624 8266 5636
rect 9493 5627 9551 5633
rect 9493 5624 9505 5627
rect 8260 5596 9505 5624
rect 8260 5584 8266 5596
rect 9493 5593 9505 5596
rect 9539 5593 9551 5627
rect 9493 5587 9551 5593
rect 9861 5627 9919 5633
rect 9861 5593 9873 5627
rect 9907 5624 9919 5627
rect 13998 5624 14004 5636
rect 9907 5596 14004 5624
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 13998 5584 14004 5596
rect 14056 5584 14062 5636
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 2832 5528 3893 5556
rect 2832 5516 2838 5528
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 3881 5519 3939 5525
rect 3970 5516 3976 5568
rect 4028 5556 4034 5568
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 4028 5528 6561 5556
rect 4028 5516 4034 5528
rect 6549 5525 6561 5528
rect 6595 5525 6607 5559
rect 7374 5556 7380 5568
rect 7335 5528 7380 5556
rect 6549 5519 6607 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 9125 5559 9183 5565
rect 9125 5525 9137 5559
rect 9171 5556 9183 5559
rect 9306 5556 9312 5568
rect 9171 5528 9312 5556
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10781 5559 10839 5565
rect 10781 5556 10793 5559
rect 10192 5528 10793 5556
rect 10192 5516 10198 5528
rect 10781 5525 10793 5528
rect 10827 5525 10839 5559
rect 10781 5519 10839 5525
rect 10870 5516 10876 5568
rect 10928 5556 10934 5568
rect 11609 5559 11667 5565
rect 11609 5556 11621 5559
rect 10928 5528 11621 5556
rect 10928 5516 10934 5528
rect 11609 5525 11621 5528
rect 11655 5525 11667 5559
rect 11609 5519 11667 5525
rect 1104 5466 16008 5488
rect 1104 5414 3480 5466
rect 3532 5414 3544 5466
rect 3596 5414 3608 5466
rect 3660 5414 3672 5466
rect 3724 5414 8478 5466
rect 8530 5414 8542 5466
rect 8594 5414 8606 5466
rect 8658 5414 8670 5466
rect 8722 5414 13475 5466
rect 13527 5414 13539 5466
rect 13591 5414 13603 5466
rect 13655 5414 13667 5466
rect 13719 5414 16008 5466
rect 1104 5392 16008 5414
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 6641 5355 6699 5361
rect 6641 5352 6653 5355
rect 3292 5324 6653 5352
rect 3292 5312 3298 5324
rect 6641 5321 6653 5324
rect 6687 5321 6699 5355
rect 6641 5315 6699 5321
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 8076 5324 8125 5352
rect 8076 5312 8082 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8113 5315 8171 5321
rect 8220 5324 8493 5352
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 5813 5287 5871 5293
rect 5813 5284 5825 5287
rect 2740 5256 5825 5284
rect 2740 5244 2746 5256
rect 5813 5253 5825 5256
rect 5859 5253 5871 5287
rect 7009 5287 7067 5293
rect 7009 5284 7021 5287
rect 5813 5247 5871 5253
rect 5920 5256 7021 5284
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 5920 5216 5948 5256
rect 7009 5253 7021 5256
rect 7055 5253 7067 5287
rect 7009 5247 7067 5253
rect 7926 5244 7932 5296
rect 7984 5284 7990 5296
rect 8220 5284 8248 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8849 5355 8907 5361
rect 8849 5352 8861 5355
rect 8481 5315 8539 5321
rect 8772 5324 8861 5352
rect 8772 5296 8800 5324
rect 8849 5321 8861 5324
rect 8895 5321 8907 5355
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8849 5315 8907 5321
rect 9048 5324 9137 5352
rect 9048 5296 9076 5324
rect 9125 5321 9137 5324
rect 9171 5321 9183 5355
rect 9125 5315 9183 5321
rect 9214 5312 9220 5364
rect 9272 5352 9278 5364
rect 9401 5355 9459 5361
rect 9401 5352 9413 5355
rect 9272 5324 9413 5352
rect 9272 5312 9278 5324
rect 9401 5321 9413 5324
rect 9447 5321 9459 5355
rect 9401 5315 9459 5321
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9640 5324 10057 5352
rect 9640 5312 9646 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10045 5315 10103 5321
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10376 5324 10885 5352
rect 10376 5312 10382 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 10873 5315 10931 5321
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 12032 5324 12173 5352
rect 12032 5312 12038 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12618 5352 12624 5364
rect 12579 5324 12624 5352
rect 12161 5315 12219 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 12894 5352 12900 5364
rect 12855 5324 12900 5352
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 7984 5256 8248 5284
rect 7984 5244 7990 5256
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 8573 5287 8631 5293
rect 8573 5284 8585 5287
rect 8352 5256 8585 5284
rect 8352 5244 8358 5256
rect 8573 5253 8585 5256
rect 8619 5253 8631 5287
rect 8573 5247 8631 5253
rect 8754 5244 8760 5296
rect 8812 5244 8818 5296
rect 9030 5244 9036 5296
rect 9088 5244 9094 5296
rect 9490 5244 9496 5296
rect 9548 5284 9554 5296
rect 9858 5284 9864 5296
rect 9548 5256 9864 5284
rect 9548 5244 9554 5256
rect 9858 5244 9864 5256
rect 9916 5244 9922 5296
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 10413 5287 10471 5293
rect 10413 5284 10425 5287
rect 10008 5256 10425 5284
rect 10008 5244 10014 5256
rect 10413 5253 10425 5256
rect 10459 5253 10471 5287
rect 10413 5247 10471 5253
rect 10594 5244 10600 5296
rect 10652 5284 10658 5296
rect 11149 5287 11207 5293
rect 11149 5284 11161 5287
rect 10652 5256 11161 5284
rect 10652 5244 10658 5256
rect 11149 5253 11161 5256
rect 11195 5253 11207 5287
rect 15286 5284 15292 5296
rect 11149 5247 11207 5253
rect 11900 5256 15292 5284
rect 8846 5216 8852 5228
rect 4120 5188 5948 5216
rect 8588 5188 8852 5216
rect 4120 5176 4126 5188
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 3326 5148 3332 5160
rect 1627 5120 3332 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 4890 5148 4896 5160
rect 4663 5120 4896 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5074 5148 5080 5160
rect 5031 5120 5080 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5350 5148 5356 5160
rect 5311 5120 5356 5148
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5626 5148 5632 5160
rect 5587 5120 5632 5148
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 5994 5148 6000 5160
rect 5955 5120 6000 5148
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6270 5148 6276 5160
rect 6231 5120 6276 5148
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7558 5148 7564 5160
rect 7239 5120 7564 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 7742 5148 7748 5160
rect 7699 5120 7748 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 7926 5148 7932 5160
rect 7887 5120 7932 5148
rect 7926 5108 7932 5120
rect 7984 5108 7990 5160
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5117 8355 5151
rect 8588 5148 8616 5188
rect 8846 5176 8852 5188
rect 8904 5176 8910 5228
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 11790 5216 11796 5228
rect 8996 5188 11796 5216
rect 8996 5176 9002 5188
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 8733 5151 8791 5157
rect 8733 5148 8745 5151
rect 8588 5120 8745 5148
rect 8297 5111 8355 5117
rect 8733 5117 8745 5120
rect 8779 5117 8791 5151
rect 8733 5111 8791 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 9355 5120 9505 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9766 5148 9772 5160
rect 9727 5120 9772 5148
rect 9493 5111 9551 5117
rect 1946 5040 1952 5092
rect 2004 5080 2010 5092
rect 8312 5080 8340 5111
rect 8938 5080 8944 5092
rect 2004 5052 5488 5080
rect 8312 5052 8944 5080
rect 2004 5040 2010 5052
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 4430 5012 4436 5024
rect 4391 4984 4436 5012
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 4798 5012 4804 5024
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5166 5012 5172 5024
rect 5127 4984 5172 5012
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5460 5021 5488 5052
rect 8938 5040 8944 5052
rect 8996 5040 9002 5092
rect 9048 5080 9076 5111
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10226 5148 10232 5160
rect 10187 5120 10232 5148
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5148 10655 5151
rect 10778 5148 10784 5160
rect 10643 5120 10784 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 11900 5157 11928 5256
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 14826 5216 14832 5228
rect 11992 5188 14832 5216
rect 11057 5151 11115 5157
rect 11057 5117 11069 5151
rect 11103 5148 11115 5151
rect 11333 5151 11391 5157
rect 11103 5120 11284 5148
rect 11103 5117 11115 5120
rect 11057 5111 11115 5117
rect 9398 5080 9404 5092
rect 9048 5052 9404 5080
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 11146 5080 11152 5092
rect 9508 5052 11152 5080
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 4981 5503 5015
rect 5445 4975 5503 4981
rect 6089 5015 6147 5021
rect 6089 4981 6101 5015
rect 6135 5012 6147 5015
rect 6270 5012 6276 5024
rect 6135 4984 6276 5012
rect 6135 4981 6147 4984
rect 6089 4975 6147 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 7466 5012 7472 5024
rect 7427 4984 7472 5012
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9508 5012 9536 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 9088 4984 9536 5012
rect 9585 5015 9643 5021
rect 9088 4972 9094 4984
rect 9585 4981 9597 5015
rect 9631 5012 9643 5015
rect 9674 5012 9680 5024
rect 9631 4984 9680 5012
rect 9631 4981 9643 4984
rect 9585 4975 9643 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 11256 5012 11284 5120
rect 11333 5117 11345 5151
rect 11379 5117 11391 5151
rect 11333 5111 11391 5117
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5117 11943 5151
rect 11885 5111 11943 5117
rect 11348 5080 11376 5111
rect 11992 5080 12020 5188
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 12342 5148 12348 5160
rect 12303 5120 12348 5148
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5117 12863 5151
rect 13078 5148 13084 5160
rect 13039 5120 13084 5148
rect 12805 5111 12863 5117
rect 12710 5080 12716 5092
rect 11348 5052 12020 5080
rect 12084 5052 12716 5080
rect 12084 5012 12112 5052
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 12820 5080 12848 5111
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 14918 5148 14924 5160
rect 13403 5120 14924 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15470 5080 15476 5092
rect 12820 5052 15476 5080
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 11256 4984 12112 5012
rect 12158 4972 12164 5024
rect 12216 5012 12222 5024
rect 13173 5015 13231 5021
rect 13173 5012 13185 5015
rect 12216 4984 13185 5012
rect 12216 4972 12222 4984
rect 13173 4981 13185 4984
rect 13219 4981 13231 5015
rect 13173 4975 13231 4981
rect 1104 4922 16008 4944
rect 1104 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 10976 4922
rect 11028 4870 11040 4922
rect 11092 4870 11104 4922
rect 11156 4870 11168 4922
rect 11220 4870 16008 4922
rect 1104 4848 16008 4870
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 6914 4808 6920 4820
rect 4948 4780 6920 4808
rect 4948 4768 4954 4780
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 9030 4808 9036 4820
rect 7800 4780 9036 4808
rect 7800 4768 7806 4780
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 9950 4808 9956 4820
rect 9640 4780 9956 4808
rect 9640 4768 9646 4780
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 14182 4808 14188 4820
rect 12400 4780 14188 4808
rect 12400 4768 12406 4780
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 4522 4700 4528 4752
rect 4580 4740 4586 4752
rect 7466 4740 7472 4752
rect 4580 4712 7472 4740
rect 4580 4700 4586 4712
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 7926 4700 7932 4752
rect 7984 4740 7990 4752
rect 9493 4743 9551 4749
rect 9493 4740 9505 4743
rect 7984 4712 9168 4740
rect 7984 4700 7990 4712
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 8110 4672 8116 4684
rect 5408 4644 8116 4672
rect 5408 4632 5414 4644
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 9140 4672 9168 4712
rect 9324 4712 9505 4740
rect 9324 4681 9352 4712
rect 9493 4709 9505 4712
rect 9539 4740 9551 4743
rect 10410 4740 10416 4752
rect 9539 4712 10416 4740
rect 9539 4709 9551 4712
rect 9493 4703 9551 4709
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 14826 4740 14832 4752
rect 10836 4712 14832 4740
rect 10836 4700 10842 4712
rect 14826 4700 14832 4712
rect 14884 4700 14890 4752
rect 9309 4675 9367 4681
rect 9140 4644 9260 4672
rect 8938 4564 8944 4616
rect 8996 4604 9002 4616
rect 8996 4576 9168 4604
rect 8996 4564 9002 4576
rect 9140 4545 9168 4576
rect 9125 4539 9183 4545
rect 9125 4505 9137 4539
rect 9171 4505 9183 4539
rect 9232 4536 9260 4644
rect 9309 4641 9321 4675
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 13814 4672 13820 4684
rect 9824 4644 13820 4672
rect 9824 4632 9830 4644
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 10962 4604 10968 4616
rect 9640 4576 10968 4604
rect 9640 4564 9646 4576
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11330 4564 11336 4616
rect 11388 4604 11394 4616
rect 11882 4604 11888 4616
rect 11388 4576 11888 4604
rect 11388 4564 11394 4576
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 15102 4604 15108 4616
rect 12768 4576 15108 4604
rect 12768 4564 12774 4576
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 12066 4536 12072 4548
rect 9232 4508 12072 4536
rect 9125 4499 9183 4505
rect 12066 4496 12072 4508
rect 12124 4496 12130 4548
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 9674 4468 9680 4480
rect 5868 4440 9680 4468
rect 5868 4428 5874 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 14550 4468 14556 4480
rect 10284 4440 14556 4468
rect 10284 4428 10290 4440
rect 14550 4428 14556 4440
rect 14608 4428 14614 4480
rect 1104 4378 16008 4400
rect 1104 4326 3480 4378
rect 3532 4326 3544 4378
rect 3596 4326 3608 4378
rect 3660 4326 3672 4378
rect 3724 4326 8478 4378
rect 8530 4326 8542 4378
rect 8594 4326 8606 4378
rect 8658 4326 8670 4378
rect 8722 4326 13475 4378
rect 13527 4326 13539 4378
rect 13591 4326 13603 4378
rect 13655 4326 13667 4378
rect 13719 4326 16008 4378
rect 1104 4304 16008 4326
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 13262 4264 13268 4276
rect 9272 4236 13268 4264
rect 9272 4224 9278 4236
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 7558 4156 7564 4208
rect 7616 4196 7622 4208
rect 7616 4168 11376 4196
rect 7616 4156 7622 4168
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 9398 4128 9404 4140
rect 7248 4100 9404 4128
rect 7248 4088 7254 4100
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 11348 4128 11376 4168
rect 11422 4156 11428 4208
rect 11480 4196 11486 4208
rect 12158 4196 12164 4208
rect 11480 4168 12164 4196
rect 11480 4156 11486 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 11514 4128 11520 4140
rect 11348 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 1104 3834 16008 3856
rect 1104 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 10976 3834
rect 11028 3782 11040 3834
rect 11092 3782 11104 3834
rect 11156 3782 11168 3834
rect 11220 3782 16008 3834
rect 1104 3760 16008 3782
rect 15013 3723 15071 3729
rect 15013 3689 15025 3723
rect 15059 3720 15071 3723
rect 15194 3720 15200 3732
rect 15059 3692 15200 3720
rect 15059 3689 15071 3692
rect 15013 3683 15071 3689
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 15470 3720 15476 3732
rect 15431 3692 15476 3720
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15197 3587 15255 3593
rect 15197 3553 15209 3587
rect 15243 3584 15255 3587
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 15243 3556 15669 3584
rect 15243 3553 15255 3556
rect 15197 3547 15255 3553
rect 15657 3553 15669 3556
rect 15703 3584 15715 3587
rect 16942 3584 16948 3596
rect 15703 3556 16948 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 15378 3380 15384 3392
rect 15339 3352 15384 3380
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 1104 3290 16008 3312
rect 1104 3238 3480 3290
rect 3532 3238 3544 3290
rect 3596 3238 3608 3290
rect 3660 3238 3672 3290
rect 3724 3238 8478 3290
rect 8530 3238 8542 3290
rect 8594 3238 8606 3290
rect 8658 3238 8670 3290
rect 8722 3238 13475 3290
rect 13527 3238 13539 3290
rect 13591 3238 13603 3290
rect 13655 3238 13667 3290
rect 13719 3238 16008 3290
rect 1104 3216 16008 3238
rect 1394 3176 1400 3188
rect 1355 3148 1400 3176
rect 1394 3136 1400 3148
rect 1452 3136 1458 3188
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3176 15255 3179
rect 15286 3176 15292 3188
rect 15243 3148 15292 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 5626 3068 5632 3120
rect 5684 3108 5690 3120
rect 9214 3108 9220 3120
rect 5684 3080 9220 3108
rect 5684 3068 5690 3080
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 14093 3111 14151 3117
rect 14093 3077 14105 3111
rect 14139 3108 14151 3111
rect 14274 3108 14280 3120
rect 14139 3080 14280 3108
rect 14139 3077 14151 3080
rect 14093 3071 14151 3077
rect 14274 3068 14280 3080
rect 14332 3108 14338 3120
rect 16482 3108 16488 3120
rect 14332 3080 16488 3108
rect 14332 3068 14338 3080
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 8202 3040 8208 3052
rect 5592 3012 8208 3040
rect 5592 3000 5598 3012
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 14921 3043 14979 3049
rect 10376 3012 12756 3040
rect 10376 3000 10382 3012
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2972 1639 2975
rect 1627 2944 1716 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 1688 2848 1716 2944
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 5626 2972 5632 2984
rect 3200 2944 5632 2972
rect 3200 2932 3206 2944
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 9122 2972 9128 2984
rect 7800 2944 9128 2972
rect 7800 2932 7806 2944
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 12728 2972 12756 3012
rect 14921 3009 14933 3043
rect 14967 3040 14979 3043
rect 14967 3012 15608 3040
rect 14967 3009 14979 3012
rect 14921 3003 14979 3009
rect 15580 2984 15608 3012
rect 15105 2975 15163 2981
rect 12728 2944 14320 2972
rect 3789 2907 3847 2913
rect 3789 2873 3801 2907
rect 3835 2873 3847 2907
rect 4062 2904 4068 2916
rect 4023 2876 4068 2904
rect 3789 2867 3847 2873
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 3694 2836 3700 2848
rect 3655 2808 3700 2836
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 3804 2836 3832 2867
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 4249 2907 4307 2913
rect 4249 2873 4261 2907
rect 4295 2904 4307 2907
rect 8846 2904 8852 2916
rect 4295 2876 8852 2904
rect 4295 2873 4307 2876
rect 4249 2867 4307 2873
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 13906 2864 13912 2916
rect 13964 2904 13970 2916
rect 14185 2907 14243 2913
rect 14185 2904 14197 2907
rect 13964 2876 14197 2904
rect 13964 2864 13970 2876
rect 14185 2873 14197 2876
rect 14231 2873 14243 2907
rect 14292 2904 14320 2944
rect 15105 2941 15117 2975
rect 15151 2972 15163 2975
rect 15194 2972 15200 2984
rect 15151 2944 15200 2972
rect 15151 2941 15163 2944
rect 15105 2935 15163 2941
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 15378 2932 15384 2984
rect 15436 2972 15442 2984
rect 15436 2944 15529 2972
rect 15436 2932 15442 2944
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 15657 2975 15715 2981
rect 15657 2972 15669 2975
rect 15620 2944 15669 2972
rect 15620 2932 15626 2944
rect 15657 2941 15669 2944
rect 15703 2941 15715 2975
rect 15657 2935 15715 2941
rect 15396 2904 15424 2932
rect 16022 2904 16028 2916
rect 14292 2876 14872 2904
rect 15396 2876 16028 2904
rect 14185 2867 14243 2873
rect 8294 2836 8300 2848
rect 3804 2808 8300 2836
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 9640 2808 9873 2836
rect 9640 2796 9646 2808
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 9861 2799 9919 2805
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 11149 2839 11207 2845
rect 11149 2836 11161 2839
rect 10928 2808 11161 2836
rect 10928 2796 10934 2808
rect 11149 2805 11161 2808
rect 11195 2805 11207 2839
rect 11790 2836 11796 2848
rect 11751 2808 11796 2836
rect 11149 2799 11207 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12618 2796 12624 2848
rect 12676 2836 12682 2848
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12676 2808 12909 2836
rect 12676 2796 12682 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 12897 2799 12955 2805
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 13817 2839 13875 2845
rect 13817 2836 13829 2839
rect 13412 2808 13829 2836
rect 13412 2796 13418 2808
rect 13817 2805 13829 2808
rect 13863 2805 13875 2839
rect 14366 2836 14372 2848
rect 14327 2808 14372 2836
rect 13817 2799 13875 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 14734 2836 14740 2848
rect 14695 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 14844 2836 14872 2876
rect 16022 2864 16028 2876
rect 16080 2864 16086 2916
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 14844 2808 15485 2836
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 1104 2746 16008 2768
rect 1104 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 10976 2746
rect 11028 2694 11040 2746
rect 11092 2694 11104 2746
rect 11156 2694 11168 2746
rect 11220 2694 16008 2746
rect 1104 2672 16008 2694
rect 2774 2632 2780 2644
rect 1412 2604 2780 2632
rect 1412 2496 1440 2604
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 4430 2632 4436 2644
rect 3620 2604 4436 2632
rect 1486 2524 1492 2576
rect 1544 2564 1550 2576
rect 2501 2567 2559 2573
rect 2501 2564 2513 2567
rect 1544 2536 2513 2564
rect 1544 2524 1550 2536
rect 2501 2533 2513 2536
rect 2547 2533 2559 2567
rect 3620 2564 3648 2604
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 7742 2632 7748 2644
rect 6196 2604 7748 2632
rect 2501 2527 2559 2533
rect 2608 2536 3648 2564
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1412 2468 1593 2496
rect 1581 2465 1593 2468
rect 1627 2465 1639 2499
rect 1581 2459 1639 2465
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2038 2496 2044 2508
rect 1995 2468 2044 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2608 2496 2636 2536
rect 3878 2524 3884 2576
rect 3936 2564 3942 2576
rect 4065 2567 4123 2573
rect 4065 2564 4077 2567
rect 3936 2536 4077 2564
rect 3936 2524 3942 2536
rect 4065 2533 4077 2536
rect 4111 2533 4123 2567
rect 4614 2564 4620 2576
rect 4575 2536 4620 2564
rect 4065 2527 4123 2533
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 5534 2564 5540 2576
rect 5495 2536 5540 2564
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 6089 2567 6147 2573
rect 6089 2564 6101 2567
rect 5684 2536 6101 2564
rect 5684 2524 5690 2536
rect 6089 2533 6101 2536
rect 6135 2533 6147 2567
rect 6089 2527 6147 2533
rect 2363 2468 2636 2496
rect 2685 2499 2743 2505
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 2958 2496 2964 2508
rect 2731 2468 2964 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 3053 2499 3111 2505
rect 3053 2465 3065 2499
rect 3099 2496 3111 2499
rect 3326 2496 3332 2508
rect 3099 2468 3332 2496
rect 3099 2465 3111 2468
rect 3053 2459 3111 2465
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 3970 2496 3976 2508
rect 3467 2468 3976 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3970 2456 3976 2468
rect 4028 2456 4034 2508
rect 5074 2496 5080 2508
rect 5035 2468 5080 2496
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5905 2499 5963 2505
rect 5905 2465 5917 2499
rect 5951 2496 5963 2499
rect 6196 2496 6224 2604
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 8757 2635 8815 2641
rect 8757 2632 8769 2635
rect 7892 2604 8769 2632
rect 7892 2592 7898 2604
rect 8757 2601 8769 2604
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 8938 2592 8944 2644
rect 8996 2592 9002 2644
rect 9214 2632 9220 2644
rect 9175 2604 9220 2632
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 9456 2604 9597 2632
rect 9456 2592 9462 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9585 2595 9643 2601
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10045 2635 10103 2641
rect 10045 2632 10057 2635
rect 10008 2604 10057 2632
rect 10008 2592 10014 2604
rect 10045 2601 10057 2604
rect 10091 2601 10103 2635
rect 10045 2595 10103 2601
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10686 2632 10692 2644
rect 10284 2604 10692 2632
rect 10284 2592 10290 2604
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10836 2604 10885 2632
rect 10836 2592 10842 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11514 2632 11520 2644
rect 11379 2604 11520 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12894 2632 12900 2644
rect 12176 2604 12900 2632
rect 6273 2567 6331 2573
rect 6273 2533 6285 2567
rect 6319 2564 6331 2567
rect 7374 2564 7380 2576
rect 6319 2536 7380 2564
rect 6319 2533 6331 2536
rect 6273 2527 6331 2533
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 7469 2567 7527 2573
rect 7469 2533 7481 2567
rect 7515 2564 7527 2567
rect 8956 2564 8984 2592
rect 10321 2567 10379 2573
rect 10321 2564 10333 2567
rect 7515 2536 8984 2564
rect 9416 2536 10333 2564
rect 7515 2533 7527 2536
rect 7469 2527 7527 2533
rect 6730 2496 6736 2508
rect 5951 2468 6224 2496
rect 6691 2468 6736 2496
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7098 2496 7104 2508
rect 7059 2468 7104 2496
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8205 2499 8263 2505
rect 7883 2468 8156 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 1026 2388 1032 2440
rect 1084 2428 1090 2440
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 1084 2400 2145 2428
rect 1084 2388 1090 2400
rect 2133 2397 2145 2400
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 2832 2400 3893 2428
rect 2832 2388 2838 2400
rect 3881 2397 3893 2400
rect 3927 2397 3939 2431
rect 5166 2428 5172 2440
rect 3881 2391 3939 2397
rect 3988 2400 5172 2428
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 256 2332 1409 2360
rect 256 2320 262 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2314 2320 2320 2372
rect 2372 2360 2378 2372
rect 3237 2363 3295 2369
rect 3237 2360 3249 2363
rect 2372 2332 3249 2360
rect 2372 2320 2378 2332
rect 3237 2329 3249 2332
rect 3283 2329 3295 2363
rect 3237 2323 3295 2329
rect 3326 2320 3332 2372
rect 3384 2360 3390 2372
rect 3988 2360 4016 2400
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 6638 2388 6644 2440
rect 6696 2428 6702 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6696 2400 6929 2428
rect 6696 2388 6702 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7064 2400 7297 2428
rect 7064 2388 7070 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 4430 2360 4436 2372
rect 3384 2332 4016 2360
rect 4391 2332 4436 2360
rect 3384 2320 3390 2332
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 4890 2360 4896 2372
rect 4851 2332 4896 2360
rect 4890 2320 4896 2332
rect 4948 2320 4954 2372
rect 5350 2360 5356 2372
rect 5311 2332 5356 2360
rect 5350 2320 5356 2332
rect 5408 2320 5414 2372
rect 5718 2360 5724 2372
rect 5679 2332 5724 2360
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 6178 2320 6184 2372
rect 6236 2360 6242 2372
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 6236 2332 6561 2360
rect 6236 2320 6242 2332
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 6549 2323 6607 2329
rect 7466 2320 7472 2372
rect 7524 2360 7530 2372
rect 7653 2363 7711 2369
rect 7653 2360 7665 2363
rect 7524 2332 7665 2360
rect 7524 2320 7530 2332
rect 7653 2329 7665 2332
rect 7699 2329 7711 2363
rect 7653 2323 7711 2329
rect 7926 2320 7932 2372
rect 7984 2360 7990 2372
rect 8021 2363 8079 2369
rect 8021 2360 8033 2363
rect 7984 2332 8033 2360
rect 7984 2320 7990 2332
rect 8021 2329 8033 2332
rect 8067 2329 8079 2363
rect 8021 2323 8079 2329
rect 566 2252 572 2304
rect 624 2292 630 2304
rect 1857 2295 1915 2301
rect 1857 2292 1869 2295
rect 624 2264 1869 2292
rect 624 2252 630 2264
rect 1857 2261 1869 2264
rect 1903 2261 1915 2295
rect 1857 2255 1915 2261
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 2004 2264 2973 2292
rect 2004 2252 2010 2264
rect 2961 2261 2973 2264
rect 3007 2261 3019 2295
rect 2961 2255 3019 2261
rect 3050 2252 3056 2304
rect 3108 2292 3114 2304
rect 6270 2292 6276 2304
rect 3108 2264 6276 2292
rect 3108 2252 3114 2264
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 8128 2292 8156 2468
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 8573 2499 8631 2505
rect 8251 2468 8524 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 8352 2332 8401 2360
rect 8352 2320 8358 2332
rect 8389 2329 8401 2332
rect 8435 2329 8447 2363
rect 8496 2360 8524 2468
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 8754 2496 8760 2508
rect 8619 2468 8760 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 8941 2499 8999 2505
rect 8941 2465 8953 2499
rect 8987 2496 8999 2499
rect 8987 2468 9076 2496
rect 8987 2465 8999 2468
rect 8941 2459 8999 2465
rect 9048 2440 9076 2468
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 9416 2505 9444 2536
rect 10321 2533 10333 2536
rect 10367 2533 10379 2567
rect 11609 2567 11667 2573
rect 11609 2564 11621 2567
rect 10321 2527 10379 2533
rect 10704 2536 11621 2564
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 9272 2468 9413 2496
rect 9272 2456 9278 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9732 2468 9781 2496
rect 9732 2456 9738 2468
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 10042 2456 10048 2508
rect 10100 2496 10106 2508
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 10100 2468 10241 2496
rect 10100 2456 10106 2468
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9088 2400 9873 2428
rect 9088 2388 9094 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 10244 2428 10272 2459
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 10704 2505 10732 2536
rect 11609 2533 11621 2536
rect 11655 2533 11667 2567
rect 12176 2564 12204 2604
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13320 2604 13461 2632
rect 13320 2592 13326 2604
rect 13449 2601 13461 2604
rect 13495 2601 13507 2635
rect 13449 2595 13507 2601
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 13909 2635 13967 2641
rect 13909 2632 13921 2635
rect 13872 2604 13921 2632
rect 13872 2592 13878 2604
rect 13909 2601 13921 2604
rect 13955 2601 13967 2635
rect 14182 2632 14188 2644
rect 14143 2604 14188 2632
rect 13909 2595 13967 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14550 2632 14556 2644
rect 14511 2604 14556 2632
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14826 2632 14832 2644
rect 14787 2604 14832 2632
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 15102 2632 15108 2644
rect 15063 2604 15108 2632
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 15344 2604 15516 2632
rect 15344 2592 15350 2604
rect 15488 2573 15516 2604
rect 12437 2567 12495 2573
rect 12437 2564 12449 2567
rect 11609 2527 11667 2533
rect 11716 2536 12204 2564
rect 12268 2536 12449 2564
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10560 2468 10701 2496
rect 10560 2456 10566 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 11054 2496 11060 2508
rect 11015 2468 11060 2496
rect 10689 2459 10747 2465
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11388 2468 11529 2496
rect 11388 2456 11394 2468
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 10244 2400 11161 2428
rect 9861 2391 9919 2397
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11716 2360 11744 2536
rect 12268 2508 12296 2536
rect 12437 2533 12449 2536
rect 12483 2533 12495 2567
rect 12437 2527 12495 2533
rect 15473 2567 15531 2573
rect 15473 2533 15485 2567
rect 15519 2533 15531 2567
rect 15473 2527 15531 2533
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11848 2468 12081 2496
rect 11848 2456 11854 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 12158 2456 12164 2508
rect 12216 2456 12222 2508
rect 12250 2456 12256 2508
rect 12308 2456 12314 2508
rect 12345 2499 12403 2505
rect 12345 2465 12357 2499
rect 12391 2496 12403 2499
rect 12391 2468 12425 2496
rect 12391 2465 12403 2468
rect 12345 2459 12403 2465
rect 12176 2428 12204 2456
rect 12360 2428 12388 2459
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 12805 2499 12863 2505
rect 12805 2496 12817 2499
rect 12676 2468 12817 2496
rect 12676 2456 12682 2468
rect 12805 2465 12817 2468
rect 12851 2465 12863 2499
rect 12805 2459 12863 2465
rect 13078 2456 13084 2508
rect 13136 2496 13142 2508
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 13136 2468 13277 2496
rect 13136 2456 13142 2468
rect 13265 2465 13277 2468
rect 13311 2465 13323 2499
rect 13265 2459 13323 2465
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12176 2400 12909 2428
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 13280 2428 13308 2459
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 13412 2468 13645 2496
rect 13412 2456 13418 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 13964 2468 14105 2496
rect 13964 2456 13970 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14274 2456 14280 2508
rect 14332 2496 14338 2508
rect 14369 2499 14427 2505
rect 14369 2496 14381 2499
rect 14332 2468 14381 2496
rect 14332 2456 14338 2468
rect 14369 2465 14381 2468
rect 14415 2465 14427 2499
rect 14369 2459 14427 2465
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14516 2468 14749 2496
rect 14516 2456 14522 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 14826 2456 14832 2508
rect 14884 2496 14890 2508
rect 15013 2499 15071 2505
rect 15013 2496 15025 2499
rect 14884 2468 15025 2496
rect 14884 2456 14890 2468
rect 15013 2465 15025 2468
rect 15059 2465 15071 2499
rect 15013 2459 15071 2465
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 15252 2468 15301 2496
rect 15252 2456 15258 2468
rect 15289 2465 15301 2468
rect 15335 2465 15347 2499
rect 15654 2496 15660 2508
rect 15615 2468 15660 2496
rect 15289 2459 15347 2465
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 13725 2431 13783 2437
rect 13725 2428 13737 2431
rect 13280 2400 13737 2428
rect 12897 2391 12955 2397
rect 13725 2397 13737 2400
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 8496 2332 11744 2360
rect 8389 2323 8447 2329
rect 12066 2320 12072 2372
rect 12124 2360 12130 2372
rect 12161 2363 12219 2369
rect 12161 2360 12173 2363
rect 12124 2332 12173 2360
rect 12124 2320 12130 2332
rect 12161 2329 12173 2332
rect 12207 2329 12219 2363
rect 12161 2323 12219 2329
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 12492 2332 12633 2360
rect 12492 2320 12498 2332
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 12621 2323 12679 2329
rect 10226 2292 10232 2304
rect 8128 2264 10232 2292
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 10410 2252 10416 2304
rect 10468 2292 10474 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10468 2264 10517 2292
rect 10468 2252 10474 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 11330 2252 11336 2304
rect 11388 2292 11394 2304
rect 12250 2292 12256 2304
rect 11388 2264 12256 2292
rect 11388 2252 11394 2264
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 12986 2252 12992 2304
rect 13044 2292 13050 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 13044 2264 13093 2292
rect 13044 2252 13050 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13081 2255 13139 2261
rect 1104 2202 16008 2224
rect 1104 2150 3480 2202
rect 3532 2150 3544 2202
rect 3596 2150 3608 2202
rect 3660 2150 3672 2202
rect 3724 2150 8478 2202
rect 8530 2150 8542 2202
rect 8594 2150 8606 2202
rect 8658 2150 8670 2202
rect 8722 2150 13475 2202
rect 13527 2150 13539 2202
rect 13591 2150 13603 2202
rect 13655 2150 13667 2202
rect 13719 2150 16008 2202
rect 1104 2128 16008 2150
rect 2038 2048 2044 2100
rect 2096 2088 2102 2100
rect 4798 2088 4804 2100
rect 2096 2060 4804 2088
rect 2096 2048 2102 2060
rect 4798 2048 4804 2060
rect 4856 2048 4862 2100
rect 8938 2048 8944 2100
rect 8996 2088 9002 2100
rect 11422 2088 11428 2100
rect 8996 2060 11428 2088
rect 8996 2048 9002 2060
rect 11422 2048 11428 2060
rect 11480 2048 11486 2100
rect 12986 2088 12992 2100
rect 12406 2060 12992 2088
rect 7098 1980 7104 2032
rect 7156 2020 7162 2032
rect 10134 2020 10140 2032
rect 7156 1992 10140 2020
rect 7156 1980 7162 1992
rect 10134 1980 10140 1992
rect 10192 1980 10198 2032
rect 10318 1980 10324 2032
rect 10376 2020 10382 2032
rect 12406 2020 12434 2060
rect 12986 2048 12992 2060
rect 13044 2048 13050 2100
rect 10376 1992 12434 2020
rect 10376 1980 10382 1992
rect 5074 1844 5080 1896
rect 5132 1884 5138 1896
rect 9306 1884 9312 1896
rect 5132 1856 9312 1884
rect 5132 1844 5138 1856
rect 9306 1844 9312 1856
rect 9364 1844 9370 1896
rect 6730 1776 6736 1828
rect 6788 1816 6794 1828
rect 10594 1816 10600 1828
rect 6788 1788 10600 1816
rect 6788 1776 6794 1788
rect 10594 1776 10600 1788
rect 10652 1776 10658 1828
rect 7650 1708 7656 1760
rect 7708 1748 7714 1760
rect 10410 1748 10416 1760
rect 7708 1720 10416 1748
rect 7708 1708 7714 1720
rect 10410 1708 10416 1720
rect 10468 1708 10474 1760
<< via1 >>
rect 8300 17892 8352 17944
rect 11980 17892 12032 17944
rect 6276 17824 6328 17876
rect 10508 17824 10560 17876
rect 7840 17756 7892 17808
rect 11796 17756 11848 17808
rect 9220 17688 9272 17740
rect 12256 17688 12308 17740
rect 7380 17620 7432 17672
rect 10324 17620 10376 17672
rect 8208 17552 8260 17604
rect 11428 17552 11480 17604
rect 4160 17484 4212 17536
rect 9312 17484 9364 17536
rect 9496 17484 9548 17536
rect 11612 17484 11664 17536
rect 15568 17484 15620 17536
rect 16120 17484 16172 17536
rect 3480 17382 3532 17434
rect 3544 17382 3596 17434
rect 3608 17382 3660 17434
rect 3672 17382 3724 17434
rect 8478 17382 8530 17434
rect 8542 17382 8594 17434
rect 8606 17382 8658 17434
rect 8670 17382 8722 17434
rect 13475 17382 13527 17434
rect 13539 17382 13591 17434
rect 13603 17382 13655 17434
rect 13667 17382 13719 17434
rect 1032 17280 1084 17332
rect 2228 17280 2280 17332
rect 3056 17280 3108 17332
rect 4344 17280 4396 17332
rect 8852 17280 8904 17332
rect 9312 17323 9364 17332
rect 9312 17289 9321 17323
rect 9321 17289 9355 17323
rect 9355 17289 9364 17323
rect 9312 17280 9364 17289
rect 9588 17280 9640 17332
rect 11612 17280 11664 17332
rect 572 17212 624 17264
rect 2780 17212 2832 17264
rect 3792 17212 3844 17264
rect 4804 17255 4856 17264
rect 4804 17221 4813 17255
rect 4813 17221 4847 17255
rect 4847 17221 4856 17255
rect 4804 17212 4856 17221
rect 5172 17255 5224 17264
rect 5172 17221 5181 17255
rect 5181 17221 5215 17255
rect 5215 17221 5224 17255
rect 5172 17212 5224 17221
rect 5632 17255 5684 17264
rect 5632 17221 5641 17255
rect 5641 17221 5675 17255
rect 5675 17221 5684 17255
rect 5632 17212 5684 17221
rect 6000 17255 6052 17264
rect 6000 17221 6009 17255
rect 6009 17221 6043 17255
rect 6043 17221 6052 17255
rect 6000 17212 6052 17221
rect 6460 17212 6512 17264
rect 6920 17255 6972 17264
rect 6920 17221 6929 17255
rect 6929 17221 6963 17255
rect 6963 17221 6972 17255
rect 7288 17255 7340 17264
rect 6920 17212 6972 17221
rect 7288 17221 7297 17255
rect 7297 17221 7331 17255
rect 7331 17221 7340 17255
rect 7288 17212 7340 17221
rect 7748 17255 7800 17264
rect 7748 17221 7757 17255
rect 7757 17221 7791 17255
rect 7791 17221 7800 17255
rect 7748 17212 7800 17221
rect 8116 17255 8168 17264
rect 8116 17221 8125 17255
rect 8125 17221 8159 17255
rect 8159 17221 8168 17255
rect 8116 17212 8168 17221
rect 1860 17144 1912 17196
rect 5080 17144 5132 17196
rect 10324 17212 10376 17264
rect 10600 17212 10652 17264
rect 15660 17255 15712 17264
rect 15660 17221 15669 17255
rect 15669 17221 15703 17255
rect 15703 17221 15712 17255
rect 15660 17212 15712 17221
rect 9772 17144 9824 17196
rect 1400 17076 1452 17128
rect 4528 17076 4580 17128
rect 8668 17076 8720 17128
rect 9680 17076 9732 17128
rect 10140 17119 10192 17128
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 11060 17144 11112 17196
rect 11336 17144 11388 17196
rect 1584 17051 1636 17060
rect 1584 17017 1593 17051
rect 1593 17017 1627 17051
rect 1627 17017 1636 17051
rect 1584 17008 1636 17017
rect 1952 17051 2004 17060
rect 1952 17017 1961 17051
rect 1961 17017 1995 17051
rect 1995 17017 2004 17051
rect 1952 17008 2004 17017
rect 2688 17051 2740 17060
rect 2688 17017 2697 17051
rect 2697 17017 2731 17051
rect 2731 17017 2740 17051
rect 2688 17008 2740 17017
rect 3240 17008 3292 17060
rect 4068 17051 4120 17060
rect 4068 17017 4077 17051
rect 4077 17017 4111 17051
rect 4111 17017 4120 17051
rect 4068 17008 4120 17017
rect 4436 17051 4488 17060
rect 4436 17017 4445 17051
rect 4445 17017 4479 17051
rect 4479 17017 4488 17051
rect 4436 17008 4488 17017
rect 4988 17051 5040 17060
rect 4988 17017 4997 17051
rect 4997 17017 5031 17051
rect 5031 17017 5040 17051
rect 4988 17008 5040 17017
rect 5356 17051 5408 17060
rect 5356 17017 5365 17051
rect 5365 17017 5399 17051
rect 5399 17017 5408 17051
rect 5356 17008 5408 17017
rect 5816 17051 5868 17060
rect 5816 17017 5825 17051
rect 5825 17017 5859 17051
rect 5859 17017 5868 17051
rect 5816 17008 5868 17017
rect 6552 17008 6604 17060
rect 6736 17051 6788 17060
rect 6736 17017 6745 17051
rect 6745 17017 6779 17051
rect 6779 17017 6788 17051
rect 6736 17008 6788 17017
rect 7472 17051 7524 17060
rect 7472 17017 7481 17051
rect 7481 17017 7515 17051
rect 7515 17017 7524 17051
rect 7472 17008 7524 17017
rect 8116 17008 8168 17060
rect 8300 17051 8352 17060
rect 8300 17017 8309 17051
rect 8309 17017 8343 17051
rect 8343 17017 8352 17051
rect 8300 17008 8352 17017
rect 5264 16940 5316 16992
rect 8024 16940 8076 16992
rect 10048 17008 10100 17060
rect 10232 17008 10284 17060
rect 11152 17076 11204 17128
rect 11888 17144 11940 17196
rect 11612 17076 11664 17128
rect 12440 17076 12492 17128
rect 12716 17076 12768 17128
rect 13176 17076 13228 17128
rect 13452 17076 13504 17128
rect 14004 17076 14056 17128
rect 14372 17076 14424 17128
rect 14464 17076 14516 17128
rect 14832 17076 14884 17128
rect 15292 17119 15344 17128
rect 15292 17085 15301 17119
rect 15301 17085 15335 17119
rect 15335 17085 15344 17119
rect 15292 17076 15344 17085
rect 15476 17051 15528 17060
rect 15476 17017 15485 17051
rect 15485 17017 15519 17051
rect 15519 17017 15528 17051
rect 15476 17008 15528 17017
rect 8852 16940 8904 16992
rect 10508 16940 10560 16992
rect 11428 16940 11480 16992
rect 11796 16940 11848 16992
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 12256 16940 12308 16992
rect 13360 16940 13412 16992
rect 14004 16983 14056 16992
rect 14004 16949 14013 16983
rect 14013 16949 14047 16983
rect 14047 16949 14056 16983
rect 14004 16940 14056 16949
rect 14556 16983 14608 16992
rect 14556 16949 14565 16983
rect 14565 16949 14599 16983
rect 14599 16949 14608 16983
rect 14556 16940 14608 16949
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 15108 16983 15160 16992
rect 15108 16949 15117 16983
rect 15117 16949 15151 16983
rect 15151 16949 15160 16983
rect 15108 16940 15160 16949
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 10976 16838 11028 16890
rect 11040 16838 11092 16890
rect 11104 16838 11156 16890
rect 11168 16838 11220 16890
rect 2780 16736 2832 16788
rect 6644 16736 6696 16788
rect 9588 16736 9640 16788
rect 204 16600 256 16652
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 3976 16668 4028 16720
rect 7748 16668 7800 16720
rect 8852 16668 8904 16720
rect 8116 16600 8168 16652
rect 10416 16736 10468 16788
rect 11336 16736 11388 16788
rect 11520 16736 11572 16788
rect 11888 16736 11940 16788
rect 12716 16736 12768 16788
rect 14372 16779 14424 16788
rect 14372 16745 14381 16779
rect 14381 16745 14415 16779
rect 14415 16745 14424 16779
rect 14372 16736 14424 16745
rect 14464 16736 14516 16788
rect 14740 16779 14792 16788
rect 14740 16745 14749 16779
rect 14749 16745 14783 16779
rect 14783 16745 14792 16779
rect 14740 16736 14792 16745
rect 10140 16668 10192 16720
rect 9772 16600 9824 16652
rect 11612 16668 11664 16720
rect 11796 16668 11848 16720
rect 10784 16600 10836 16652
rect 12164 16600 12216 16652
rect 10876 16532 10928 16584
rect 8944 16464 8996 16516
rect 10140 16464 10192 16516
rect 10232 16464 10284 16516
rect 15016 16532 15068 16584
rect 15568 16600 15620 16652
rect 15752 16600 15804 16652
rect 16948 16532 17000 16584
rect 9404 16396 9456 16448
rect 10416 16396 10468 16448
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 3480 16294 3532 16346
rect 3544 16294 3596 16346
rect 3608 16294 3660 16346
rect 3672 16294 3724 16346
rect 8478 16294 8530 16346
rect 8542 16294 8594 16346
rect 8606 16294 8658 16346
rect 8670 16294 8722 16346
rect 13475 16294 13527 16346
rect 13539 16294 13591 16346
rect 13603 16294 13655 16346
rect 13667 16294 13719 16346
rect 9680 16192 9732 16244
rect 12624 16192 12676 16244
rect 15016 16192 15068 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 15752 16124 15804 16176
rect 16488 15988 16540 16040
rect 13084 15852 13136 15904
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 10976 15750 11028 15802
rect 11040 15750 11092 15802
rect 11104 15750 11156 15802
rect 11168 15750 11220 15802
rect 15568 15691 15620 15700
rect 15568 15657 15577 15691
rect 15577 15657 15611 15691
rect 15611 15657 15620 15691
rect 15568 15648 15620 15657
rect 3480 15206 3532 15258
rect 3544 15206 3596 15258
rect 3608 15206 3660 15258
rect 3672 15206 3724 15258
rect 8478 15206 8530 15258
rect 8542 15206 8594 15258
rect 8606 15206 8658 15258
rect 8670 15206 8722 15258
rect 13475 15206 13527 15258
rect 13539 15206 13591 15258
rect 13603 15206 13655 15258
rect 13667 15206 13719 15258
rect 1584 15104 1636 15156
rect 4528 15147 4580 15156
rect 4528 15113 4537 15147
rect 4537 15113 4571 15147
rect 4571 15113 4580 15147
rect 4528 15104 4580 15113
rect 5264 15104 5316 15156
rect 4988 15036 5040 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 1768 14832 1820 14884
rect 7104 14832 7156 14884
rect 7564 14832 7616 14884
rect 7288 14764 7340 14816
rect 9404 14764 9456 14816
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 10976 14662 11028 14714
rect 11040 14662 11092 14714
rect 11104 14662 11156 14714
rect 11168 14662 11220 14714
rect 7472 14560 7524 14612
rect 9956 14424 10008 14476
rect 3480 14118 3532 14170
rect 3544 14118 3596 14170
rect 3608 14118 3660 14170
rect 3672 14118 3724 14170
rect 8478 14118 8530 14170
rect 8542 14118 8594 14170
rect 8606 14118 8658 14170
rect 8670 14118 8722 14170
rect 13475 14118 13527 14170
rect 13539 14118 13591 14170
rect 13603 14118 13655 14170
rect 13667 14118 13719 14170
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 10976 13574 11028 13626
rect 11040 13574 11092 13626
rect 11104 13574 11156 13626
rect 11168 13574 11220 13626
rect 15476 13472 15528 13524
rect 3976 13404 4028 13456
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 5540 13336 5592 13388
rect 15200 13336 15252 13388
rect 3148 13132 3200 13184
rect 9588 13200 9640 13252
rect 7012 13132 7064 13184
rect 15200 13175 15252 13184
rect 15200 13141 15209 13175
rect 15209 13141 15243 13175
rect 15243 13141 15252 13175
rect 15200 13132 15252 13141
rect 3480 13030 3532 13082
rect 3544 13030 3596 13082
rect 3608 13030 3660 13082
rect 3672 13030 3724 13082
rect 8478 13030 8530 13082
rect 8542 13030 8594 13082
rect 8606 13030 8658 13082
rect 8670 13030 8722 13082
rect 13475 13030 13527 13082
rect 13539 13030 13591 13082
rect 13603 13030 13655 13082
rect 13667 13030 13719 13082
rect 6368 12724 6420 12776
rect 5540 12588 5592 12640
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 10976 12486 11028 12538
rect 11040 12486 11092 12538
rect 11104 12486 11156 12538
rect 11168 12486 11220 12538
rect 9588 12316 9640 12368
rect 15660 12359 15712 12368
rect 15660 12325 15669 12359
rect 15669 12325 15703 12359
rect 15703 12325 15712 12359
rect 15660 12316 15712 12325
rect 6920 12248 6972 12300
rect 7380 12248 7432 12300
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 7472 12044 7524 12096
rect 3480 11942 3532 11994
rect 3544 11942 3596 11994
rect 3608 11942 3660 11994
rect 3672 11942 3724 11994
rect 8478 11942 8530 11994
rect 8542 11942 8594 11994
rect 8606 11942 8658 11994
rect 8670 11942 8722 11994
rect 13475 11942 13527 11994
rect 13539 11942 13591 11994
rect 13603 11942 13655 11994
rect 13667 11942 13719 11994
rect 9588 11840 9640 11892
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 7104 11568 7156 11620
rect 7748 11568 7800 11620
rect 12532 11636 12584 11688
rect 9312 11568 9364 11620
rect 3240 11500 3292 11552
rect 6368 11500 6420 11552
rect 8116 11500 8168 11552
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 10976 11398 11028 11450
rect 11040 11398 11092 11450
rect 11104 11398 11156 11450
rect 11168 11398 11220 11450
rect 5540 11296 5592 11348
rect 7104 11160 7156 11212
rect 7288 11160 7340 11212
rect 8576 11296 8628 11348
rect 9036 11296 9088 11348
rect 7564 11228 7616 11280
rect 7748 11228 7800 11280
rect 8116 11160 8168 11212
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 7012 11024 7064 11076
rect 7288 11067 7340 11076
rect 7288 11033 7297 11067
rect 7297 11033 7331 11067
rect 7331 11033 7340 11067
rect 7288 11024 7340 11033
rect 7564 10956 7616 11008
rect 8300 10956 8352 11008
rect 8944 10956 8996 11008
rect 15200 10956 15252 11008
rect 3480 10854 3532 10906
rect 3544 10854 3596 10906
rect 3608 10854 3660 10906
rect 3672 10854 3724 10906
rect 8478 10854 8530 10906
rect 8542 10854 8594 10906
rect 8606 10854 8658 10906
rect 8670 10854 8722 10906
rect 13475 10854 13527 10906
rect 13539 10854 13591 10906
rect 13603 10854 13655 10906
rect 13667 10854 13719 10906
rect 3240 10616 3292 10668
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 7656 10616 7708 10668
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 10876 10752 10928 10804
rect 3148 10548 3200 10600
rect 8944 10548 8996 10600
rect 8116 10480 8168 10532
rect 8392 10480 8444 10532
rect 8300 10412 8352 10464
rect 9588 10480 9640 10532
rect 10048 10548 10100 10600
rect 10416 10591 10468 10600
rect 10416 10557 10425 10591
rect 10425 10557 10459 10591
rect 10459 10557 10468 10591
rect 10416 10548 10468 10557
rect 10876 10548 10928 10600
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 9404 10412 9456 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 10508 10412 10560 10464
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 10976 10310 11028 10362
rect 11040 10310 11092 10362
rect 11104 10310 11156 10362
rect 11168 10310 11220 10362
rect 9128 10208 9180 10260
rect 10232 10208 10284 10260
rect 1584 10183 1636 10192
rect 1584 10149 1593 10183
rect 1593 10149 1627 10183
rect 1627 10149 1636 10183
rect 1584 10140 1636 10149
rect 3148 10140 3200 10192
rect 8300 10140 8352 10192
rect 8852 10140 8904 10192
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 9036 10072 9088 10124
rect 9588 10072 9640 10124
rect 7104 10004 7156 10056
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 10600 9936 10652 9988
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 7564 9868 7616 9920
rect 9312 9868 9364 9920
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 3480 9766 3532 9818
rect 3544 9766 3596 9818
rect 3608 9766 3660 9818
rect 3672 9766 3724 9818
rect 8478 9766 8530 9818
rect 8542 9766 8594 9818
rect 8606 9766 8658 9818
rect 8670 9766 8722 9818
rect 13475 9766 13527 9818
rect 13539 9766 13591 9818
rect 13603 9766 13655 9818
rect 13667 9766 13719 9818
rect 7104 9707 7156 9716
rect 7104 9673 7113 9707
rect 7113 9673 7147 9707
rect 7147 9673 7156 9707
rect 7104 9664 7156 9673
rect 7380 9528 7432 9580
rect 8300 9528 8352 9580
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 9588 9460 9640 9512
rect 9956 9392 10008 9444
rect 8300 9367 8352 9376
rect 8300 9333 8309 9367
rect 8309 9333 8343 9367
rect 8343 9333 8352 9367
rect 8300 9324 8352 9333
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 10976 9222 11028 9274
rect 11040 9222 11092 9274
rect 11104 9222 11156 9274
rect 11168 9222 11220 9274
rect 7288 9120 7340 9172
rect 8300 9052 8352 9104
rect 12532 9095 12584 9104
rect 12532 9061 12541 9095
rect 12541 9061 12575 9095
rect 12575 9061 12584 9095
rect 12532 9052 12584 9061
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 7564 8916 7616 8968
rect 4160 8780 4212 8832
rect 13268 8780 13320 8832
rect 3480 8678 3532 8730
rect 3544 8678 3596 8730
rect 3608 8678 3660 8730
rect 3672 8678 3724 8730
rect 8478 8678 8530 8730
rect 8542 8678 8594 8730
rect 8606 8678 8658 8730
rect 8670 8678 8722 8730
rect 13475 8678 13527 8730
rect 13539 8678 13591 8730
rect 13603 8678 13655 8730
rect 13667 8678 13719 8730
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 10976 8134 11028 8186
rect 11040 8134 11092 8186
rect 11104 8134 11156 8186
rect 11168 8134 11220 8186
rect 3480 7590 3532 7642
rect 3544 7590 3596 7642
rect 3608 7590 3660 7642
rect 3672 7590 3724 7642
rect 8478 7590 8530 7642
rect 8542 7590 8594 7642
rect 8606 7590 8658 7642
rect 8670 7590 8722 7642
rect 13475 7590 13527 7642
rect 13539 7590 13591 7642
rect 13603 7590 13655 7642
rect 13667 7590 13719 7642
rect 5448 7352 5500 7404
rect 9036 7352 9088 7404
rect 4160 7284 4212 7336
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 10976 7046 11028 7098
rect 11040 7046 11092 7098
rect 11104 7046 11156 7098
rect 11168 7046 11220 7098
rect 3480 6502 3532 6554
rect 3544 6502 3596 6554
rect 3608 6502 3660 6554
rect 3672 6502 3724 6554
rect 8478 6502 8530 6554
rect 8542 6502 8594 6554
rect 8606 6502 8658 6554
rect 8670 6502 8722 6554
rect 13475 6502 13527 6554
rect 13539 6502 13591 6554
rect 13603 6502 13655 6554
rect 13667 6502 13719 6554
rect 6552 6060 6604 6112
rect 9588 6060 9640 6112
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 10976 5958 11028 6010
rect 11040 5958 11092 6010
rect 11104 5958 11156 6010
rect 11168 5958 11220 6010
rect 3884 5856 3936 5908
rect 6644 5720 6696 5772
rect 7840 5856 7892 5908
rect 9128 5856 9180 5908
rect 7932 5788 7984 5840
rect 10048 5788 10100 5840
rect 14556 5856 14608 5908
rect 15108 5788 15160 5840
rect 11796 5763 11848 5772
rect 7012 5652 7064 5704
rect 11796 5729 11805 5763
rect 11805 5729 11839 5763
rect 11839 5729 11848 5763
rect 11796 5720 11848 5729
rect 13268 5652 13320 5704
rect 4620 5584 4672 5636
rect 8208 5584 8260 5636
rect 14004 5584 14056 5636
rect 2780 5516 2832 5568
rect 3976 5516 4028 5568
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 9312 5516 9364 5568
rect 10140 5516 10192 5568
rect 10876 5516 10928 5568
rect 3480 5414 3532 5466
rect 3544 5414 3596 5466
rect 3608 5414 3660 5466
rect 3672 5414 3724 5466
rect 8478 5414 8530 5466
rect 8542 5414 8594 5466
rect 8606 5414 8658 5466
rect 8670 5414 8722 5466
rect 13475 5414 13527 5466
rect 13539 5414 13591 5466
rect 13603 5414 13655 5466
rect 13667 5414 13719 5466
rect 3240 5312 3292 5364
rect 8024 5312 8076 5364
rect 2688 5244 2740 5296
rect 4068 5176 4120 5228
rect 7932 5244 7984 5296
rect 9220 5312 9272 5364
rect 9588 5312 9640 5364
rect 10324 5312 10376 5364
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 11980 5312 12032 5364
rect 12624 5355 12676 5364
rect 12624 5321 12633 5355
rect 12633 5321 12667 5355
rect 12667 5321 12676 5355
rect 12624 5312 12676 5321
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 8300 5244 8352 5296
rect 8760 5244 8812 5296
rect 9036 5244 9088 5296
rect 9496 5244 9548 5296
rect 9864 5244 9916 5296
rect 9956 5244 10008 5296
rect 10600 5244 10652 5296
rect 3332 5108 3384 5160
rect 4896 5108 4948 5160
rect 5080 5108 5132 5160
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 6276 5151 6328 5160
rect 6276 5117 6285 5151
rect 6285 5117 6319 5151
rect 6319 5117 6328 5151
rect 6276 5108 6328 5117
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7564 5108 7616 5160
rect 7748 5108 7800 5160
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 8852 5176 8904 5228
rect 8944 5176 8996 5228
rect 11796 5176 11848 5228
rect 9772 5151 9824 5160
rect 1952 5040 2004 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 8944 5040 8996 5092
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 10232 5151 10284 5160
rect 10232 5117 10241 5151
rect 10241 5117 10275 5151
rect 10275 5117 10284 5151
rect 10232 5108 10284 5117
rect 10784 5108 10836 5160
rect 15292 5244 15344 5296
rect 9404 5040 9456 5092
rect 6276 4972 6328 5024
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 9036 4972 9088 5024
rect 11152 5040 11204 5092
rect 9680 4972 9732 5024
rect 14832 5176 14884 5228
rect 12348 5151 12400 5160
rect 12348 5117 12357 5151
rect 12357 5117 12391 5151
rect 12391 5117 12400 5151
rect 12348 5108 12400 5117
rect 13084 5151 13136 5160
rect 12716 5040 12768 5092
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 14924 5108 14976 5160
rect 15476 5040 15528 5092
rect 12164 4972 12216 5024
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 10976 4870 11028 4922
rect 11040 4870 11092 4922
rect 11104 4870 11156 4922
rect 11168 4870 11220 4922
rect 4896 4768 4948 4820
rect 6920 4768 6972 4820
rect 7748 4768 7800 4820
rect 9036 4768 9088 4820
rect 9588 4768 9640 4820
rect 9956 4768 10008 4820
rect 12348 4768 12400 4820
rect 14188 4768 14240 4820
rect 4528 4700 4580 4752
rect 7472 4700 7524 4752
rect 7932 4700 7984 4752
rect 5356 4632 5408 4684
rect 8116 4632 8168 4684
rect 10416 4700 10468 4752
rect 10784 4700 10836 4752
rect 14832 4700 14884 4752
rect 8944 4564 8996 4616
rect 9772 4632 9824 4684
rect 13820 4632 13872 4684
rect 9588 4564 9640 4616
rect 10968 4564 11020 4616
rect 11336 4564 11388 4616
rect 11888 4564 11940 4616
rect 12716 4564 12768 4616
rect 15108 4564 15160 4616
rect 12072 4496 12124 4548
rect 5816 4428 5868 4480
rect 9680 4428 9732 4480
rect 10232 4428 10284 4480
rect 14556 4428 14608 4480
rect 3480 4326 3532 4378
rect 3544 4326 3596 4378
rect 3608 4326 3660 4378
rect 3672 4326 3724 4378
rect 8478 4326 8530 4378
rect 8542 4326 8594 4378
rect 8606 4326 8658 4378
rect 8670 4326 8722 4378
rect 13475 4326 13527 4378
rect 13539 4326 13591 4378
rect 13603 4326 13655 4378
rect 13667 4326 13719 4378
rect 9220 4224 9272 4276
rect 13268 4224 13320 4276
rect 7564 4156 7616 4208
rect 7196 4088 7248 4140
rect 9404 4088 9456 4140
rect 11428 4156 11480 4208
rect 12164 4156 12216 4208
rect 11520 4088 11572 4140
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 10976 3782 11028 3834
rect 11040 3782 11092 3834
rect 11104 3782 11156 3834
rect 11168 3782 11220 3834
rect 15200 3680 15252 3732
rect 15476 3723 15528 3732
rect 15476 3689 15485 3723
rect 15485 3689 15519 3723
rect 15519 3689 15528 3723
rect 15476 3680 15528 3689
rect 16948 3544 17000 3596
rect 15384 3383 15436 3392
rect 15384 3349 15393 3383
rect 15393 3349 15427 3383
rect 15427 3349 15436 3383
rect 15384 3340 15436 3349
rect 3480 3238 3532 3290
rect 3544 3238 3596 3290
rect 3608 3238 3660 3290
rect 3672 3238 3724 3290
rect 8478 3238 8530 3290
rect 8542 3238 8594 3290
rect 8606 3238 8658 3290
rect 8670 3238 8722 3290
rect 13475 3238 13527 3290
rect 13539 3238 13591 3290
rect 13603 3238 13655 3290
rect 13667 3238 13719 3290
rect 1400 3179 1452 3188
rect 1400 3145 1409 3179
rect 1409 3145 1443 3179
rect 1443 3145 1452 3179
rect 1400 3136 1452 3145
rect 15292 3136 15344 3188
rect 5632 3068 5684 3120
rect 9220 3068 9272 3120
rect 14280 3068 14332 3120
rect 16488 3068 16540 3120
rect 5540 3000 5592 3052
rect 8208 3000 8260 3052
rect 10324 3000 10376 3052
rect 3148 2932 3200 2984
rect 5632 2932 5684 2984
rect 7748 2932 7800 2984
rect 9128 2932 9180 2984
rect 4068 2907 4120 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 4068 2873 4077 2907
rect 4077 2873 4111 2907
rect 4111 2873 4120 2907
rect 4068 2864 4120 2873
rect 8852 2864 8904 2916
rect 13912 2864 13964 2916
rect 15200 2932 15252 2984
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 15568 2932 15620 2984
rect 8300 2796 8352 2848
rect 9588 2796 9640 2848
rect 10876 2796 10928 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 12624 2796 12676 2848
rect 13360 2796 13412 2848
rect 14372 2839 14424 2848
rect 14372 2805 14381 2839
rect 14381 2805 14415 2839
rect 14415 2805 14424 2839
rect 14372 2796 14424 2805
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 16028 2864 16080 2916
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 10976 2694 11028 2746
rect 11040 2694 11092 2746
rect 11104 2694 11156 2746
rect 11168 2694 11220 2746
rect 2780 2592 2832 2644
rect 1492 2524 1544 2576
rect 4436 2592 4488 2644
rect 2044 2456 2096 2508
rect 3884 2524 3936 2576
rect 4620 2567 4672 2576
rect 4620 2533 4629 2567
rect 4629 2533 4663 2567
rect 4663 2533 4672 2567
rect 4620 2524 4672 2533
rect 5540 2567 5592 2576
rect 5540 2533 5549 2567
rect 5549 2533 5583 2567
rect 5583 2533 5592 2567
rect 5540 2524 5592 2533
rect 5632 2524 5684 2576
rect 2964 2456 3016 2508
rect 3332 2456 3384 2508
rect 3976 2456 4028 2508
rect 5080 2499 5132 2508
rect 5080 2465 5089 2499
rect 5089 2465 5123 2499
rect 5123 2465 5132 2499
rect 5080 2456 5132 2465
rect 7748 2592 7800 2644
rect 7840 2592 7892 2644
rect 8944 2592 8996 2644
rect 9220 2635 9272 2644
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 9404 2592 9456 2644
rect 9956 2592 10008 2644
rect 10232 2592 10284 2644
rect 10692 2592 10744 2644
rect 10784 2592 10836 2644
rect 11520 2592 11572 2644
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 7380 2524 7432 2576
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 1032 2388 1084 2440
rect 2780 2388 2832 2440
rect 204 2320 256 2372
rect 2320 2320 2372 2372
rect 3332 2320 3384 2372
rect 5172 2388 5224 2440
rect 6644 2388 6696 2440
rect 7012 2388 7064 2440
rect 4436 2363 4488 2372
rect 4436 2329 4445 2363
rect 4445 2329 4479 2363
rect 4479 2329 4488 2363
rect 4436 2320 4488 2329
rect 4896 2363 4948 2372
rect 4896 2329 4905 2363
rect 4905 2329 4939 2363
rect 4939 2329 4948 2363
rect 4896 2320 4948 2329
rect 5356 2363 5408 2372
rect 5356 2329 5365 2363
rect 5365 2329 5399 2363
rect 5399 2329 5408 2363
rect 5356 2320 5408 2329
rect 5724 2363 5776 2372
rect 5724 2329 5733 2363
rect 5733 2329 5767 2363
rect 5767 2329 5776 2363
rect 5724 2320 5776 2329
rect 6184 2320 6236 2372
rect 7472 2320 7524 2372
rect 7932 2320 7984 2372
rect 572 2252 624 2304
rect 1952 2252 2004 2304
rect 3056 2252 3108 2304
rect 6276 2252 6328 2304
rect 8300 2320 8352 2372
rect 8760 2456 8812 2508
rect 9220 2456 9272 2508
rect 9680 2456 9732 2508
rect 10048 2456 10100 2508
rect 9036 2388 9088 2440
rect 10508 2456 10560 2508
rect 12900 2592 12952 2644
rect 13268 2592 13320 2644
rect 13820 2592 13872 2644
rect 14188 2635 14240 2644
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 14556 2635 14608 2644
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 15108 2635 15160 2644
rect 15108 2601 15117 2635
rect 15117 2601 15151 2635
rect 15151 2601 15160 2635
rect 15108 2592 15160 2601
rect 15292 2592 15344 2644
rect 11060 2499 11112 2508
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 11060 2456 11112 2465
rect 11336 2456 11388 2508
rect 11796 2456 11848 2508
rect 12164 2456 12216 2508
rect 12256 2456 12308 2508
rect 12624 2456 12676 2508
rect 13084 2456 13136 2508
rect 13360 2456 13412 2508
rect 13912 2456 13964 2508
rect 14280 2456 14332 2508
rect 14464 2456 14516 2508
rect 14832 2456 14884 2508
rect 15200 2456 15252 2508
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 12072 2320 12124 2372
rect 12440 2320 12492 2372
rect 10232 2252 10284 2304
rect 10416 2252 10468 2304
rect 11336 2252 11388 2304
rect 12256 2252 12308 2304
rect 12992 2252 13044 2304
rect 3480 2150 3532 2202
rect 3544 2150 3596 2202
rect 3608 2150 3660 2202
rect 3672 2150 3724 2202
rect 8478 2150 8530 2202
rect 8542 2150 8594 2202
rect 8606 2150 8658 2202
rect 8670 2150 8722 2202
rect 13475 2150 13527 2202
rect 13539 2150 13591 2202
rect 13603 2150 13655 2202
rect 13667 2150 13719 2202
rect 2044 2048 2096 2100
rect 4804 2048 4856 2100
rect 8944 2048 8996 2100
rect 11428 2048 11480 2100
rect 7104 1980 7156 2032
rect 10140 1980 10192 2032
rect 10324 1980 10376 2032
rect 12992 2048 13044 2100
rect 5080 1844 5132 1896
rect 9312 1844 9364 1896
rect 6736 1776 6788 1828
rect 10600 1776 10652 1828
rect 7656 1708 7708 1760
rect 10416 1708 10468 1760
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1858 19200 1914 20000
rect 2226 19200 2282 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3514 19200 3570 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4802 19200 4858 20000
rect 5170 19200 5226 20000
rect 5630 19200 5686 20000
rect 5998 19200 6054 20000
rect 6458 19200 6514 20000
rect 6826 19200 6882 20000
rect 7286 19200 7342 20000
rect 7746 19200 7802 20000
rect 8114 19200 8170 20000
rect 8574 19200 8630 20000
rect 8942 19200 8998 20000
rect 9402 19200 9458 20000
rect 9770 19200 9826 20000
rect 10230 19200 10286 20000
rect 10690 19200 10746 20000
rect 11058 19200 11114 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12346 19200 12402 20000
rect 12714 19200 12770 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 14002 19200 14058 20000
rect 14462 19200 14518 20000
rect 14830 19200 14886 20000
rect 15290 19200 15346 20000
rect 15658 19200 15714 20000
rect 16118 19200 16174 20000
rect 16486 19200 16542 20000
rect 16946 19200 17002 20000
rect 216 16658 244 19200
rect 584 17270 612 19200
rect 1044 17338 1072 19200
rect 1032 17332 1084 17338
rect 1032 17274 1084 17280
rect 572 17264 624 17270
rect 572 17206 624 17212
rect 1412 17134 1440 19200
rect 1674 18320 1730 18329
rect 1674 18255 1730 18264
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1584 17060 1636 17066
rect 1584 17002 1636 17008
rect 204 16652 256 16658
rect 204 16594 256 16600
rect 1596 15162 1624 17002
rect 1688 16658 1716 18255
rect 1872 17202 1900 19200
rect 2240 17338 2268 19200
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2700 17252 2728 19200
rect 3068 17338 3096 19200
rect 3528 17626 3556 19200
rect 3988 17626 4016 19200
rect 3528 17598 3832 17626
rect 3988 17598 4200 17626
rect 3454 17436 3750 17456
rect 3510 17434 3534 17436
rect 3590 17434 3614 17436
rect 3670 17434 3694 17436
rect 3532 17382 3534 17434
rect 3596 17382 3608 17434
rect 3670 17382 3672 17434
rect 3510 17380 3534 17382
rect 3590 17380 3614 17382
rect 3670 17380 3694 17382
rect 3454 17360 3750 17380
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3804 17270 3832 17598
rect 4172 17542 4200 17598
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4356 17338 4384 19200
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4816 17270 4844 19200
rect 5184 17270 5212 19200
rect 5644 17270 5672 19200
rect 6012 17270 6040 19200
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 2780 17264 2832 17270
rect 2700 17224 2780 17252
rect 2780 17206 2832 17212
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1398 15056 1454 15065
rect 1398 14991 1400 15000
rect 1452 14991 1454 15000
rect 1400 14962 1452 14968
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1400 11688 1452 11694
rect 1398 11656 1400 11665
rect 1452 11656 1454 11665
rect 1398 11591 1454 11600
rect 1584 10192 1636 10198
rect 1584 10134 1636 10140
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1398 8392 1454 8401
rect 1398 8327 1400 8336
rect 1452 8327 1454 8336
rect 1400 8298 1452 8304
rect 1504 6914 1532 9998
rect 1596 8430 1624 10134
rect 1780 10062 1808 14826
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1412 6886 1532 6914
rect 1412 3194 1440 6886
rect 1964 5098 1992 17002
rect 2700 5302 2728 17002
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2792 13394 2820 16730
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 10606 3188 13126
rect 3252 12434 3280 17002
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 3454 16348 3750 16368
rect 3510 16346 3534 16348
rect 3590 16346 3614 16348
rect 3670 16346 3694 16348
rect 3532 16294 3534 16346
rect 3596 16294 3608 16346
rect 3670 16294 3672 16346
rect 3510 16292 3534 16294
rect 3590 16292 3614 16294
rect 3670 16292 3694 16294
rect 3454 16272 3750 16292
rect 3454 15260 3750 15280
rect 3510 15258 3534 15260
rect 3590 15258 3614 15260
rect 3670 15258 3694 15260
rect 3532 15206 3534 15258
rect 3596 15206 3608 15258
rect 3670 15206 3672 15258
rect 3510 15204 3534 15206
rect 3590 15204 3614 15206
rect 3670 15204 3694 15206
rect 3454 15184 3750 15204
rect 3454 14172 3750 14192
rect 3510 14170 3534 14172
rect 3590 14170 3614 14172
rect 3670 14170 3694 14172
rect 3532 14118 3534 14170
rect 3596 14118 3608 14170
rect 3670 14118 3672 14170
rect 3510 14116 3534 14118
rect 3590 14116 3614 14118
rect 3670 14116 3694 14118
rect 3454 14096 3750 14116
rect 3988 13462 4016 16662
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3454 13084 3750 13104
rect 3510 13082 3534 13084
rect 3590 13082 3614 13084
rect 3670 13082 3694 13084
rect 3532 13030 3534 13082
rect 3596 13030 3608 13082
rect 3670 13030 3672 13082
rect 3510 13028 3534 13030
rect 3590 13028 3614 13030
rect 3670 13028 3694 13030
rect 3454 13008 3750 13028
rect 3252 12406 3372 12434
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 10674 3280 11494
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 10198 3188 10542
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3344 7834 3372 12406
rect 3454 11996 3750 12016
rect 3510 11994 3534 11996
rect 3590 11994 3614 11996
rect 3670 11994 3694 11996
rect 3532 11942 3534 11994
rect 3596 11942 3608 11994
rect 3670 11942 3672 11994
rect 3510 11940 3534 11942
rect 3590 11940 3614 11942
rect 3670 11940 3694 11942
rect 3454 11920 3750 11940
rect 3454 10908 3750 10928
rect 3510 10906 3534 10908
rect 3590 10906 3614 10908
rect 3670 10906 3694 10908
rect 3532 10854 3534 10906
rect 3596 10854 3608 10906
rect 3670 10854 3672 10906
rect 3510 10852 3534 10854
rect 3590 10852 3614 10854
rect 3670 10852 3694 10854
rect 3454 10832 3750 10852
rect 3454 9820 3750 9840
rect 3510 9818 3534 9820
rect 3590 9818 3614 9820
rect 3670 9818 3694 9820
rect 3532 9766 3534 9818
rect 3596 9766 3608 9818
rect 3670 9766 3672 9818
rect 3510 9764 3534 9766
rect 3590 9764 3614 9766
rect 3670 9764 3694 9766
rect 3454 9744 3750 9764
rect 3454 8732 3750 8752
rect 3510 8730 3534 8732
rect 3590 8730 3614 8732
rect 3670 8730 3694 8732
rect 3532 8678 3534 8730
rect 3596 8678 3608 8730
rect 3670 8678 3672 8730
rect 3510 8676 3534 8678
rect 3590 8676 3614 8678
rect 3670 8676 3694 8678
rect 3454 8656 3750 8676
rect 3252 7806 3372 7834
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1492 5024 1544 5030
rect 1490 4992 1492 5001
rect 1544 4992 1546 5001
rect 1490 4927 1546 4936
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1492 2576 1544 2582
rect 1492 2518 1544 2524
rect 1032 2440 1084 2446
rect 1032 2382 1084 2388
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 800 244 2314
rect 572 2304 624 2310
rect 572 2246 624 2252
rect 584 800 612 2246
rect 1044 800 1072 2382
rect 1504 800 1532 2518
rect 1688 1737 1716 2790
rect 2792 2650 2820 5510
rect 3252 5370 3280 7806
rect 3454 7644 3750 7664
rect 3510 7642 3534 7644
rect 3590 7642 3614 7644
rect 3670 7642 3694 7644
rect 3532 7590 3534 7642
rect 3596 7590 3608 7642
rect 3670 7590 3672 7642
rect 3510 7588 3534 7590
rect 3590 7588 3614 7590
rect 3670 7588 3694 7590
rect 3454 7568 3750 7588
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3344 5166 3372 7142
rect 3454 6556 3750 6576
rect 3510 6554 3534 6556
rect 3590 6554 3614 6556
rect 3670 6554 3694 6556
rect 3532 6502 3534 6554
rect 3596 6502 3608 6554
rect 3670 6502 3672 6554
rect 3510 6500 3534 6502
rect 3590 6500 3614 6502
rect 3670 6500 3694 6502
rect 3454 6480 3750 6500
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3454 5468 3750 5488
rect 3510 5466 3534 5468
rect 3590 5466 3614 5468
rect 3670 5466 3694 5468
rect 3532 5414 3534 5466
rect 3596 5414 3608 5466
rect 3670 5414 3672 5466
rect 3510 5412 3534 5414
rect 3590 5412 3614 5414
rect 3670 5412 3694 5414
rect 3454 5392 3750 5412
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3454 4380 3750 4400
rect 3510 4378 3534 4380
rect 3590 4378 3614 4380
rect 3670 4378 3694 4380
rect 3532 4326 3534 4378
rect 3596 4326 3608 4378
rect 3670 4326 3672 4378
rect 3510 4324 3534 4326
rect 3590 4324 3614 4326
rect 3670 4324 3694 4326
rect 3454 4304 3750 4324
rect 3454 3292 3750 3312
rect 3510 3290 3534 3292
rect 3590 3290 3614 3292
rect 3670 3290 3694 3292
rect 3532 3238 3534 3290
rect 3596 3238 3608 3290
rect 3670 3238 3672 3290
rect 3510 3236 3534 3238
rect 3590 3236 3614 3238
rect 3670 3236 3694 3238
rect 3454 3216 3750 3236
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2964 2508 3016 2514
rect 3016 2468 3096 2496
rect 2964 2450 3016 2456
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1674 1728 1730 1737
rect 1674 1663 1730 1672
rect 1964 1170 1992 2246
rect 2056 2106 2084 2450
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 1872 1142 1992 1170
rect 1872 800 1900 1142
rect 2332 800 2360 2314
rect 2792 800 2820 2382
rect 3068 2310 3096 2468
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3160 800 3188 2926
rect 3700 2848 3752 2854
rect 3752 2808 3832 2836
rect 3700 2790 3752 2796
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3344 2378 3372 2450
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3454 2204 3750 2224
rect 3510 2202 3534 2204
rect 3590 2202 3614 2204
rect 3670 2202 3694 2204
rect 3532 2150 3534 2202
rect 3596 2150 3608 2202
rect 3670 2150 3672 2202
rect 3510 2148 3534 2150
rect 3590 2148 3614 2150
rect 3670 2148 3694 2150
rect 3454 2128 3750 2148
rect 3804 898 3832 2808
rect 3896 2582 3924 5850
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 3988 2514 4016 5510
rect 4080 5234 4108 17002
rect 4448 12434 4476 17002
rect 4540 15162 4568 17070
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 5000 15094 5028 17002
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4448 12406 4568 12434
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 7342 4200 8774
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 3620 870 3832 898
rect 3620 800 3648 870
rect 4080 800 4108 2858
rect 4448 2650 4476 4966
rect 4540 4758 4568 12406
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4632 2582 4660 5578
rect 5092 5166 5120 17138
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 15162 5304 16934
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5368 12434 5396 17002
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 12646 5580 13330
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5368 12406 5488 12434
rect 5460 7410 5488 12406
rect 5552 11354 5580 12582
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4448 800 4476 2314
rect 4816 2106 4844 4966
rect 4908 4826 4936 5102
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 4908 800 4936 2314
rect 5092 1902 5120 2450
rect 5184 2446 5212 4966
rect 5368 4690 5396 5102
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5644 3126 5672 5102
rect 5828 4486 5856 17002
rect 5953 16892 6249 16912
rect 6009 16890 6033 16892
rect 6089 16890 6113 16892
rect 6169 16890 6193 16892
rect 6031 16838 6033 16890
rect 6095 16838 6107 16890
rect 6169 16838 6171 16890
rect 6009 16836 6033 16838
rect 6089 16836 6113 16838
rect 6169 16836 6193 16838
rect 5953 16816 6249 16836
rect 5953 15804 6249 15824
rect 6009 15802 6033 15804
rect 6089 15802 6113 15804
rect 6169 15802 6193 15804
rect 6031 15750 6033 15802
rect 6095 15750 6107 15802
rect 6169 15750 6171 15802
rect 6009 15748 6033 15750
rect 6089 15748 6113 15750
rect 6169 15748 6193 15750
rect 5953 15728 6249 15748
rect 5953 14716 6249 14736
rect 6009 14714 6033 14716
rect 6089 14714 6113 14716
rect 6169 14714 6193 14716
rect 6031 14662 6033 14714
rect 6095 14662 6107 14714
rect 6169 14662 6171 14714
rect 6009 14660 6033 14662
rect 6089 14660 6113 14662
rect 6169 14660 6193 14662
rect 5953 14640 6249 14660
rect 5953 13628 6249 13648
rect 6009 13626 6033 13628
rect 6089 13626 6113 13628
rect 6169 13626 6193 13628
rect 6031 13574 6033 13626
rect 6095 13574 6107 13626
rect 6169 13574 6171 13626
rect 6009 13572 6033 13574
rect 6089 13572 6113 13574
rect 6169 13572 6193 13574
rect 5953 13552 6249 13572
rect 5953 12540 6249 12560
rect 6009 12538 6033 12540
rect 6089 12538 6113 12540
rect 6169 12538 6193 12540
rect 6031 12486 6033 12538
rect 6095 12486 6107 12538
rect 6169 12486 6171 12538
rect 6009 12484 6033 12486
rect 6089 12484 6113 12486
rect 6169 12484 6193 12486
rect 5953 12464 6249 12484
rect 5953 11452 6249 11472
rect 6009 11450 6033 11452
rect 6089 11450 6113 11452
rect 6169 11450 6193 11452
rect 6031 11398 6033 11450
rect 6095 11398 6107 11450
rect 6169 11398 6171 11450
rect 6009 11396 6033 11398
rect 6089 11396 6113 11398
rect 6169 11396 6193 11398
rect 5953 11376 6249 11396
rect 5953 10364 6249 10384
rect 6009 10362 6033 10364
rect 6089 10362 6113 10364
rect 6169 10362 6193 10364
rect 6031 10310 6033 10362
rect 6095 10310 6107 10362
rect 6169 10310 6171 10362
rect 6009 10308 6033 10310
rect 6089 10308 6113 10310
rect 6169 10308 6193 10310
rect 5953 10288 6249 10308
rect 5953 9276 6249 9296
rect 6009 9274 6033 9276
rect 6089 9274 6113 9276
rect 6169 9274 6193 9276
rect 6031 9222 6033 9274
rect 6095 9222 6107 9274
rect 6169 9222 6171 9274
rect 6009 9220 6033 9222
rect 6089 9220 6113 9222
rect 6169 9220 6193 9222
rect 5953 9200 6249 9220
rect 5953 8188 6249 8208
rect 6009 8186 6033 8188
rect 6089 8186 6113 8188
rect 6169 8186 6193 8188
rect 6031 8134 6033 8186
rect 6095 8134 6107 8186
rect 6169 8134 6171 8186
rect 6009 8132 6033 8134
rect 6089 8132 6113 8134
rect 6169 8132 6193 8134
rect 5953 8112 6249 8132
rect 5953 7100 6249 7120
rect 6009 7098 6033 7100
rect 6089 7098 6113 7100
rect 6169 7098 6193 7100
rect 6031 7046 6033 7098
rect 6095 7046 6107 7098
rect 6169 7046 6171 7098
rect 6009 7044 6033 7046
rect 6089 7044 6113 7046
rect 6169 7044 6193 7046
rect 5953 7024 6249 7044
rect 5953 6012 6249 6032
rect 6009 6010 6033 6012
rect 6089 6010 6113 6012
rect 6169 6010 6193 6012
rect 6031 5958 6033 6010
rect 6095 5958 6107 6010
rect 6169 5958 6171 6010
rect 6009 5956 6033 5958
rect 6089 5956 6113 5958
rect 6169 5956 6193 5958
rect 5953 5936 6249 5956
rect 6288 5166 6316 17818
rect 6472 17270 6500 19200
rect 6840 17898 6868 19200
rect 6840 17870 6960 17898
rect 6932 17270 6960 17870
rect 7300 17270 7328 19200
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 7288 17264 7340 17270
rect 7288 17206 7340 17212
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6380 11558 6408 12718
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6564 6118 6592 17002
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6656 5778 6684 16730
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6748 5273 6776 17002
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6734 5264 6790 5273
rect 6734 5199 6790 5208
rect 6000 5160 6052 5166
rect 5998 5128 6000 5137
rect 6276 5160 6328 5166
rect 6052 5128 6054 5137
rect 6276 5102 6328 5108
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 5998 5063 6054 5072
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5953 4924 6249 4944
rect 6009 4922 6033 4924
rect 6089 4922 6113 4924
rect 6169 4922 6193 4924
rect 6031 4870 6033 4922
rect 6095 4870 6107 4922
rect 6169 4870 6171 4922
rect 6009 4868 6033 4870
rect 6089 4868 6113 4870
rect 6169 4868 6193 4870
rect 5953 4848 6249 4868
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5953 3836 6249 3856
rect 6009 3834 6033 3836
rect 6089 3834 6113 3836
rect 6169 3834 6193 3836
rect 6031 3782 6033 3834
rect 6095 3782 6107 3834
rect 6169 3782 6171 3834
rect 6009 3780 6033 3782
rect 6089 3780 6113 3782
rect 6169 3780 6193 3782
rect 5953 3760 6249 3780
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5552 2582 5580 2994
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2582 5672 2926
rect 5953 2748 6249 2768
rect 6009 2746 6033 2748
rect 6089 2746 6113 2748
rect 6169 2746 6193 2748
rect 6031 2694 6033 2746
rect 6095 2694 6107 2746
rect 6169 2694 6171 2746
rect 6009 2692 6033 2694
rect 6089 2692 6113 2694
rect 6169 2692 6193 2694
rect 5953 2672 6249 2692
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 5080 1896 5132 1902
rect 5080 1838 5132 1844
rect 5368 800 5396 2314
rect 5736 800 5764 2314
rect 6196 800 6224 2314
rect 6288 2310 6316 4966
rect 6840 4729 6868 5102
rect 6932 4826 6960 12242
rect 7024 12238 7052 13126
rect 7116 12434 7144 14826
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7116 12406 7236 12434
rect 7208 12238 7236 12406
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7024 11082 7052 12174
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7116 11218 7144 11562
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10674 7052 11018
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7116 10554 7144 11154
rect 7024 10526 7144 10554
rect 7024 5710 7052 10526
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7116 9722 7144 9998
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6826 4720 6882 4729
rect 6826 4655 6882 4664
rect 7208 4146 7236 12174
rect 7300 11218 7328 14758
rect 7392 12306 7420 17614
rect 7760 17270 7788 19200
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 14618 7512 17002
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 12434 7604 14826
rect 7576 12406 7696 12434
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7300 10010 7328 11018
rect 7300 9982 7420 10010
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7300 9178 7328 9862
rect 7392 9586 7420 9982
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7484 9518 7512 12038
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7576 11014 7604 11222
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7668 10674 7696 12406
rect 7760 11626 7788 16662
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7576 8974 7604 9862
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7392 2582 7420 5510
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4758 7512 4966
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7576 4214 7604 5102
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6656 800 6684 2382
rect 6748 1834 6776 2450
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6736 1828 6788 1834
rect 6736 1770 6788 1776
rect 7024 800 7052 2382
rect 7116 2038 7144 2450
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7104 2032 7156 2038
rect 7104 1974 7156 1980
rect 7484 800 7512 2314
rect 7668 1766 7696 10610
rect 7760 5794 7788 11222
rect 7852 5914 7880 17750
rect 8128 17270 8156 19200
rect 8588 18170 8616 19200
rect 8588 18142 8892 18170
rect 8300 17944 8352 17950
rect 8300 17886 8352 17892
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 7930 16688 7986 16697
rect 7930 16623 7986 16632
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7944 5846 7972 16623
rect 7932 5840 7984 5846
rect 7760 5766 7880 5794
rect 7932 5782 7984 5788
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7760 4826 7788 5102
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 2650 7788 2926
rect 7852 2650 7880 5766
rect 7930 5672 7986 5681
rect 7930 5607 7986 5616
rect 7944 5302 7972 5607
rect 8036 5370 8064 16934
rect 8128 16658 8156 17002
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11218 8156 11494
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8220 10554 8248 17546
rect 8312 17066 8340 17886
rect 8452 17436 8748 17456
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8530 17382 8532 17434
rect 8594 17382 8606 17434
rect 8668 17382 8670 17434
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8452 17360 8748 17380
rect 8864 17338 8892 18142
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8680 16969 8708 17070
rect 8852 16992 8904 16998
rect 8666 16960 8722 16969
rect 8852 16934 8904 16940
rect 8666 16895 8722 16904
rect 8864 16726 8892 16934
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 8956 16522 8984 19200
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8452 16348 8748 16368
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8530 16294 8532 16346
rect 8594 16294 8606 16346
rect 8668 16294 8670 16346
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8452 16272 8748 16292
rect 8452 15260 8748 15280
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8530 15206 8532 15258
rect 8594 15206 8606 15258
rect 8668 15206 8670 15258
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8452 15184 8748 15204
rect 8452 14172 8748 14192
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8530 14118 8532 14170
rect 8594 14118 8606 14170
rect 8668 14118 8670 14170
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8452 14096 8748 14116
rect 8452 13084 8748 13104
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8530 13030 8532 13082
rect 8594 13030 8606 13082
rect 8668 13030 8670 13082
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8452 13008 8748 13028
rect 8452 11996 8748 12016
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8530 11942 8532 11994
rect 8594 11942 8606 11994
rect 8668 11942 8670 11994
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8452 11920 8748 11940
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 11354 8616 11630
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8312 10690 8340 10950
rect 8452 10908 8748 10928
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8530 10854 8532 10906
rect 8594 10854 8606 10906
rect 8668 10854 8670 10906
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8452 10832 8748 10852
rect 8312 10662 8432 10690
rect 8128 10538 8248 10554
rect 8404 10538 8432 10662
rect 8956 10606 8984 10950
rect 9048 10674 9076 11290
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8116 10532 8248 10538
rect 8168 10526 8248 10532
rect 8392 10532 8444 10538
rect 8116 10474 8168 10480
rect 8392 10474 8444 10480
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7944 4758 7972 5102
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 8128 4690 8156 10474
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10198 8340 10406
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8404 10010 8432 10474
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8312 9982 8432 10010
rect 8312 9586 8340 9982
rect 8452 9820 8748 9840
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8530 9766 8532 9818
rect 8594 9766 8606 9818
rect 8668 9766 8670 9818
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8452 9744 8748 9764
rect 8864 9586 8892 10134
rect 9048 10130 9076 10610
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10266 9168 10406
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 9110 8340 9318
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8452 8732 8748 8752
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8530 8678 8532 8730
rect 8594 8678 8606 8730
rect 8668 8678 8670 8730
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8452 8656 8748 8676
rect 8452 7644 8748 7664
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8530 7590 8532 7642
rect 8594 7590 8606 7642
rect 8668 7590 8670 7642
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8452 7568 8748 7588
rect 9232 7562 9260 17682
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 17338 9352 17478
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9416 16454 9444 19200
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9324 9926 9352 11562
rect 9416 10470 9444 14758
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9508 9674 9536 17478
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9600 16794 9628 17274
rect 9784 17202 9812 19200
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9692 16250 9720 17070
rect 9784 16658 9812 17138
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 10060 16574 10088 17002
rect 10152 16726 10180 17070
rect 10244 17066 10272 19200
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10336 17270 10364 17614
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 9876 16546 10088 16574
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9600 12374 9628 13194
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9600 11898 9628 12310
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9600 10130 9628 10474
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 8864 7534 9260 7562
rect 9416 9646 9536 9674
rect 8452 6556 8748 6576
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8530 6502 8532 6554
rect 8594 6502 8606 6554
rect 8668 6502 8670 6554
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8452 6480 8748 6500
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8220 3058 8248 5578
rect 8452 5468 8748 5488
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8530 5414 8532 5466
rect 8594 5414 8606 5466
rect 8668 5414 8670 5466
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8452 5392 8748 5412
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8312 2854 8340 5238
rect 8772 4468 8800 5238
rect 8864 5234 8892 7534
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 5302 9076 7346
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 5098 8984 5170
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 4826 9076 4966
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8772 4440 8892 4468
rect 8452 4380 8748 4400
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8530 4326 8532 4378
rect 8594 4326 8606 4378
rect 8668 4326 8670 4378
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8452 4304 8748 4324
rect 8452 3292 8748 3312
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8530 3238 8532 3290
rect 8594 3238 8606 3290
rect 8668 3238 8670 3290
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8452 3216 8748 3236
rect 8864 2922 8892 4440
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8956 2650 8984 4558
rect 9140 2990 9168 5850
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 4282 9260 5306
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9232 2650 9260 3062
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 8300 2372 8352 2378
rect 8772 2360 8800 2450
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8772 2332 8984 2360
rect 8300 2314 8352 2320
rect 7656 1760 7708 1766
rect 7656 1702 7708 1708
rect 7944 800 7972 2314
rect 8312 800 8340 2314
rect 8452 2204 8748 2224
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8530 2150 8532 2202
rect 8594 2150 8606 2202
rect 8668 2150 8670 2202
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8452 2128 8748 2148
rect 8956 2106 8984 2332
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9048 1986 9076 2382
rect 8772 1958 9076 1986
rect 8772 800 8800 1958
rect 9232 800 9260 2450
rect 9324 1902 9352 5510
rect 9416 5098 9444 9646
rect 9600 9518 9628 9862
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9494 5672 9550 5681
rect 9494 5607 9550 5616
rect 9508 5302 9536 5607
rect 9600 5370 9628 6054
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9876 5302 9904 16546
rect 10152 16522 10180 16662
rect 10244 16522 10272 17002
rect 10322 16960 10378 16969
rect 10322 16895 10378 16904
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 12434 9996 14418
rect 9968 12406 10272 12434
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 10606 10088 11086
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 9450 9996 10406
rect 10244 10266 10272 12406
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10060 5846 10088 9998
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9864 5296 9916 5302
rect 9956 5296 10008 5302
rect 9864 5238 9916 5244
rect 9954 5264 9956 5273
rect 10008 5264 10010 5273
rect 9954 5199 10010 5208
rect 9772 5160 9824 5166
rect 9494 5128 9550 5137
rect 9404 5092 9456 5098
rect 9772 5102 9824 5108
rect 9494 5063 9550 5072
rect 9404 5034 9456 5040
rect 9508 4978 9536 5063
rect 9680 5024 9732 5030
rect 9508 4950 9628 4978
rect 9680 4966 9732 4972
rect 9600 4826 9628 4950
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9494 4720 9550 4729
rect 9550 4678 9628 4706
rect 9494 4655 9550 4664
rect 9600 4622 9628 4678
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9692 4486 9720 4966
rect 9784 4690 9812 5102
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9416 2650 9444 4082
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9600 2496 9628 2790
rect 9968 2650 9996 4762
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9680 2508 9732 2514
rect 9600 2468 9680 2496
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 9600 800 9628 2468
rect 9680 2450 9732 2456
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10060 800 10088 2450
rect 10152 2038 10180 5510
rect 10244 5250 10272 10202
rect 10336 5370 10364 16895
rect 10428 16794 10456 17070
rect 10520 16998 10548 17818
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10428 16454 10456 16730
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10244 5222 10364 5250
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4486 10272 5102
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10336 3058 10364 5222
rect 10428 4758 10456 10542
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10520 2774 10548 10406
rect 10612 9994 10640 17206
rect 10704 17082 10732 19200
rect 11072 17202 11100 19200
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11152 17128 11204 17134
rect 10704 17076 11152 17082
rect 10704 17070 11204 17076
rect 10704 17054 11192 17070
rect 10950 16892 11246 16912
rect 11006 16890 11030 16892
rect 11086 16890 11110 16892
rect 11166 16890 11190 16892
rect 11028 16838 11030 16890
rect 11092 16838 11104 16890
rect 11166 16838 11168 16890
rect 11006 16836 11030 16838
rect 11086 16836 11110 16838
rect 11166 16836 11190 16838
rect 10950 16816 11246 16836
rect 11348 16794 11376 17138
rect 11440 16998 11468 17546
rect 11532 17082 11560 19200
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11624 17338 11652 17478
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11612 17128 11664 17134
rect 11532 17076 11612 17082
rect 11532 17070 11664 17076
rect 11532 17054 11652 17070
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11532 16794 11560 17054
rect 11808 16998 11836 17750
rect 11900 17202 11928 19200
rect 11980 17944 12032 17950
rect 11980 17886 12032 17892
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11900 16794 11928 17138
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11612 16720 11664 16726
rect 10782 16688 10838 16697
rect 11612 16662 11664 16668
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 10782 16623 10784 16632
rect 10836 16623 10838 16632
rect 10784 16594 10836 16600
rect 10876 16584 10928 16590
rect 11624 16574 11652 16662
rect 11624 16546 11744 16574
rect 10876 16526 10928 16532
rect 10888 10810 10916 16526
rect 10950 15804 11246 15824
rect 11006 15802 11030 15804
rect 11086 15802 11110 15804
rect 11166 15802 11190 15804
rect 11028 15750 11030 15802
rect 11092 15750 11104 15802
rect 11166 15750 11168 15802
rect 11006 15748 11030 15750
rect 11086 15748 11110 15750
rect 11166 15748 11190 15750
rect 10950 15728 11246 15748
rect 10950 14716 11246 14736
rect 11006 14714 11030 14716
rect 11086 14714 11110 14716
rect 11166 14714 11190 14716
rect 11028 14662 11030 14714
rect 11092 14662 11104 14714
rect 11166 14662 11168 14714
rect 11006 14660 11030 14662
rect 11086 14660 11110 14662
rect 11166 14660 11190 14662
rect 10950 14640 11246 14660
rect 10950 13628 11246 13648
rect 11006 13626 11030 13628
rect 11086 13626 11110 13628
rect 11166 13626 11190 13628
rect 11028 13574 11030 13626
rect 11092 13574 11104 13626
rect 11166 13574 11168 13626
rect 11006 13572 11030 13574
rect 11086 13572 11110 13574
rect 11166 13572 11190 13574
rect 10950 13552 11246 13572
rect 10950 12540 11246 12560
rect 11006 12538 11030 12540
rect 11086 12538 11110 12540
rect 11166 12538 11190 12540
rect 11028 12486 11030 12538
rect 11092 12486 11104 12538
rect 11166 12486 11168 12538
rect 11006 12484 11030 12486
rect 11086 12484 11110 12486
rect 11166 12484 11190 12486
rect 10950 12464 11246 12484
rect 10950 11452 11246 11472
rect 11006 11450 11030 11452
rect 11086 11450 11110 11452
rect 11166 11450 11190 11452
rect 11028 11398 11030 11450
rect 11092 11398 11104 11450
rect 11166 11398 11168 11450
rect 11006 11396 11030 11398
rect 11086 11396 11110 11398
rect 11166 11396 11190 11398
rect 10950 11376 11246 11396
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10606 10916 10746
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10950 10364 11246 10384
rect 11006 10362 11030 10364
rect 11086 10362 11110 10364
rect 11166 10362 11190 10364
rect 11028 10310 11030 10362
rect 11092 10310 11104 10362
rect 11166 10310 11168 10362
rect 11006 10308 11030 10310
rect 11086 10308 11110 10310
rect 11166 10308 11190 10310
rect 10950 10288 11246 10308
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10950 9276 11246 9296
rect 11006 9274 11030 9276
rect 11086 9274 11110 9276
rect 11166 9274 11190 9276
rect 11028 9222 11030 9274
rect 11092 9222 11104 9274
rect 11166 9222 11168 9274
rect 11006 9220 11030 9222
rect 11086 9220 11110 9222
rect 11166 9220 11190 9222
rect 10950 9200 11246 9220
rect 10950 8188 11246 8208
rect 11006 8186 11030 8188
rect 11086 8186 11110 8188
rect 11166 8186 11190 8188
rect 11028 8134 11030 8186
rect 11092 8134 11104 8186
rect 11166 8134 11168 8186
rect 11006 8132 11030 8134
rect 11086 8132 11110 8134
rect 11166 8132 11190 8134
rect 10950 8112 11246 8132
rect 10950 7100 11246 7120
rect 11006 7098 11030 7100
rect 11086 7098 11110 7100
rect 11166 7098 11190 7100
rect 11028 7046 11030 7098
rect 11092 7046 11104 7098
rect 11166 7046 11168 7098
rect 11006 7044 11030 7046
rect 11086 7044 11110 7046
rect 11166 7044 11190 7046
rect 10950 7024 11246 7044
rect 10950 6012 11246 6032
rect 11006 6010 11030 6012
rect 11086 6010 11110 6012
rect 11166 6010 11190 6012
rect 11028 5958 11030 6010
rect 11092 5958 11104 6010
rect 11166 5958 11168 6010
rect 11006 5956 11030 5958
rect 11086 5956 11110 5958
rect 11166 5956 11190 5958
rect 10950 5936 11246 5956
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10336 2746 10548 2774
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10244 2310 10272 2586
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10336 2038 10364 2746
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10140 2032 10192 2038
rect 10140 1974 10192 1980
rect 10324 2032 10376 2038
rect 10324 1974 10376 1980
rect 10428 1766 10456 2246
rect 10416 1760 10468 1766
rect 10416 1702 10468 1708
rect 10520 800 10548 2450
rect 10612 1834 10640 5238
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10796 4758 10824 5102
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10888 4162 10916 5510
rect 11716 5370 11744 16546
rect 11808 5778 11836 16662
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11992 5370 12020 17886
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12268 16998 12296 17682
rect 12360 17218 12388 19200
rect 12360 17190 12480 17218
rect 12452 17134 12480 17190
rect 12728 17134 12756 19200
rect 13188 17134 13216 19200
rect 13556 17762 13584 19200
rect 13372 17734 13584 17762
rect 13372 17218 13400 17734
rect 13449 17436 13745 17456
rect 13505 17434 13529 17436
rect 13585 17434 13609 17436
rect 13665 17434 13689 17436
rect 13527 17382 13529 17434
rect 13591 17382 13603 17434
rect 13665 17382 13667 17434
rect 13505 17380 13529 17382
rect 13585 17380 13609 17382
rect 13665 17380 13689 17382
rect 13449 17360 13745 17380
rect 13372 17190 13492 17218
rect 13464 17134 13492 17190
rect 14016 17134 14044 19200
rect 14476 17134 14504 19200
rect 14844 17134 14872 19200
rect 15304 17134 15332 19200
rect 15672 17626 15700 19200
rect 15672 17598 15792 17626
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15658 17504 15714 17513
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14464 17128 14516 17134
rect 14832 17128 14884 17134
rect 14464 17070 14516 17076
rect 14752 17076 14832 17082
rect 14752 17070 14884 17076
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12176 16658 12204 16934
rect 12728 16794 12756 17070
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12544 9110 12572 11630
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12636 5370 12664 16186
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11808 5137 11836 5170
rect 12348 5160 12400 5166
rect 11794 5128 11850 5137
rect 11152 5092 11204 5098
rect 11204 5052 11376 5080
rect 12348 5102 12400 5108
rect 12438 5128 12494 5137
rect 11794 5063 11850 5072
rect 11152 5034 11204 5040
rect 10950 4924 11246 4944
rect 11006 4922 11030 4924
rect 11086 4922 11110 4924
rect 11166 4922 11190 4924
rect 11028 4870 11030 4922
rect 11092 4870 11104 4922
rect 11166 4870 11168 4922
rect 11006 4868 11030 4870
rect 11086 4868 11110 4870
rect 11166 4868 11190 4870
rect 10950 4848 11246 4868
rect 11348 4622 11376 5052
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 10704 4134 10916 4162
rect 10704 2650 10732 4134
rect 10980 4026 11008 4558
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 10796 3998 11008 4026
rect 10796 2650 10824 3998
rect 10950 3836 11246 3856
rect 11006 3834 11030 3836
rect 11086 3834 11110 3836
rect 11166 3834 11190 3836
rect 11028 3782 11030 3834
rect 11092 3782 11104 3834
rect 11166 3782 11168 3834
rect 11006 3780 11030 3782
rect 11086 3780 11110 3782
rect 11166 3780 11190 3782
rect 10950 3760 11246 3780
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10888 2496 10916 2790
rect 10950 2748 11246 2768
rect 11006 2746 11030 2748
rect 11086 2746 11110 2748
rect 11166 2746 11190 2748
rect 11028 2694 11030 2746
rect 11092 2694 11104 2746
rect 11166 2694 11168 2746
rect 11006 2692 11030 2694
rect 11086 2692 11110 2694
rect 11166 2692 11190 2694
rect 10950 2672 11246 2692
rect 11060 2508 11112 2514
rect 10888 2468 11060 2496
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 10888 800 10916 2468
rect 11060 2450 11112 2456
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11348 2310 11376 2450
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11348 800 11376 2246
rect 11440 2106 11468 4150
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11532 2650 11560 4082
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11808 2514 11836 2790
rect 11900 2650 11928 4558
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11428 2100 11480 2106
rect 11428 2042 11480 2048
rect 11808 800 11836 2450
rect 12084 2378 12112 4490
rect 12176 4214 12204 4966
rect 12360 4826 12388 5102
rect 12438 5063 12494 5072
rect 12716 5092 12768 5098
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 12176 800 12204 2450
rect 12268 2310 12296 2450
rect 12452 2378 12480 5063
rect 12716 5034 12768 5040
rect 12728 4622 12756 5034
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12636 2514 12664 2790
rect 12912 2650 12940 5306
rect 13096 5166 13124 15846
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13280 8838 13308 8978
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 7449 13308 8774
rect 13266 7440 13322 7449
rect 13266 7375 13322 7384
rect 13372 6914 13400 16934
rect 13449 16348 13745 16368
rect 13505 16346 13529 16348
rect 13585 16346 13609 16348
rect 13665 16346 13689 16348
rect 13527 16294 13529 16346
rect 13591 16294 13603 16346
rect 13665 16294 13667 16346
rect 13505 16292 13529 16294
rect 13585 16292 13609 16294
rect 13665 16292 13689 16294
rect 13449 16272 13745 16292
rect 13449 15260 13745 15280
rect 13505 15258 13529 15260
rect 13585 15258 13609 15260
rect 13665 15258 13689 15260
rect 13527 15206 13529 15258
rect 13591 15206 13603 15258
rect 13665 15206 13667 15258
rect 13505 15204 13529 15206
rect 13585 15204 13609 15206
rect 13665 15204 13689 15206
rect 13449 15184 13745 15204
rect 13449 14172 13745 14192
rect 13505 14170 13529 14172
rect 13585 14170 13609 14172
rect 13665 14170 13689 14172
rect 13527 14118 13529 14170
rect 13591 14118 13603 14170
rect 13665 14118 13667 14170
rect 13505 14116 13529 14118
rect 13585 14116 13609 14118
rect 13665 14116 13689 14118
rect 13449 14096 13745 14116
rect 13449 13084 13745 13104
rect 13505 13082 13529 13084
rect 13585 13082 13609 13084
rect 13665 13082 13689 13084
rect 13527 13030 13529 13082
rect 13591 13030 13603 13082
rect 13665 13030 13667 13082
rect 13505 13028 13529 13030
rect 13585 13028 13609 13030
rect 13665 13028 13689 13030
rect 13449 13008 13745 13028
rect 13449 11996 13745 12016
rect 13505 11994 13529 11996
rect 13585 11994 13609 11996
rect 13665 11994 13689 11996
rect 13527 11942 13529 11994
rect 13591 11942 13603 11994
rect 13665 11942 13667 11994
rect 13505 11940 13529 11942
rect 13585 11940 13609 11942
rect 13665 11940 13689 11942
rect 13449 11920 13745 11940
rect 13449 10908 13745 10928
rect 13505 10906 13529 10908
rect 13585 10906 13609 10908
rect 13665 10906 13689 10908
rect 13527 10854 13529 10906
rect 13591 10854 13603 10906
rect 13665 10854 13667 10906
rect 13505 10852 13529 10854
rect 13585 10852 13609 10854
rect 13665 10852 13689 10854
rect 13449 10832 13745 10852
rect 13449 9820 13745 9840
rect 13505 9818 13529 9820
rect 13585 9818 13609 9820
rect 13665 9818 13689 9820
rect 13527 9766 13529 9818
rect 13591 9766 13603 9818
rect 13665 9766 13667 9818
rect 13505 9764 13529 9766
rect 13585 9764 13609 9766
rect 13665 9764 13689 9766
rect 13449 9744 13745 9764
rect 13449 8732 13745 8752
rect 13505 8730 13529 8732
rect 13585 8730 13609 8732
rect 13665 8730 13689 8732
rect 13527 8678 13529 8730
rect 13591 8678 13603 8730
rect 13665 8678 13667 8730
rect 13505 8676 13529 8678
rect 13585 8676 13609 8678
rect 13665 8676 13689 8678
rect 13449 8656 13745 8676
rect 13449 7644 13745 7664
rect 13505 7642 13529 7644
rect 13585 7642 13609 7644
rect 13665 7642 13689 7644
rect 13527 7590 13529 7642
rect 13591 7590 13603 7642
rect 13665 7590 13667 7642
rect 13505 7588 13529 7590
rect 13585 7588 13609 7590
rect 13665 7588 13689 7590
rect 13449 7568 13745 7588
rect 13280 6886 13400 6914
rect 13280 5710 13308 6886
rect 13449 6556 13745 6576
rect 13505 6554 13529 6556
rect 13585 6554 13609 6556
rect 13665 6554 13689 6556
rect 13527 6502 13529 6554
rect 13591 6502 13603 6554
rect 13665 6502 13667 6554
rect 13505 6500 13529 6502
rect 13585 6500 13609 6502
rect 13665 6500 13689 6502
rect 13449 6480 13745 6500
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 14016 5642 14044 16934
rect 14384 16794 14412 17070
rect 14476 16794 14504 17070
rect 14752 17054 14872 17070
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14568 5914 14596 16934
rect 14752 16794 14780 17054
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 13449 5468 13745 5488
rect 13505 5466 13529 5468
rect 13585 5466 13609 5468
rect 13665 5466 13689 5468
rect 13527 5414 13529 5466
rect 13591 5414 13603 5466
rect 13665 5414 13667 5466
rect 13505 5412 13529 5414
rect 13585 5412 13609 5414
rect 13665 5412 13689 5414
rect 13449 5392 13745 5412
rect 14844 5234 14872 16934
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14936 5166 14964 16390
rect 15028 16250 15056 16526
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15120 5846 15148 16934
rect 15304 16250 15332 17070
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15488 13530 15516 17002
rect 15580 16658 15608 17478
rect 15658 17439 15714 17448
rect 15672 17270 15700 17439
rect 15660 17264 15712 17270
rect 15660 17206 15712 17212
rect 15764 16658 15792 17598
rect 16132 17542 16160 19200
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15580 15706 15608 16594
rect 15764 16182 15792 16594
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 16500 16046 16528 19200
rect 16960 16590 16988 19200
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15212 13190 15240 13330
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15212 11014 15240 13126
rect 15658 12472 15714 12481
rect 15658 12407 15714 12416
rect 15672 12374 15700 12407
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13449 4380 13745 4400
rect 13505 4378 13529 4380
rect 13585 4378 13609 4380
rect 13665 4378 13689 4380
rect 13527 4326 13529 4378
rect 13591 4326 13603 4378
rect 13665 4326 13667 4378
rect 13505 4324 13529 4326
rect 13585 4324 13609 4326
rect 13665 4324 13689 4326
rect 13449 4304 13745 4324
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13280 2650 13308 4218
rect 13449 3292 13745 3312
rect 13505 3290 13529 3292
rect 13585 3290 13609 3292
rect 13665 3290 13689 3292
rect 13527 3238 13529 3290
rect 13591 3238 13603 3290
rect 13665 3238 13667 3290
rect 13505 3236 13529 3238
rect 13585 3236 13609 3238
rect 13665 3236 13689 3238
rect 13449 3216 13745 3236
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13372 2514 13400 2790
rect 13832 2650 13860 4626
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13924 2514 13952 2858
rect 14200 2650 14228 4762
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14292 2514 14320 3062
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14384 2530 14412 2790
rect 14568 2650 14596 4422
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14752 2530 14780 2790
rect 14844 2650 14872 4694
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15120 2650 15148 4558
rect 15212 3738 15240 10950
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15212 3074 15240 3674
rect 15304 3194 15332 5238
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15488 3738 15516 5034
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15212 3046 15332 3074
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 14384 2514 14504 2530
rect 14752 2514 14872 2530
rect 15212 2514 15240 2926
rect 15304 2650 15332 3046
rect 15396 2990 15424 3334
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14384 2508 14516 2514
rect 14384 2502 14464 2508
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12636 800 12664 2450
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13004 2106 13032 2246
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 13096 800 13124 2450
rect 13372 1986 13400 2450
rect 13449 2204 13745 2224
rect 13505 2202 13529 2204
rect 13585 2202 13609 2204
rect 13665 2202 13689 2204
rect 13527 2150 13529 2202
rect 13591 2150 13603 2202
rect 13665 2150 13667 2202
rect 13505 2148 13529 2150
rect 13585 2148 13609 2150
rect 13665 2148 13689 2150
rect 13449 2128 13745 2148
rect 13372 1958 13492 1986
rect 13464 800 13492 1958
rect 13924 800 13952 2450
rect 14384 800 14412 2502
rect 14464 2450 14516 2456
rect 14752 2508 14884 2514
rect 14752 2502 14832 2508
rect 14752 800 14780 2502
rect 14832 2450 14884 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15212 800 15240 2450
rect 15580 2394 15608 2926
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 15658 2544 15714 2553
rect 15658 2479 15660 2488
rect 15712 2479 15714 2488
rect 15660 2450 15712 2456
rect 15580 2366 15700 2394
rect 15672 800 15700 2366
rect 16040 800 16068 2858
rect 16500 800 16528 3062
rect 16960 800 16988 3538
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
<< via2 >>
rect 1674 18264 1730 18320
rect 3454 17434 3510 17436
rect 3534 17434 3590 17436
rect 3614 17434 3670 17436
rect 3694 17434 3750 17436
rect 3454 17382 3480 17434
rect 3480 17382 3510 17434
rect 3534 17382 3544 17434
rect 3544 17382 3590 17434
rect 3614 17382 3660 17434
rect 3660 17382 3670 17434
rect 3694 17382 3724 17434
rect 3724 17382 3750 17434
rect 3454 17380 3510 17382
rect 3534 17380 3590 17382
rect 3614 17380 3670 17382
rect 3694 17380 3750 17382
rect 1398 15020 1454 15056
rect 1398 15000 1400 15020
rect 1400 15000 1452 15020
rect 1452 15000 1454 15020
rect 1398 11636 1400 11656
rect 1400 11636 1452 11656
rect 1452 11636 1454 11656
rect 1398 11600 1454 11636
rect 1398 8356 1454 8392
rect 1398 8336 1400 8356
rect 1400 8336 1452 8356
rect 1452 8336 1454 8356
rect 3454 16346 3510 16348
rect 3534 16346 3590 16348
rect 3614 16346 3670 16348
rect 3694 16346 3750 16348
rect 3454 16294 3480 16346
rect 3480 16294 3510 16346
rect 3534 16294 3544 16346
rect 3544 16294 3590 16346
rect 3614 16294 3660 16346
rect 3660 16294 3670 16346
rect 3694 16294 3724 16346
rect 3724 16294 3750 16346
rect 3454 16292 3510 16294
rect 3534 16292 3590 16294
rect 3614 16292 3670 16294
rect 3694 16292 3750 16294
rect 3454 15258 3510 15260
rect 3534 15258 3590 15260
rect 3614 15258 3670 15260
rect 3694 15258 3750 15260
rect 3454 15206 3480 15258
rect 3480 15206 3510 15258
rect 3534 15206 3544 15258
rect 3544 15206 3590 15258
rect 3614 15206 3660 15258
rect 3660 15206 3670 15258
rect 3694 15206 3724 15258
rect 3724 15206 3750 15258
rect 3454 15204 3510 15206
rect 3534 15204 3590 15206
rect 3614 15204 3670 15206
rect 3694 15204 3750 15206
rect 3454 14170 3510 14172
rect 3534 14170 3590 14172
rect 3614 14170 3670 14172
rect 3694 14170 3750 14172
rect 3454 14118 3480 14170
rect 3480 14118 3510 14170
rect 3534 14118 3544 14170
rect 3544 14118 3590 14170
rect 3614 14118 3660 14170
rect 3660 14118 3670 14170
rect 3694 14118 3724 14170
rect 3724 14118 3750 14170
rect 3454 14116 3510 14118
rect 3534 14116 3590 14118
rect 3614 14116 3670 14118
rect 3694 14116 3750 14118
rect 3454 13082 3510 13084
rect 3534 13082 3590 13084
rect 3614 13082 3670 13084
rect 3694 13082 3750 13084
rect 3454 13030 3480 13082
rect 3480 13030 3510 13082
rect 3534 13030 3544 13082
rect 3544 13030 3590 13082
rect 3614 13030 3660 13082
rect 3660 13030 3670 13082
rect 3694 13030 3724 13082
rect 3724 13030 3750 13082
rect 3454 13028 3510 13030
rect 3534 13028 3590 13030
rect 3614 13028 3670 13030
rect 3694 13028 3750 13030
rect 3454 11994 3510 11996
rect 3534 11994 3590 11996
rect 3614 11994 3670 11996
rect 3694 11994 3750 11996
rect 3454 11942 3480 11994
rect 3480 11942 3510 11994
rect 3534 11942 3544 11994
rect 3544 11942 3590 11994
rect 3614 11942 3660 11994
rect 3660 11942 3670 11994
rect 3694 11942 3724 11994
rect 3724 11942 3750 11994
rect 3454 11940 3510 11942
rect 3534 11940 3590 11942
rect 3614 11940 3670 11942
rect 3694 11940 3750 11942
rect 3454 10906 3510 10908
rect 3534 10906 3590 10908
rect 3614 10906 3670 10908
rect 3694 10906 3750 10908
rect 3454 10854 3480 10906
rect 3480 10854 3510 10906
rect 3534 10854 3544 10906
rect 3544 10854 3590 10906
rect 3614 10854 3660 10906
rect 3660 10854 3670 10906
rect 3694 10854 3724 10906
rect 3724 10854 3750 10906
rect 3454 10852 3510 10854
rect 3534 10852 3590 10854
rect 3614 10852 3670 10854
rect 3694 10852 3750 10854
rect 3454 9818 3510 9820
rect 3534 9818 3590 9820
rect 3614 9818 3670 9820
rect 3694 9818 3750 9820
rect 3454 9766 3480 9818
rect 3480 9766 3510 9818
rect 3534 9766 3544 9818
rect 3544 9766 3590 9818
rect 3614 9766 3660 9818
rect 3660 9766 3670 9818
rect 3694 9766 3724 9818
rect 3724 9766 3750 9818
rect 3454 9764 3510 9766
rect 3534 9764 3590 9766
rect 3614 9764 3670 9766
rect 3694 9764 3750 9766
rect 3454 8730 3510 8732
rect 3534 8730 3590 8732
rect 3614 8730 3670 8732
rect 3694 8730 3750 8732
rect 3454 8678 3480 8730
rect 3480 8678 3510 8730
rect 3534 8678 3544 8730
rect 3544 8678 3590 8730
rect 3614 8678 3660 8730
rect 3660 8678 3670 8730
rect 3694 8678 3724 8730
rect 3724 8678 3750 8730
rect 3454 8676 3510 8678
rect 3534 8676 3590 8678
rect 3614 8676 3670 8678
rect 3694 8676 3750 8678
rect 1490 4972 1492 4992
rect 1492 4972 1544 4992
rect 1544 4972 1546 4992
rect 1490 4936 1546 4972
rect 3454 7642 3510 7644
rect 3534 7642 3590 7644
rect 3614 7642 3670 7644
rect 3694 7642 3750 7644
rect 3454 7590 3480 7642
rect 3480 7590 3510 7642
rect 3534 7590 3544 7642
rect 3544 7590 3590 7642
rect 3614 7590 3660 7642
rect 3660 7590 3670 7642
rect 3694 7590 3724 7642
rect 3724 7590 3750 7642
rect 3454 7588 3510 7590
rect 3534 7588 3590 7590
rect 3614 7588 3670 7590
rect 3694 7588 3750 7590
rect 3454 6554 3510 6556
rect 3534 6554 3590 6556
rect 3614 6554 3670 6556
rect 3694 6554 3750 6556
rect 3454 6502 3480 6554
rect 3480 6502 3510 6554
rect 3534 6502 3544 6554
rect 3544 6502 3590 6554
rect 3614 6502 3660 6554
rect 3660 6502 3670 6554
rect 3694 6502 3724 6554
rect 3724 6502 3750 6554
rect 3454 6500 3510 6502
rect 3534 6500 3590 6502
rect 3614 6500 3670 6502
rect 3694 6500 3750 6502
rect 3454 5466 3510 5468
rect 3534 5466 3590 5468
rect 3614 5466 3670 5468
rect 3694 5466 3750 5468
rect 3454 5414 3480 5466
rect 3480 5414 3510 5466
rect 3534 5414 3544 5466
rect 3544 5414 3590 5466
rect 3614 5414 3660 5466
rect 3660 5414 3670 5466
rect 3694 5414 3724 5466
rect 3724 5414 3750 5466
rect 3454 5412 3510 5414
rect 3534 5412 3590 5414
rect 3614 5412 3670 5414
rect 3694 5412 3750 5414
rect 3454 4378 3510 4380
rect 3534 4378 3590 4380
rect 3614 4378 3670 4380
rect 3694 4378 3750 4380
rect 3454 4326 3480 4378
rect 3480 4326 3510 4378
rect 3534 4326 3544 4378
rect 3544 4326 3590 4378
rect 3614 4326 3660 4378
rect 3660 4326 3670 4378
rect 3694 4326 3724 4378
rect 3724 4326 3750 4378
rect 3454 4324 3510 4326
rect 3534 4324 3590 4326
rect 3614 4324 3670 4326
rect 3694 4324 3750 4326
rect 3454 3290 3510 3292
rect 3534 3290 3590 3292
rect 3614 3290 3670 3292
rect 3694 3290 3750 3292
rect 3454 3238 3480 3290
rect 3480 3238 3510 3290
rect 3534 3238 3544 3290
rect 3544 3238 3590 3290
rect 3614 3238 3660 3290
rect 3660 3238 3670 3290
rect 3694 3238 3724 3290
rect 3724 3238 3750 3290
rect 3454 3236 3510 3238
rect 3534 3236 3590 3238
rect 3614 3236 3670 3238
rect 3694 3236 3750 3238
rect 1674 1672 1730 1728
rect 3454 2202 3510 2204
rect 3534 2202 3590 2204
rect 3614 2202 3670 2204
rect 3694 2202 3750 2204
rect 3454 2150 3480 2202
rect 3480 2150 3510 2202
rect 3534 2150 3544 2202
rect 3544 2150 3590 2202
rect 3614 2150 3660 2202
rect 3660 2150 3670 2202
rect 3694 2150 3724 2202
rect 3724 2150 3750 2202
rect 3454 2148 3510 2150
rect 3534 2148 3590 2150
rect 3614 2148 3670 2150
rect 3694 2148 3750 2150
rect 5953 16890 6009 16892
rect 6033 16890 6089 16892
rect 6113 16890 6169 16892
rect 6193 16890 6249 16892
rect 5953 16838 5979 16890
rect 5979 16838 6009 16890
rect 6033 16838 6043 16890
rect 6043 16838 6089 16890
rect 6113 16838 6159 16890
rect 6159 16838 6169 16890
rect 6193 16838 6223 16890
rect 6223 16838 6249 16890
rect 5953 16836 6009 16838
rect 6033 16836 6089 16838
rect 6113 16836 6169 16838
rect 6193 16836 6249 16838
rect 5953 15802 6009 15804
rect 6033 15802 6089 15804
rect 6113 15802 6169 15804
rect 6193 15802 6249 15804
rect 5953 15750 5979 15802
rect 5979 15750 6009 15802
rect 6033 15750 6043 15802
rect 6043 15750 6089 15802
rect 6113 15750 6159 15802
rect 6159 15750 6169 15802
rect 6193 15750 6223 15802
rect 6223 15750 6249 15802
rect 5953 15748 6009 15750
rect 6033 15748 6089 15750
rect 6113 15748 6169 15750
rect 6193 15748 6249 15750
rect 5953 14714 6009 14716
rect 6033 14714 6089 14716
rect 6113 14714 6169 14716
rect 6193 14714 6249 14716
rect 5953 14662 5979 14714
rect 5979 14662 6009 14714
rect 6033 14662 6043 14714
rect 6043 14662 6089 14714
rect 6113 14662 6159 14714
rect 6159 14662 6169 14714
rect 6193 14662 6223 14714
rect 6223 14662 6249 14714
rect 5953 14660 6009 14662
rect 6033 14660 6089 14662
rect 6113 14660 6169 14662
rect 6193 14660 6249 14662
rect 5953 13626 6009 13628
rect 6033 13626 6089 13628
rect 6113 13626 6169 13628
rect 6193 13626 6249 13628
rect 5953 13574 5979 13626
rect 5979 13574 6009 13626
rect 6033 13574 6043 13626
rect 6043 13574 6089 13626
rect 6113 13574 6159 13626
rect 6159 13574 6169 13626
rect 6193 13574 6223 13626
rect 6223 13574 6249 13626
rect 5953 13572 6009 13574
rect 6033 13572 6089 13574
rect 6113 13572 6169 13574
rect 6193 13572 6249 13574
rect 5953 12538 6009 12540
rect 6033 12538 6089 12540
rect 6113 12538 6169 12540
rect 6193 12538 6249 12540
rect 5953 12486 5979 12538
rect 5979 12486 6009 12538
rect 6033 12486 6043 12538
rect 6043 12486 6089 12538
rect 6113 12486 6159 12538
rect 6159 12486 6169 12538
rect 6193 12486 6223 12538
rect 6223 12486 6249 12538
rect 5953 12484 6009 12486
rect 6033 12484 6089 12486
rect 6113 12484 6169 12486
rect 6193 12484 6249 12486
rect 5953 11450 6009 11452
rect 6033 11450 6089 11452
rect 6113 11450 6169 11452
rect 6193 11450 6249 11452
rect 5953 11398 5979 11450
rect 5979 11398 6009 11450
rect 6033 11398 6043 11450
rect 6043 11398 6089 11450
rect 6113 11398 6159 11450
rect 6159 11398 6169 11450
rect 6193 11398 6223 11450
rect 6223 11398 6249 11450
rect 5953 11396 6009 11398
rect 6033 11396 6089 11398
rect 6113 11396 6169 11398
rect 6193 11396 6249 11398
rect 5953 10362 6009 10364
rect 6033 10362 6089 10364
rect 6113 10362 6169 10364
rect 6193 10362 6249 10364
rect 5953 10310 5979 10362
rect 5979 10310 6009 10362
rect 6033 10310 6043 10362
rect 6043 10310 6089 10362
rect 6113 10310 6159 10362
rect 6159 10310 6169 10362
rect 6193 10310 6223 10362
rect 6223 10310 6249 10362
rect 5953 10308 6009 10310
rect 6033 10308 6089 10310
rect 6113 10308 6169 10310
rect 6193 10308 6249 10310
rect 5953 9274 6009 9276
rect 6033 9274 6089 9276
rect 6113 9274 6169 9276
rect 6193 9274 6249 9276
rect 5953 9222 5979 9274
rect 5979 9222 6009 9274
rect 6033 9222 6043 9274
rect 6043 9222 6089 9274
rect 6113 9222 6159 9274
rect 6159 9222 6169 9274
rect 6193 9222 6223 9274
rect 6223 9222 6249 9274
rect 5953 9220 6009 9222
rect 6033 9220 6089 9222
rect 6113 9220 6169 9222
rect 6193 9220 6249 9222
rect 5953 8186 6009 8188
rect 6033 8186 6089 8188
rect 6113 8186 6169 8188
rect 6193 8186 6249 8188
rect 5953 8134 5979 8186
rect 5979 8134 6009 8186
rect 6033 8134 6043 8186
rect 6043 8134 6089 8186
rect 6113 8134 6159 8186
rect 6159 8134 6169 8186
rect 6193 8134 6223 8186
rect 6223 8134 6249 8186
rect 5953 8132 6009 8134
rect 6033 8132 6089 8134
rect 6113 8132 6169 8134
rect 6193 8132 6249 8134
rect 5953 7098 6009 7100
rect 6033 7098 6089 7100
rect 6113 7098 6169 7100
rect 6193 7098 6249 7100
rect 5953 7046 5979 7098
rect 5979 7046 6009 7098
rect 6033 7046 6043 7098
rect 6043 7046 6089 7098
rect 6113 7046 6159 7098
rect 6159 7046 6169 7098
rect 6193 7046 6223 7098
rect 6223 7046 6249 7098
rect 5953 7044 6009 7046
rect 6033 7044 6089 7046
rect 6113 7044 6169 7046
rect 6193 7044 6249 7046
rect 5953 6010 6009 6012
rect 6033 6010 6089 6012
rect 6113 6010 6169 6012
rect 6193 6010 6249 6012
rect 5953 5958 5979 6010
rect 5979 5958 6009 6010
rect 6033 5958 6043 6010
rect 6043 5958 6089 6010
rect 6113 5958 6159 6010
rect 6159 5958 6169 6010
rect 6193 5958 6223 6010
rect 6223 5958 6249 6010
rect 5953 5956 6009 5958
rect 6033 5956 6089 5958
rect 6113 5956 6169 5958
rect 6193 5956 6249 5958
rect 6734 5208 6790 5264
rect 5998 5108 6000 5128
rect 6000 5108 6052 5128
rect 6052 5108 6054 5128
rect 5998 5072 6054 5108
rect 5953 4922 6009 4924
rect 6033 4922 6089 4924
rect 6113 4922 6169 4924
rect 6193 4922 6249 4924
rect 5953 4870 5979 4922
rect 5979 4870 6009 4922
rect 6033 4870 6043 4922
rect 6043 4870 6089 4922
rect 6113 4870 6159 4922
rect 6159 4870 6169 4922
rect 6193 4870 6223 4922
rect 6223 4870 6249 4922
rect 5953 4868 6009 4870
rect 6033 4868 6089 4870
rect 6113 4868 6169 4870
rect 6193 4868 6249 4870
rect 5953 3834 6009 3836
rect 6033 3834 6089 3836
rect 6113 3834 6169 3836
rect 6193 3834 6249 3836
rect 5953 3782 5979 3834
rect 5979 3782 6009 3834
rect 6033 3782 6043 3834
rect 6043 3782 6089 3834
rect 6113 3782 6159 3834
rect 6159 3782 6169 3834
rect 6193 3782 6223 3834
rect 6223 3782 6249 3834
rect 5953 3780 6009 3782
rect 6033 3780 6089 3782
rect 6113 3780 6169 3782
rect 6193 3780 6249 3782
rect 5953 2746 6009 2748
rect 6033 2746 6089 2748
rect 6113 2746 6169 2748
rect 6193 2746 6249 2748
rect 5953 2694 5979 2746
rect 5979 2694 6009 2746
rect 6033 2694 6043 2746
rect 6043 2694 6089 2746
rect 6113 2694 6159 2746
rect 6159 2694 6169 2746
rect 6193 2694 6223 2746
rect 6223 2694 6249 2746
rect 5953 2692 6009 2694
rect 6033 2692 6089 2694
rect 6113 2692 6169 2694
rect 6193 2692 6249 2694
rect 6826 4664 6882 4720
rect 7930 16632 7986 16688
rect 7930 5616 7986 5672
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8478 17434
rect 8478 17382 8508 17434
rect 8532 17382 8542 17434
rect 8542 17382 8588 17434
rect 8612 17382 8658 17434
rect 8658 17382 8668 17434
rect 8692 17382 8722 17434
rect 8722 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8666 16904 8722 16960
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8478 16346
rect 8478 16294 8508 16346
rect 8532 16294 8542 16346
rect 8542 16294 8588 16346
rect 8612 16294 8658 16346
rect 8658 16294 8668 16346
rect 8692 16294 8722 16346
rect 8722 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8478 15258
rect 8478 15206 8508 15258
rect 8532 15206 8542 15258
rect 8542 15206 8588 15258
rect 8612 15206 8658 15258
rect 8658 15206 8668 15258
rect 8692 15206 8722 15258
rect 8722 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8478 14170
rect 8478 14118 8508 14170
rect 8532 14118 8542 14170
rect 8542 14118 8588 14170
rect 8612 14118 8658 14170
rect 8658 14118 8668 14170
rect 8692 14118 8722 14170
rect 8722 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8478 13082
rect 8478 13030 8508 13082
rect 8532 13030 8542 13082
rect 8542 13030 8588 13082
rect 8612 13030 8658 13082
rect 8658 13030 8668 13082
rect 8692 13030 8722 13082
rect 8722 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8478 11994
rect 8478 11942 8508 11994
rect 8532 11942 8542 11994
rect 8542 11942 8588 11994
rect 8612 11942 8658 11994
rect 8658 11942 8668 11994
rect 8692 11942 8722 11994
rect 8722 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8478 10906
rect 8478 10854 8508 10906
rect 8532 10854 8542 10906
rect 8542 10854 8588 10906
rect 8612 10854 8658 10906
rect 8658 10854 8668 10906
rect 8692 10854 8722 10906
rect 8722 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8478 9818
rect 8478 9766 8508 9818
rect 8532 9766 8542 9818
rect 8542 9766 8588 9818
rect 8612 9766 8658 9818
rect 8658 9766 8668 9818
rect 8692 9766 8722 9818
rect 8722 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8478 8730
rect 8478 8678 8508 8730
rect 8532 8678 8542 8730
rect 8542 8678 8588 8730
rect 8612 8678 8658 8730
rect 8658 8678 8668 8730
rect 8692 8678 8722 8730
rect 8722 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8478 7642
rect 8478 7590 8508 7642
rect 8532 7590 8542 7642
rect 8542 7590 8588 7642
rect 8612 7590 8658 7642
rect 8658 7590 8668 7642
rect 8692 7590 8722 7642
rect 8722 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8478 6554
rect 8478 6502 8508 6554
rect 8532 6502 8542 6554
rect 8542 6502 8588 6554
rect 8612 6502 8658 6554
rect 8658 6502 8668 6554
rect 8692 6502 8722 6554
rect 8722 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8478 5466
rect 8478 5414 8508 5466
rect 8532 5414 8542 5466
rect 8542 5414 8588 5466
rect 8612 5414 8658 5466
rect 8658 5414 8668 5466
rect 8692 5414 8722 5466
rect 8722 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8478 4378
rect 8478 4326 8508 4378
rect 8532 4326 8542 4378
rect 8542 4326 8588 4378
rect 8612 4326 8658 4378
rect 8658 4326 8668 4378
rect 8692 4326 8722 4378
rect 8722 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8478 3290
rect 8478 3238 8508 3290
rect 8532 3238 8542 3290
rect 8542 3238 8588 3290
rect 8612 3238 8658 3290
rect 8658 3238 8668 3290
rect 8692 3238 8722 3290
rect 8722 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8478 2202
rect 8478 2150 8508 2202
rect 8532 2150 8542 2202
rect 8542 2150 8588 2202
rect 8612 2150 8658 2202
rect 8658 2150 8668 2202
rect 8692 2150 8722 2202
rect 8722 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9494 5616 9550 5672
rect 10322 16904 10378 16960
rect 9954 5244 9956 5264
rect 9956 5244 10008 5264
rect 10008 5244 10010 5264
rect 9954 5208 10010 5244
rect 9494 5072 9550 5128
rect 9494 4664 9550 4720
rect 10950 16890 11006 16892
rect 11030 16890 11086 16892
rect 11110 16890 11166 16892
rect 11190 16890 11246 16892
rect 10950 16838 10976 16890
rect 10976 16838 11006 16890
rect 11030 16838 11040 16890
rect 11040 16838 11086 16890
rect 11110 16838 11156 16890
rect 11156 16838 11166 16890
rect 11190 16838 11220 16890
rect 11220 16838 11246 16890
rect 10950 16836 11006 16838
rect 11030 16836 11086 16838
rect 11110 16836 11166 16838
rect 11190 16836 11246 16838
rect 10782 16652 10838 16688
rect 10782 16632 10784 16652
rect 10784 16632 10836 16652
rect 10836 16632 10838 16652
rect 10950 15802 11006 15804
rect 11030 15802 11086 15804
rect 11110 15802 11166 15804
rect 11190 15802 11246 15804
rect 10950 15750 10976 15802
rect 10976 15750 11006 15802
rect 11030 15750 11040 15802
rect 11040 15750 11086 15802
rect 11110 15750 11156 15802
rect 11156 15750 11166 15802
rect 11190 15750 11220 15802
rect 11220 15750 11246 15802
rect 10950 15748 11006 15750
rect 11030 15748 11086 15750
rect 11110 15748 11166 15750
rect 11190 15748 11246 15750
rect 10950 14714 11006 14716
rect 11030 14714 11086 14716
rect 11110 14714 11166 14716
rect 11190 14714 11246 14716
rect 10950 14662 10976 14714
rect 10976 14662 11006 14714
rect 11030 14662 11040 14714
rect 11040 14662 11086 14714
rect 11110 14662 11156 14714
rect 11156 14662 11166 14714
rect 11190 14662 11220 14714
rect 11220 14662 11246 14714
rect 10950 14660 11006 14662
rect 11030 14660 11086 14662
rect 11110 14660 11166 14662
rect 11190 14660 11246 14662
rect 10950 13626 11006 13628
rect 11030 13626 11086 13628
rect 11110 13626 11166 13628
rect 11190 13626 11246 13628
rect 10950 13574 10976 13626
rect 10976 13574 11006 13626
rect 11030 13574 11040 13626
rect 11040 13574 11086 13626
rect 11110 13574 11156 13626
rect 11156 13574 11166 13626
rect 11190 13574 11220 13626
rect 11220 13574 11246 13626
rect 10950 13572 11006 13574
rect 11030 13572 11086 13574
rect 11110 13572 11166 13574
rect 11190 13572 11246 13574
rect 10950 12538 11006 12540
rect 11030 12538 11086 12540
rect 11110 12538 11166 12540
rect 11190 12538 11246 12540
rect 10950 12486 10976 12538
rect 10976 12486 11006 12538
rect 11030 12486 11040 12538
rect 11040 12486 11086 12538
rect 11110 12486 11156 12538
rect 11156 12486 11166 12538
rect 11190 12486 11220 12538
rect 11220 12486 11246 12538
rect 10950 12484 11006 12486
rect 11030 12484 11086 12486
rect 11110 12484 11166 12486
rect 11190 12484 11246 12486
rect 10950 11450 11006 11452
rect 11030 11450 11086 11452
rect 11110 11450 11166 11452
rect 11190 11450 11246 11452
rect 10950 11398 10976 11450
rect 10976 11398 11006 11450
rect 11030 11398 11040 11450
rect 11040 11398 11086 11450
rect 11110 11398 11156 11450
rect 11156 11398 11166 11450
rect 11190 11398 11220 11450
rect 11220 11398 11246 11450
rect 10950 11396 11006 11398
rect 11030 11396 11086 11398
rect 11110 11396 11166 11398
rect 11190 11396 11246 11398
rect 10950 10362 11006 10364
rect 11030 10362 11086 10364
rect 11110 10362 11166 10364
rect 11190 10362 11246 10364
rect 10950 10310 10976 10362
rect 10976 10310 11006 10362
rect 11030 10310 11040 10362
rect 11040 10310 11086 10362
rect 11110 10310 11156 10362
rect 11156 10310 11166 10362
rect 11190 10310 11220 10362
rect 11220 10310 11246 10362
rect 10950 10308 11006 10310
rect 11030 10308 11086 10310
rect 11110 10308 11166 10310
rect 11190 10308 11246 10310
rect 10950 9274 11006 9276
rect 11030 9274 11086 9276
rect 11110 9274 11166 9276
rect 11190 9274 11246 9276
rect 10950 9222 10976 9274
rect 10976 9222 11006 9274
rect 11030 9222 11040 9274
rect 11040 9222 11086 9274
rect 11110 9222 11156 9274
rect 11156 9222 11166 9274
rect 11190 9222 11220 9274
rect 11220 9222 11246 9274
rect 10950 9220 11006 9222
rect 11030 9220 11086 9222
rect 11110 9220 11166 9222
rect 11190 9220 11246 9222
rect 10950 8186 11006 8188
rect 11030 8186 11086 8188
rect 11110 8186 11166 8188
rect 11190 8186 11246 8188
rect 10950 8134 10976 8186
rect 10976 8134 11006 8186
rect 11030 8134 11040 8186
rect 11040 8134 11086 8186
rect 11110 8134 11156 8186
rect 11156 8134 11166 8186
rect 11190 8134 11220 8186
rect 11220 8134 11246 8186
rect 10950 8132 11006 8134
rect 11030 8132 11086 8134
rect 11110 8132 11166 8134
rect 11190 8132 11246 8134
rect 10950 7098 11006 7100
rect 11030 7098 11086 7100
rect 11110 7098 11166 7100
rect 11190 7098 11246 7100
rect 10950 7046 10976 7098
rect 10976 7046 11006 7098
rect 11030 7046 11040 7098
rect 11040 7046 11086 7098
rect 11110 7046 11156 7098
rect 11156 7046 11166 7098
rect 11190 7046 11220 7098
rect 11220 7046 11246 7098
rect 10950 7044 11006 7046
rect 11030 7044 11086 7046
rect 11110 7044 11166 7046
rect 11190 7044 11246 7046
rect 10950 6010 11006 6012
rect 11030 6010 11086 6012
rect 11110 6010 11166 6012
rect 11190 6010 11246 6012
rect 10950 5958 10976 6010
rect 10976 5958 11006 6010
rect 11030 5958 11040 6010
rect 11040 5958 11086 6010
rect 11110 5958 11156 6010
rect 11156 5958 11166 6010
rect 11190 5958 11220 6010
rect 11220 5958 11246 6010
rect 10950 5956 11006 5958
rect 11030 5956 11086 5958
rect 11110 5956 11166 5958
rect 11190 5956 11246 5958
rect 13449 17434 13505 17436
rect 13529 17434 13585 17436
rect 13609 17434 13665 17436
rect 13689 17434 13745 17436
rect 13449 17382 13475 17434
rect 13475 17382 13505 17434
rect 13529 17382 13539 17434
rect 13539 17382 13585 17434
rect 13609 17382 13655 17434
rect 13655 17382 13665 17434
rect 13689 17382 13719 17434
rect 13719 17382 13745 17434
rect 13449 17380 13505 17382
rect 13529 17380 13585 17382
rect 13609 17380 13665 17382
rect 13689 17380 13745 17382
rect 11794 5072 11850 5128
rect 10950 4922 11006 4924
rect 11030 4922 11086 4924
rect 11110 4922 11166 4924
rect 11190 4922 11246 4924
rect 10950 4870 10976 4922
rect 10976 4870 11006 4922
rect 11030 4870 11040 4922
rect 11040 4870 11086 4922
rect 11110 4870 11156 4922
rect 11156 4870 11166 4922
rect 11190 4870 11220 4922
rect 11220 4870 11246 4922
rect 10950 4868 11006 4870
rect 11030 4868 11086 4870
rect 11110 4868 11166 4870
rect 11190 4868 11246 4870
rect 10950 3834 11006 3836
rect 11030 3834 11086 3836
rect 11110 3834 11166 3836
rect 11190 3834 11246 3836
rect 10950 3782 10976 3834
rect 10976 3782 11006 3834
rect 11030 3782 11040 3834
rect 11040 3782 11086 3834
rect 11110 3782 11156 3834
rect 11156 3782 11166 3834
rect 11190 3782 11220 3834
rect 11220 3782 11246 3834
rect 10950 3780 11006 3782
rect 11030 3780 11086 3782
rect 11110 3780 11166 3782
rect 11190 3780 11246 3782
rect 10950 2746 11006 2748
rect 11030 2746 11086 2748
rect 11110 2746 11166 2748
rect 11190 2746 11246 2748
rect 10950 2694 10976 2746
rect 10976 2694 11006 2746
rect 11030 2694 11040 2746
rect 11040 2694 11086 2746
rect 11110 2694 11156 2746
rect 11156 2694 11166 2746
rect 11190 2694 11220 2746
rect 11220 2694 11246 2746
rect 10950 2692 11006 2694
rect 11030 2692 11086 2694
rect 11110 2692 11166 2694
rect 11190 2692 11246 2694
rect 12438 5072 12494 5128
rect 13266 7384 13322 7440
rect 13449 16346 13505 16348
rect 13529 16346 13585 16348
rect 13609 16346 13665 16348
rect 13689 16346 13745 16348
rect 13449 16294 13475 16346
rect 13475 16294 13505 16346
rect 13529 16294 13539 16346
rect 13539 16294 13585 16346
rect 13609 16294 13655 16346
rect 13655 16294 13665 16346
rect 13689 16294 13719 16346
rect 13719 16294 13745 16346
rect 13449 16292 13505 16294
rect 13529 16292 13585 16294
rect 13609 16292 13665 16294
rect 13689 16292 13745 16294
rect 13449 15258 13505 15260
rect 13529 15258 13585 15260
rect 13609 15258 13665 15260
rect 13689 15258 13745 15260
rect 13449 15206 13475 15258
rect 13475 15206 13505 15258
rect 13529 15206 13539 15258
rect 13539 15206 13585 15258
rect 13609 15206 13655 15258
rect 13655 15206 13665 15258
rect 13689 15206 13719 15258
rect 13719 15206 13745 15258
rect 13449 15204 13505 15206
rect 13529 15204 13585 15206
rect 13609 15204 13665 15206
rect 13689 15204 13745 15206
rect 13449 14170 13505 14172
rect 13529 14170 13585 14172
rect 13609 14170 13665 14172
rect 13689 14170 13745 14172
rect 13449 14118 13475 14170
rect 13475 14118 13505 14170
rect 13529 14118 13539 14170
rect 13539 14118 13585 14170
rect 13609 14118 13655 14170
rect 13655 14118 13665 14170
rect 13689 14118 13719 14170
rect 13719 14118 13745 14170
rect 13449 14116 13505 14118
rect 13529 14116 13585 14118
rect 13609 14116 13665 14118
rect 13689 14116 13745 14118
rect 13449 13082 13505 13084
rect 13529 13082 13585 13084
rect 13609 13082 13665 13084
rect 13689 13082 13745 13084
rect 13449 13030 13475 13082
rect 13475 13030 13505 13082
rect 13529 13030 13539 13082
rect 13539 13030 13585 13082
rect 13609 13030 13655 13082
rect 13655 13030 13665 13082
rect 13689 13030 13719 13082
rect 13719 13030 13745 13082
rect 13449 13028 13505 13030
rect 13529 13028 13585 13030
rect 13609 13028 13665 13030
rect 13689 13028 13745 13030
rect 13449 11994 13505 11996
rect 13529 11994 13585 11996
rect 13609 11994 13665 11996
rect 13689 11994 13745 11996
rect 13449 11942 13475 11994
rect 13475 11942 13505 11994
rect 13529 11942 13539 11994
rect 13539 11942 13585 11994
rect 13609 11942 13655 11994
rect 13655 11942 13665 11994
rect 13689 11942 13719 11994
rect 13719 11942 13745 11994
rect 13449 11940 13505 11942
rect 13529 11940 13585 11942
rect 13609 11940 13665 11942
rect 13689 11940 13745 11942
rect 13449 10906 13505 10908
rect 13529 10906 13585 10908
rect 13609 10906 13665 10908
rect 13689 10906 13745 10908
rect 13449 10854 13475 10906
rect 13475 10854 13505 10906
rect 13529 10854 13539 10906
rect 13539 10854 13585 10906
rect 13609 10854 13655 10906
rect 13655 10854 13665 10906
rect 13689 10854 13719 10906
rect 13719 10854 13745 10906
rect 13449 10852 13505 10854
rect 13529 10852 13585 10854
rect 13609 10852 13665 10854
rect 13689 10852 13745 10854
rect 13449 9818 13505 9820
rect 13529 9818 13585 9820
rect 13609 9818 13665 9820
rect 13689 9818 13745 9820
rect 13449 9766 13475 9818
rect 13475 9766 13505 9818
rect 13529 9766 13539 9818
rect 13539 9766 13585 9818
rect 13609 9766 13655 9818
rect 13655 9766 13665 9818
rect 13689 9766 13719 9818
rect 13719 9766 13745 9818
rect 13449 9764 13505 9766
rect 13529 9764 13585 9766
rect 13609 9764 13665 9766
rect 13689 9764 13745 9766
rect 13449 8730 13505 8732
rect 13529 8730 13585 8732
rect 13609 8730 13665 8732
rect 13689 8730 13745 8732
rect 13449 8678 13475 8730
rect 13475 8678 13505 8730
rect 13529 8678 13539 8730
rect 13539 8678 13585 8730
rect 13609 8678 13655 8730
rect 13655 8678 13665 8730
rect 13689 8678 13719 8730
rect 13719 8678 13745 8730
rect 13449 8676 13505 8678
rect 13529 8676 13585 8678
rect 13609 8676 13665 8678
rect 13689 8676 13745 8678
rect 13449 7642 13505 7644
rect 13529 7642 13585 7644
rect 13609 7642 13665 7644
rect 13689 7642 13745 7644
rect 13449 7590 13475 7642
rect 13475 7590 13505 7642
rect 13529 7590 13539 7642
rect 13539 7590 13585 7642
rect 13609 7590 13655 7642
rect 13655 7590 13665 7642
rect 13689 7590 13719 7642
rect 13719 7590 13745 7642
rect 13449 7588 13505 7590
rect 13529 7588 13585 7590
rect 13609 7588 13665 7590
rect 13689 7588 13745 7590
rect 13449 6554 13505 6556
rect 13529 6554 13585 6556
rect 13609 6554 13665 6556
rect 13689 6554 13745 6556
rect 13449 6502 13475 6554
rect 13475 6502 13505 6554
rect 13529 6502 13539 6554
rect 13539 6502 13585 6554
rect 13609 6502 13655 6554
rect 13655 6502 13665 6554
rect 13689 6502 13719 6554
rect 13719 6502 13745 6554
rect 13449 6500 13505 6502
rect 13529 6500 13585 6502
rect 13609 6500 13665 6502
rect 13689 6500 13745 6502
rect 13449 5466 13505 5468
rect 13529 5466 13585 5468
rect 13609 5466 13665 5468
rect 13689 5466 13745 5468
rect 13449 5414 13475 5466
rect 13475 5414 13505 5466
rect 13529 5414 13539 5466
rect 13539 5414 13585 5466
rect 13609 5414 13655 5466
rect 13655 5414 13665 5466
rect 13689 5414 13719 5466
rect 13719 5414 13745 5466
rect 13449 5412 13505 5414
rect 13529 5412 13585 5414
rect 13609 5412 13665 5414
rect 13689 5412 13745 5414
rect 15658 17448 15714 17504
rect 15658 12416 15714 12472
rect 13449 4378 13505 4380
rect 13529 4378 13585 4380
rect 13609 4378 13665 4380
rect 13689 4378 13745 4380
rect 13449 4326 13475 4378
rect 13475 4326 13505 4378
rect 13529 4326 13539 4378
rect 13539 4326 13585 4378
rect 13609 4326 13655 4378
rect 13655 4326 13665 4378
rect 13689 4326 13719 4378
rect 13719 4326 13745 4378
rect 13449 4324 13505 4326
rect 13529 4324 13585 4326
rect 13609 4324 13665 4326
rect 13689 4324 13745 4326
rect 13449 3290 13505 3292
rect 13529 3290 13585 3292
rect 13609 3290 13665 3292
rect 13689 3290 13745 3292
rect 13449 3238 13475 3290
rect 13475 3238 13505 3290
rect 13529 3238 13539 3290
rect 13539 3238 13585 3290
rect 13609 3238 13655 3290
rect 13655 3238 13665 3290
rect 13689 3238 13719 3290
rect 13719 3238 13745 3290
rect 13449 3236 13505 3238
rect 13529 3236 13585 3238
rect 13609 3236 13665 3238
rect 13689 3236 13745 3238
rect 13449 2202 13505 2204
rect 13529 2202 13585 2204
rect 13609 2202 13665 2204
rect 13689 2202 13745 2204
rect 13449 2150 13475 2202
rect 13475 2150 13505 2202
rect 13529 2150 13539 2202
rect 13539 2150 13585 2202
rect 13609 2150 13655 2202
rect 13655 2150 13665 2202
rect 13689 2150 13719 2202
rect 13719 2150 13745 2202
rect 13449 2148 13505 2150
rect 13529 2148 13585 2150
rect 13609 2148 13665 2150
rect 13689 2148 13745 2150
rect 15658 2508 15714 2544
rect 15658 2488 15660 2508
rect 15660 2488 15712 2508
rect 15712 2488 15714 2508
<< metal3 >>
rect 0 18322 800 18352
rect 1669 18322 1735 18325
rect 0 18320 1735 18322
rect 0 18264 1674 18320
rect 1730 18264 1735 18320
rect 0 18262 1735 18264
rect 0 18232 800 18262
rect 1669 18259 1735 18262
rect 15653 17506 15719 17509
rect 16400 17506 17200 17536
rect 15653 17504 17200 17506
rect 15653 17448 15658 17504
rect 15714 17448 17200 17504
rect 15653 17446 17200 17448
rect 15653 17443 15719 17446
rect 3442 17440 3762 17441
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3762 17440
rect 3442 17375 3762 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 13437 17440 13757 17441
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 16400 17416 17200 17446
rect 13437 17375 13757 17376
rect 8661 16962 8727 16965
rect 10317 16962 10383 16965
rect 8661 16960 10383 16962
rect 8661 16904 8666 16960
rect 8722 16904 10322 16960
rect 10378 16904 10383 16960
rect 8661 16902 10383 16904
rect 8661 16899 8727 16902
rect 10317 16899 10383 16902
rect 5941 16896 6261 16897
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 16831 6261 16832
rect 10938 16896 11258 16897
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11258 16896
rect 10938 16831 11258 16832
rect 7925 16690 7991 16693
rect 10777 16690 10843 16693
rect 7925 16688 10843 16690
rect 7925 16632 7930 16688
rect 7986 16632 10782 16688
rect 10838 16632 10843 16688
rect 7925 16630 10843 16632
rect 7925 16627 7991 16630
rect 10777 16627 10843 16630
rect 3442 16352 3762 16353
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3762 16352
rect 3442 16287 3762 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 13437 16352 13757 16353
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 16287 13757 16288
rect 5941 15808 6261 15809
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 15743 6261 15744
rect 10938 15808 11258 15809
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11258 15808
rect 10938 15743 11258 15744
rect 3442 15264 3762 15265
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3762 15264
rect 3442 15199 3762 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 13437 15264 13757 15265
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 15199 13757 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 5941 14720 6261 14721
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 14655 6261 14656
rect 10938 14720 11258 14721
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11258 14720
rect 10938 14655 11258 14656
rect 3442 14176 3762 14177
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3762 14176
rect 3442 14111 3762 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 13437 14176 13757 14177
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 14111 13757 14112
rect 5941 13632 6261 13633
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 13567 6261 13568
rect 10938 13632 11258 13633
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11258 13632
rect 10938 13567 11258 13568
rect 3442 13088 3762 13089
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3762 13088
rect 3442 13023 3762 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 13437 13088 13757 13089
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 13023 13757 13024
rect 5941 12544 6261 12545
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 12479 6261 12480
rect 10938 12544 11258 12545
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11258 12544
rect 10938 12479 11258 12480
rect 15653 12474 15719 12477
rect 16400 12474 17200 12504
rect 15653 12472 17200 12474
rect 15653 12416 15658 12472
rect 15714 12416 17200 12472
rect 15653 12414 17200 12416
rect 15653 12411 15719 12414
rect 16400 12384 17200 12414
rect 3442 12000 3762 12001
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3762 12000
rect 3442 11935 3762 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 13437 12000 13757 12001
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 11935 13757 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 5941 11456 6261 11457
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 11391 6261 11392
rect 10938 11456 11258 11457
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11258 11456
rect 10938 11391 11258 11392
rect 3442 10912 3762 10913
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3762 10912
rect 3442 10847 3762 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 13437 10912 13757 10913
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 10847 13757 10848
rect 5941 10368 6261 10369
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 10303 6261 10304
rect 10938 10368 11258 10369
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11258 10368
rect 10938 10303 11258 10304
rect 3442 9824 3762 9825
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3762 9824
rect 3442 9759 3762 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 13437 9824 13757 9825
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 9759 13757 9760
rect 5941 9280 6261 9281
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 9215 6261 9216
rect 10938 9280 11258 9281
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11258 9280
rect 10938 9215 11258 9216
rect 3442 8736 3762 8737
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3762 8736
rect 3442 8671 3762 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 13437 8736 13757 8737
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 8671 13757 8672
rect 0 8394 800 8424
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 5941 8192 6261 8193
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 8127 6261 8128
rect 10938 8192 11258 8193
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11258 8192
rect 10938 8127 11258 8128
rect 3442 7648 3762 7649
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3762 7648
rect 3442 7583 3762 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 13437 7648 13757 7649
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 7583 13757 7584
rect 13261 7442 13327 7445
rect 16400 7442 17200 7472
rect 13261 7440 17200 7442
rect 13261 7384 13266 7440
rect 13322 7384 17200 7440
rect 13261 7382 17200 7384
rect 13261 7379 13327 7382
rect 16400 7352 17200 7382
rect 5941 7104 6261 7105
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 7039 6261 7040
rect 10938 7104 11258 7105
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11258 7104
rect 10938 7039 11258 7040
rect 3442 6560 3762 6561
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3762 6560
rect 3442 6495 3762 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 13437 6560 13757 6561
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 6495 13757 6496
rect 5941 6016 6261 6017
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 5951 6261 5952
rect 10938 6016 11258 6017
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11258 6016
rect 10938 5951 11258 5952
rect 7925 5674 7991 5677
rect 9489 5674 9555 5677
rect 7925 5672 9555 5674
rect 7925 5616 7930 5672
rect 7986 5616 9494 5672
rect 9550 5616 9555 5672
rect 7925 5614 9555 5616
rect 7925 5611 7991 5614
rect 9489 5611 9555 5614
rect 3442 5472 3762 5473
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3762 5472
rect 3442 5407 3762 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 13437 5472 13757 5473
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 5407 13757 5408
rect 6729 5266 6795 5269
rect 9949 5266 10015 5269
rect 6729 5264 10015 5266
rect 6729 5208 6734 5264
rect 6790 5208 9954 5264
rect 10010 5208 10015 5264
rect 6729 5206 10015 5208
rect 6729 5203 6795 5206
rect 9949 5203 10015 5206
rect 5993 5130 6059 5133
rect 9489 5130 9555 5133
rect 5993 5128 9555 5130
rect 5993 5072 5998 5128
rect 6054 5072 9494 5128
rect 9550 5072 9555 5128
rect 5993 5070 9555 5072
rect 5993 5067 6059 5070
rect 9489 5067 9555 5070
rect 11789 5130 11855 5133
rect 12433 5130 12499 5133
rect 11789 5128 12499 5130
rect 11789 5072 11794 5128
rect 11850 5072 12438 5128
rect 12494 5072 12499 5128
rect 11789 5070 12499 5072
rect 11789 5067 11855 5070
rect 12433 5067 12499 5070
rect 0 4994 800 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 800 4934
rect 1485 4931 1551 4934
rect 5941 4928 6261 4929
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 4863 6261 4864
rect 10938 4928 11258 4929
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11258 4928
rect 10938 4863 11258 4864
rect 6821 4722 6887 4725
rect 9489 4722 9555 4725
rect 6821 4720 9555 4722
rect 6821 4664 6826 4720
rect 6882 4664 9494 4720
rect 9550 4664 9555 4720
rect 6821 4662 9555 4664
rect 6821 4659 6887 4662
rect 9489 4659 9555 4662
rect 3442 4384 3762 4385
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3762 4384
rect 3442 4319 3762 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 13437 4384 13757 4385
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 4319 13757 4320
rect 5941 3840 6261 3841
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 3775 6261 3776
rect 10938 3840 11258 3841
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11258 3840
rect 10938 3775 11258 3776
rect 3442 3296 3762 3297
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3762 3296
rect 3442 3231 3762 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 13437 3296 13757 3297
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 13437 3231 13757 3232
rect 5941 2752 6261 2753
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2687 6261 2688
rect 10938 2752 11258 2753
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11258 2752
rect 10938 2687 11258 2688
rect 15653 2546 15719 2549
rect 16400 2546 17200 2576
rect 15653 2544 17200 2546
rect 15653 2488 15658 2544
rect 15714 2488 17200 2544
rect 15653 2486 17200 2488
rect 15653 2483 15719 2486
rect 16400 2456 17200 2486
rect 3442 2208 3762 2209
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3762 2208
rect 3442 2143 3762 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 13437 2208 13757 2209
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2143 13757 2144
rect 0 1730 800 1760
rect 1669 1730 1735 1733
rect 0 1728 1735 1730
rect 0 1672 1674 1728
rect 1730 1672 1735 1728
rect 0 1670 1735 1672
rect 0 1640 800 1670
rect 1669 1667 1735 1670
<< via3 >>
rect 3450 17436 3514 17440
rect 3450 17380 3454 17436
rect 3454 17380 3510 17436
rect 3510 17380 3514 17436
rect 3450 17376 3514 17380
rect 3530 17436 3594 17440
rect 3530 17380 3534 17436
rect 3534 17380 3590 17436
rect 3590 17380 3594 17436
rect 3530 17376 3594 17380
rect 3610 17436 3674 17440
rect 3610 17380 3614 17436
rect 3614 17380 3670 17436
rect 3670 17380 3674 17436
rect 3610 17376 3674 17380
rect 3690 17436 3754 17440
rect 3690 17380 3694 17436
rect 3694 17380 3750 17436
rect 3750 17380 3754 17436
rect 3690 17376 3754 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 13445 17436 13509 17440
rect 13445 17380 13449 17436
rect 13449 17380 13505 17436
rect 13505 17380 13509 17436
rect 13445 17376 13509 17380
rect 13525 17436 13589 17440
rect 13525 17380 13529 17436
rect 13529 17380 13585 17436
rect 13585 17380 13589 17436
rect 13525 17376 13589 17380
rect 13605 17436 13669 17440
rect 13605 17380 13609 17436
rect 13609 17380 13665 17436
rect 13665 17380 13669 17436
rect 13605 17376 13669 17380
rect 13685 17436 13749 17440
rect 13685 17380 13689 17436
rect 13689 17380 13745 17436
rect 13745 17380 13749 17436
rect 13685 17376 13749 17380
rect 5949 16892 6013 16896
rect 5949 16836 5953 16892
rect 5953 16836 6009 16892
rect 6009 16836 6013 16892
rect 5949 16832 6013 16836
rect 6029 16892 6093 16896
rect 6029 16836 6033 16892
rect 6033 16836 6089 16892
rect 6089 16836 6093 16892
rect 6029 16832 6093 16836
rect 6109 16892 6173 16896
rect 6109 16836 6113 16892
rect 6113 16836 6169 16892
rect 6169 16836 6173 16892
rect 6109 16832 6173 16836
rect 6189 16892 6253 16896
rect 6189 16836 6193 16892
rect 6193 16836 6249 16892
rect 6249 16836 6253 16892
rect 6189 16832 6253 16836
rect 10946 16892 11010 16896
rect 10946 16836 10950 16892
rect 10950 16836 11006 16892
rect 11006 16836 11010 16892
rect 10946 16832 11010 16836
rect 11026 16892 11090 16896
rect 11026 16836 11030 16892
rect 11030 16836 11086 16892
rect 11086 16836 11090 16892
rect 11026 16832 11090 16836
rect 11106 16892 11170 16896
rect 11106 16836 11110 16892
rect 11110 16836 11166 16892
rect 11166 16836 11170 16892
rect 11106 16832 11170 16836
rect 11186 16892 11250 16896
rect 11186 16836 11190 16892
rect 11190 16836 11246 16892
rect 11246 16836 11250 16892
rect 11186 16832 11250 16836
rect 3450 16348 3514 16352
rect 3450 16292 3454 16348
rect 3454 16292 3510 16348
rect 3510 16292 3514 16348
rect 3450 16288 3514 16292
rect 3530 16348 3594 16352
rect 3530 16292 3534 16348
rect 3534 16292 3590 16348
rect 3590 16292 3594 16348
rect 3530 16288 3594 16292
rect 3610 16348 3674 16352
rect 3610 16292 3614 16348
rect 3614 16292 3670 16348
rect 3670 16292 3674 16348
rect 3610 16288 3674 16292
rect 3690 16348 3754 16352
rect 3690 16292 3694 16348
rect 3694 16292 3750 16348
rect 3750 16292 3754 16348
rect 3690 16288 3754 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 13445 16348 13509 16352
rect 13445 16292 13449 16348
rect 13449 16292 13505 16348
rect 13505 16292 13509 16348
rect 13445 16288 13509 16292
rect 13525 16348 13589 16352
rect 13525 16292 13529 16348
rect 13529 16292 13585 16348
rect 13585 16292 13589 16348
rect 13525 16288 13589 16292
rect 13605 16348 13669 16352
rect 13605 16292 13609 16348
rect 13609 16292 13665 16348
rect 13665 16292 13669 16348
rect 13605 16288 13669 16292
rect 13685 16348 13749 16352
rect 13685 16292 13689 16348
rect 13689 16292 13745 16348
rect 13745 16292 13749 16348
rect 13685 16288 13749 16292
rect 5949 15804 6013 15808
rect 5949 15748 5953 15804
rect 5953 15748 6009 15804
rect 6009 15748 6013 15804
rect 5949 15744 6013 15748
rect 6029 15804 6093 15808
rect 6029 15748 6033 15804
rect 6033 15748 6089 15804
rect 6089 15748 6093 15804
rect 6029 15744 6093 15748
rect 6109 15804 6173 15808
rect 6109 15748 6113 15804
rect 6113 15748 6169 15804
rect 6169 15748 6173 15804
rect 6109 15744 6173 15748
rect 6189 15804 6253 15808
rect 6189 15748 6193 15804
rect 6193 15748 6249 15804
rect 6249 15748 6253 15804
rect 6189 15744 6253 15748
rect 10946 15804 11010 15808
rect 10946 15748 10950 15804
rect 10950 15748 11006 15804
rect 11006 15748 11010 15804
rect 10946 15744 11010 15748
rect 11026 15804 11090 15808
rect 11026 15748 11030 15804
rect 11030 15748 11086 15804
rect 11086 15748 11090 15804
rect 11026 15744 11090 15748
rect 11106 15804 11170 15808
rect 11106 15748 11110 15804
rect 11110 15748 11166 15804
rect 11166 15748 11170 15804
rect 11106 15744 11170 15748
rect 11186 15804 11250 15808
rect 11186 15748 11190 15804
rect 11190 15748 11246 15804
rect 11246 15748 11250 15804
rect 11186 15744 11250 15748
rect 3450 15260 3514 15264
rect 3450 15204 3454 15260
rect 3454 15204 3510 15260
rect 3510 15204 3514 15260
rect 3450 15200 3514 15204
rect 3530 15260 3594 15264
rect 3530 15204 3534 15260
rect 3534 15204 3590 15260
rect 3590 15204 3594 15260
rect 3530 15200 3594 15204
rect 3610 15260 3674 15264
rect 3610 15204 3614 15260
rect 3614 15204 3670 15260
rect 3670 15204 3674 15260
rect 3610 15200 3674 15204
rect 3690 15260 3754 15264
rect 3690 15204 3694 15260
rect 3694 15204 3750 15260
rect 3750 15204 3754 15260
rect 3690 15200 3754 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 13445 15260 13509 15264
rect 13445 15204 13449 15260
rect 13449 15204 13505 15260
rect 13505 15204 13509 15260
rect 13445 15200 13509 15204
rect 13525 15260 13589 15264
rect 13525 15204 13529 15260
rect 13529 15204 13585 15260
rect 13585 15204 13589 15260
rect 13525 15200 13589 15204
rect 13605 15260 13669 15264
rect 13605 15204 13609 15260
rect 13609 15204 13665 15260
rect 13665 15204 13669 15260
rect 13605 15200 13669 15204
rect 13685 15260 13749 15264
rect 13685 15204 13689 15260
rect 13689 15204 13745 15260
rect 13745 15204 13749 15260
rect 13685 15200 13749 15204
rect 5949 14716 6013 14720
rect 5949 14660 5953 14716
rect 5953 14660 6009 14716
rect 6009 14660 6013 14716
rect 5949 14656 6013 14660
rect 6029 14716 6093 14720
rect 6029 14660 6033 14716
rect 6033 14660 6089 14716
rect 6089 14660 6093 14716
rect 6029 14656 6093 14660
rect 6109 14716 6173 14720
rect 6109 14660 6113 14716
rect 6113 14660 6169 14716
rect 6169 14660 6173 14716
rect 6109 14656 6173 14660
rect 6189 14716 6253 14720
rect 6189 14660 6193 14716
rect 6193 14660 6249 14716
rect 6249 14660 6253 14716
rect 6189 14656 6253 14660
rect 10946 14716 11010 14720
rect 10946 14660 10950 14716
rect 10950 14660 11006 14716
rect 11006 14660 11010 14716
rect 10946 14656 11010 14660
rect 11026 14716 11090 14720
rect 11026 14660 11030 14716
rect 11030 14660 11086 14716
rect 11086 14660 11090 14716
rect 11026 14656 11090 14660
rect 11106 14716 11170 14720
rect 11106 14660 11110 14716
rect 11110 14660 11166 14716
rect 11166 14660 11170 14716
rect 11106 14656 11170 14660
rect 11186 14716 11250 14720
rect 11186 14660 11190 14716
rect 11190 14660 11246 14716
rect 11246 14660 11250 14716
rect 11186 14656 11250 14660
rect 3450 14172 3514 14176
rect 3450 14116 3454 14172
rect 3454 14116 3510 14172
rect 3510 14116 3514 14172
rect 3450 14112 3514 14116
rect 3530 14172 3594 14176
rect 3530 14116 3534 14172
rect 3534 14116 3590 14172
rect 3590 14116 3594 14172
rect 3530 14112 3594 14116
rect 3610 14172 3674 14176
rect 3610 14116 3614 14172
rect 3614 14116 3670 14172
rect 3670 14116 3674 14172
rect 3610 14112 3674 14116
rect 3690 14172 3754 14176
rect 3690 14116 3694 14172
rect 3694 14116 3750 14172
rect 3750 14116 3754 14172
rect 3690 14112 3754 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 13445 14172 13509 14176
rect 13445 14116 13449 14172
rect 13449 14116 13505 14172
rect 13505 14116 13509 14172
rect 13445 14112 13509 14116
rect 13525 14172 13589 14176
rect 13525 14116 13529 14172
rect 13529 14116 13585 14172
rect 13585 14116 13589 14172
rect 13525 14112 13589 14116
rect 13605 14172 13669 14176
rect 13605 14116 13609 14172
rect 13609 14116 13665 14172
rect 13665 14116 13669 14172
rect 13605 14112 13669 14116
rect 13685 14172 13749 14176
rect 13685 14116 13689 14172
rect 13689 14116 13745 14172
rect 13745 14116 13749 14172
rect 13685 14112 13749 14116
rect 5949 13628 6013 13632
rect 5949 13572 5953 13628
rect 5953 13572 6009 13628
rect 6009 13572 6013 13628
rect 5949 13568 6013 13572
rect 6029 13628 6093 13632
rect 6029 13572 6033 13628
rect 6033 13572 6089 13628
rect 6089 13572 6093 13628
rect 6029 13568 6093 13572
rect 6109 13628 6173 13632
rect 6109 13572 6113 13628
rect 6113 13572 6169 13628
rect 6169 13572 6173 13628
rect 6109 13568 6173 13572
rect 6189 13628 6253 13632
rect 6189 13572 6193 13628
rect 6193 13572 6249 13628
rect 6249 13572 6253 13628
rect 6189 13568 6253 13572
rect 10946 13628 11010 13632
rect 10946 13572 10950 13628
rect 10950 13572 11006 13628
rect 11006 13572 11010 13628
rect 10946 13568 11010 13572
rect 11026 13628 11090 13632
rect 11026 13572 11030 13628
rect 11030 13572 11086 13628
rect 11086 13572 11090 13628
rect 11026 13568 11090 13572
rect 11106 13628 11170 13632
rect 11106 13572 11110 13628
rect 11110 13572 11166 13628
rect 11166 13572 11170 13628
rect 11106 13568 11170 13572
rect 11186 13628 11250 13632
rect 11186 13572 11190 13628
rect 11190 13572 11246 13628
rect 11246 13572 11250 13628
rect 11186 13568 11250 13572
rect 3450 13084 3514 13088
rect 3450 13028 3454 13084
rect 3454 13028 3510 13084
rect 3510 13028 3514 13084
rect 3450 13024 3514 13028
rect 3530 13084 3594 13088
rect 3530 13028 3534 13084
rect 3534 13028 3590 13084
rect 3590 13028 3594 13084
rect 3530 13024 3594 13028
rect 3610 13084 3674 13088
rect 3610 13028 3614 13084
rect 3614 13028 3670 13084
rect 3670 13028 3674 13084
rect 3610 13024 3674 13028
rect 3690 13084 3754 13088
rect 3690 13028 3694 13084
rect 3694 13028 3750 13084
rect 3750 13028 3754 13084
rect 3690 13024 3754 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 13445 13084 13509 13088
rect 13445 13028 13449 13084
rect 13449 13028 13505 13084
rect 13505 13028 13509 13084
rect 13445 13024 13509 13028
rect 13525 13084 13589 13088
rect 13525 13028 13529 13084
rect 13529 13028 13585 13084
rect 13585 13028 13589 13084
rect 13525 13024 13589 13028
rect 13605 13084 13669 13088
rect 13605 13028 13609 13084
rect 13609 13028 13665 13084
rect 13665 13028 13669 13084
rect 13605 13024 13669 13028
rect 13685 13084 13749 13088
rect 13685 13028 13689 13084
rect 13689 13028 13745 13084
rect 13745 13028 13749 13084
rect 13685 13024 13749 13028
rect 5949 12540 6013 12544
rect 5949 12484 5953 12540
rect 5953 12484 6009 12540
rect 6009 12484 6013 12540
rect 5949 12480 6013 12484
rect 6029 12540 6093 12544
rect 6029 12484 6033 12540
rect 6033 12484 6089 12540
rect 6089 12484 6093 12540
rect 6029 12480 6093 12484
rect 6109 12540 6173 12544
rect 6109 12484 6113 12540
rect 6113 12484 6169 12540
rect 6169 12484 6173 12540
rect 6109 12480 6173 12484
rect 6189 12540 6253 12544
rect 6189 12484 6193 12540
rect 6193 12484 6249 12540
rect 6249 12484 6253 12540
rect 6189 12480 6253 12484
rect 10946 12540 11010 12544
rect 10946 12484 10950 12540
rect 10950 12484 11006 12540
rect 11006 12484 11010 12540
rect 10946 12480 11010 12484
rect 11026 12540 11090 12544
rect 11026 12484 11030 12540
rect 11030 12484 11086 12540
rect 11086 12484 11090 12540
rect 11026 12480 11090 12484
rect 11106 12540 11170 12544
rect 11106 12484 11110 12540
rect 11110 12484 11166 12540
rect 11166 12484 11170 12540
rect 11106 12480 11170 12484
rect 11186 12540 11250 12544
rect 11186 12484 11190 12540
rect 11190 12484 11246 12540
rect 11246 12484 11250 12540
rect 11186 12480 11250 12484
rect 3450 11996 3514 12000
rect 3450 11940 3454 11996
rect 3454 11940 3510 11996
rect 3510 11940 3514 11996
rect 3450 11936 3514 11940
rect 3530 11996 3594 12000
rect 3530 11940 3534 11996
rect 3534 11940 3590 11996
rect 3590 11940 3594 11996
rect 3530 11936 3594 11940
rect 3610 11996 3674 12000
rect 3610 11940 3614 11996
rect 3614 11940 3670 11996
rect 3670 11940 3674 11996
rect 3610 11936 3674 11940
rect 3690 11996 3754 12000
rect 3690 11940 3694 11996
rect 3694 11940 3750 11996
rect 3750 11940 3754 11996
rect 3690 11936 3754 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 13445 11996 13509 12000
rect 13445 11940 13449 11996
rect 13449 11940 13505 11996
rect 13505 11940 13509 11996
rect 13445 11936 13509 11940
rect 13525 11996 13589 12000
rect 13525 11940 13529 11996
rect 13529 11940 13585 11996
rect 13585 11940 13589 11996
rect 13525 11936 13589 11940
rect 13605 11996 13669 12000
rect 13605 11940 13609 11996
rect 13609 11940 13665 11996
rect 13665 11940 13669 11996
rect 13605 11936 13669 11940
rect 13685 11996 13749 12000
rect 13685 11940 13689 11996
rect 13689 11940 13745 11996
rect 13745 11940 13749 11996
rect 13685 11936 13749 11940
rect 5949 11452 6013 11456
rect 5949 11396 5953 11452
rect 5953 11396 6009 11452
rect 6009 11396 6013 11452
rect 5949 11392 6013 11396
rect 6029 11452 6093 11456
rect 6029 11396 6033 11452
rect 6033 11396 6089 11452
rect 6089 11396 6093 11452
rect 6029 11392 6093 11396
rect 6109 11452 6173 11456
rect 6109 11396 6113 11452
rect 6113 11396 6169 11452
rect 6169 11396 6173 11452
rect 6109 11392 6173 11396
rect 6189 11452 6253 11456
rect 6189 11396 6193 11452
rect 6193 11396 6249 11452
rect 6249 11396 6253 11452
rect 6189 11392 6253 11396
rect 10946 11452 11010 11456
rect 10946 11396 10950 11452
rect 10950 11396 11006 11452
rect 11006 11396 11010 11452
rect 10946 11392 11010 11396
rect 11026 11452 11090 11456
rect 11026 11396 11030 11452
rect 11030 11396 11086 11452
rect 11086 11396 11090 11452
rect 11026 11392 11090 11396
rect 11106 11452 11170 11456
rect 11106 11396 11110 11452
rect 11110 11396 11166 11452
rect 11166 11396 11170 11452
rect 11106 11392 11170 11396
rect 11186 11452 11250 11456
rect 11186 11396 11190 11452
rect 11190 11396 11246 11452
rect 11246 11396 11250 11452
rect 11186 11392 11250 11396
rect 3450 10908 3514 10912
rect 3450 10852 3454 10908
rect 3454 10852 3510 10908
rect 3510 10852 3514 10908
rect 3450 10848 3514 10852
rect 3530 10908 3594 10912
rect 3530 10852 3534 10908
rect 3534 10852 3590 10908
rect 3590 10852 3594 10908
rect 3530 10848 3594 10852
rect 3610 10908 3674 10912
rect 3610 10852 3614 10908
rect 3614 10852 3670 10908
rect 3670 10852 3674 10908
rect 3610 10848 3674 10852
rect 3690 10908 3754 10912
rect 3690 10852 3694 10908
rect 3694 10852 3750 10908
rect 3750 10852 3754 10908
rect 3690 10848 3754 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 13445 10908 13509 10912
rect 13445 10852 13449 10908
rect 13449 10852 13505 10908
rect 13505 10852 13509 10908
rect 13445 10848 13509 10852
rect 13525 10908 13589 10912
rect 13525 10852 13529 10908
rect 13529 10852 13585 10908
rect 13585 10852 13589 10908
rect 13525 10848 13589 10852
rect 13605 10908 13669 10912
rect 13605 10852 13609 10908
rect 13609 10852 13665 10908
rect 13665 10852 13669 10908
rect 13605 10848 13669 10852
rect 13685 10908 13749 10912
rect 13685 10852 13689 10908
rect 13689 10852 13745 10908
rect 13745 10852 13749 10908
rect 13685 10848 13749 10852
rect 5949 10364 6013 10368
rect 5949 10308 5953 10364
rect 5953 10308 6009 10364
rect 6009 10308 6013 10364
rect 5949 10304 6013 10308
rect 6029 10364 6093 10368
rect 6029 10308 6033 10364
rect 6033 10308 6089 10364
rect 6089 10308 6093 10364
rect 6029 10304 6093 10308
rect 6109 10364 6173 10368
rect 6109 10308 6113 10364
rect 6113 10308 6169 10364
rect 6169 10308 6173 10364
rect 6109 10304 6173 10308
rect 6189 10364 6253 10368
rect 6189 10308 6193 10364
rect 6193 10308 6249 10364
rect 6249 10308 6253 10364
rect 6189 10304 6253 10308
rect 10946 10364 11010 10368
rect 10946 10308 10950 10364
rect 10950 10308 11006 10364
rect 11006 10308 11010 10364
rect 10946 10304 11010 10308
rect 11026 10364 11090 10368
rect 11026 10308 11030 10364
rect 11030 10308 11086 10364
rect 11086 10308 11090 10364
rect 11026 10304 11090 10308
rect 11106 10364 11170 10368
rect 11106 10308 11110 10364
rect 11110 10308 11166 10364
rect 11166 10308 11170 10364
rect 11106 10304 11170 10308
rect 11186 10364 11250 10368
rect 11186 10308 11190 10364
rect 11190 10308 11246 10364
rect 11246 10308 11250 10364
rect 11186 10304 11250 10308
rect 3450 9820 3514 9824
rect 3450 9764 3454 9820
rect 3454 9764 3510 9820
rect 3510 9764 3514 9820
rect 3450 9760 3514 9764
rect 3530 9820 3594 9824
rect 3530 9764 3534 9820
rect 3534 9764 3590 9820
rect 3590 9764 3594 9820
rect 3530 9760 3594 9764
rect 3610 9820 3674 9824
rect 3610 9764 3614 9820
rect 3614 9764 3670 9820
rect 3670 9764 3674 9820
rect 3610 9760 3674 9764
rect 3690 9820 3754 9824
rect 3690 9764 3694 9820
rect 3694 9764 3750 9820
rect 3750 9764 3754 9820
rect 3690 9760 3754 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 13445 9820 13509 9824
rect 13445 9764 13449 9820
rect 13449 9764 13505 9820
rect 13505 9764 13509 9820
rect 13445 9760 13509 9764
rect 13525 9820 13589 9824
rect 13525 9764 13529 9820
rect 13529 9764 13585 9820
rect 13585 9764 13589 9820
rect 13525 9760 13589 9764
rect 13605 9820 13669 9824
rect 13605 9764 13609 9820
rect 13609 9764 13665 9820
rect 13665 9764 13669 9820
rect 13605 9760 13669 9764
rect 13685 9820 13749 9824
rect 13685 9764 13689 9820
rect 13689 9764 13745 9820
rect 13745 9764 13749 9820
rect 13685 9760 13749 9764
rect 5949 9276 6013 9280
rect 5949 9220 5953 9276
rect 5953 9220 6009 9276
rect 6009 9220 6013 9276
rect 5949 9216 6013 9220
rect 6029 9276 6093 9280
rect 6029 9220 6033 9276
rect 6033 9220 6089 9276
rect 6089 9220 6093 9276
rect 6029 9216 6093 9220
rect 6109 9276 6173 9280
rect 6109 9220 6113 9276
rect 6113 9220 6169 9276
rect 6169 9220 6173 9276
rect 6109 9216 6173 9220
rect 6189 9276 6253 9280
rect 6189 9220 6193 9276
rect 6193 9220 6249 9276
rect 6249 9220 6253 9276
rect 6189 9216 6253 9220
rect 10946 9276 11010 9280
rect 10946 9220 10950 9276
rect 10950 9220 11006 9276
rect 11006 9220 11010 9276
rect 10946 9216 11010 9220
rect 11026 9276 11090 9280
rect 11026 9220 11030 9276
rect 11030 9220 11086 9276
rect 11086 9220 11090 9276
rect 11026 9216 11090 9220
rect 11106 9276 11170 9280
rect 11106 9220 11110 9276
rect 11110 9220 11166 9276
rect 11166 9220 11170 9276
rect 11106 9216 11170 9220
rect 11186 9276 11250 9280
rect 11186 9220 11190 9276
rect 11190 9220 11246 9276
rect 11246 9220 11250 9276
rect 11186 9216 11250 9220
rect 3450 8732 3514 8736
rect 3450 8676 3454 8732
rect 3454 8676 3510 8732
rect 3510 8676 3514 8732
rect 3450 8672 3514 8676
rect 3530 8732 3594 8736
rect 3530 8676 3534 8732
rect 3534 8676 3590 8732
rect 3590 8676 3594 8732
rect 3530 8672 3594 8676
rect 3610 8732 3674 8736
rect 3610 8676 3614 8732
rect 3614 8676 3670 8732
rect 3670 8676 3674 8732
rect 3610 8672 3674 8676
rect 3690 8732 3754 8736
rect 3690 8676 3694 8732
rect 3694 8676 3750 8732
rect 3750 8676 3754 8732
rect 3690 8672 3754 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 13445 8732 13509 8736
rect 13445 8676 13449 8732
rect 13449 8676 13505 8732
rect 13505 8676 13509 8732
rect 13445 8672 13509 8676
rect 13525 8732 13589 8736
rect 13525 8676 13529 8732
rect 13529 8676 13585 8732
rect 13585 8676 13589 8732
rect 13525 8672 13589 8676
rect 13605 8732 13669 8736
rect 13605 8676 13609 8732
rect 13609 8676 13665 8732
rect 13665 8676 13669 8732
rect 13605 8672 13669 8676
rect 13685 8732 13749 8736
rect 13685 8676 13689 8732
rect 13689 8676 13745 8732
rect 13745 8676 13749 8732
rect 13685 8672 13749 8676
rect 5949 8188 6013 8192
rect 5949 8132 5953 8188
rect 5953 8132 6009 8188
rect 6009 8132 6013 8188
rect 5949 8128 6013 8132
rect 6029 8188 6093 8192
rect 6029 8132 6033 8188
rect 6033 8132 6089 8188
rect 6089 8132 6093 8188
rect 6029 8128 6093 8132
rect 6109 8188 6173 8192
rect 6109 8132 6113 8188
rect 6113 8132 6169 8188
rect 6169 8132 6173 8188
rect 6109 8128 6173 8132
rect 6189 8188 6253 8192
rect 6189 8132 6193 8188
rect 6193 8132 6249 8188
rect 6249 8132 6253 8188
rect 6189 8128 6253 8132
rect 10946 8188 11010 8192
rect 10946 8132 10950 8188
rect 10950 8132 11006 8188
rect 11006 8132 11010 8188
rect 10946 8128 11010 8132
rect 11026 8188 11090 8192
rect 11026 8132 11030 8188
rect 11030 8132 11086 8188
rect 11086 8132 11090 8188
rect 11026 8128 11090 8132
rect 11106 8188 11170 8192
rect 11106 8132 11110 8188
rect 11110 8132 11166 8188
rect 11166 8132 11170 8188
rect 11106 8128 11170 8132
rect 11186 8188 11250 8192
rect 11186 8132 11190 8188
rect 11190 8132 11246 8188
rect 11246 8132 11250 8188
rect 11186 8128 11250 8132
rect 3450 7644 3514 7648
rect 3450 7588 3454 7644
rect 3454 7588 3510 7644
rect 3510 7588 3514 7644
rect 3450 7584 3514 7588
rect 3530 7644 3594 7648
rect 3530 7588 3534 7644
rect 3534 7588 3590 7644
rect 3590 7588 3594 7644
rect 3530 7584 3594 7588
rect 3610 7644 3674 7648
rect 3610 7588 3614 7644
rect 3614 7588 3670 7644
rect 3670 7588 3674 7644
rect 3610 7584 3674 7588
rect 3690 7644 3754 7648
rect 3690 7588 3694 7644
rect 3694 7588 3750 7644
rect 3750 7588 3754 7644
rect 3690 7584 3754 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 13445 7644 13509 7648
rect 13445 7588 13449 7644
rect 13449 7588 13505 7644
rect 13505 7588 13509 7644
rect 13445 7584 13509 7588
rect 13525 7644 13589 7648
rect 13525 7588 13529 7644
rect 13529 7588 13585 7644
rect 13585 7588 13589 7644
rect 13525 7584 13589 7588
rect 13605 7644 13669 7648
rect 13605 7588 13609 7644
rect 13609 7588 13665 7644
rect 13665 7588 13669 7644
rect 13605 7584 13669 7588
rect 13685 7644 13749 7648
rect 13685 7588 13689 7644
rect 13689 7588 13745 7644
rect 13745 7588 13749 7644
rect 13685 7584 13749 7588
rect 5949 7100 6013 7104
rect 5949 7044 5953 7100
rect 5953 7044 6009 7100
rect 6009 7044 6013 7100
rect 5949 7040 6013 7044
rect 6029 7100 6093 7104
rect 6029 7044 6033 7100
rect 6033 7044 6089 7100
rect 6089 7044 6093 7100
rect 6029 7040 6093 7044
rect 6109 7100 6173 7104
rect 6109 7044 6113 7100
rect 6113 7044 6169 7100
rect 6169 7044 6173 7100
rect 6109 7040 6173 7044
rect 6189 7100 6253 7104
rect 6189 7044 6193 7100
rect 6193 7044 6249 7100
rect 6249 7044 6253 7100
rect 6189 7040 6253 7044
rect 10946 7100 11010 7104
rect 10946 7044 10950 7100
rect 10950 7044 11006 7100
rect 11006 7044 11010 7100
rect 10946 7040 11010 7044
rect 11026 7100 11090 7104
rect 11026 7044 11030 7100
rect 11030 7044 11086 7100
rect 11086 7044 11090 7100
rect 11026 7040 11090 7044
rect 11106 7100 11170 7104
rect 11106 7044 11110 7100
rect 11110 7044 11166 7100
rect 11166 7044 11170 7100
rect 11106 7040 11170 7044
rect 11186 7100 11250 7104
rect 11186 7044 11190 7100
rect 11190 7044 11246 7100
rect 11246 7044 11250 7100
rect 11186 7040 11250 7044
rect 3450 6556 3514 6560
rect 3450 6500 3454 6556
rect 3454 6500 3510 6556
rect 3510 6500 3514 6556
rect 3450 6496 3514 6500
rect 3530 6556 3594 6560
rect 3530 6500 3534 6556
rect 3534 6500 3590 6556
rect 3590 6500 3594 6556
rect 3530 6496 3594 6500
rect 3610 6556 3674 6560
rect 3610 6500 3614 6556
rect 3614 6500 3670 6556
rect 3670 6500 3674 6556
rect 3610 6496 3674 6500
rect 3690 6556 3754 6560
rect 3690 6500 3694 6556
rect 3694 6500 3750 6556
rect 3750 6500 3754 6556
rect 3690 6496 3754 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 13445 6556 13509 6560
rect 13445 6500 13449 6556
rect 13449 6500 13505 6556
rect 13505 6500 13509 6556
rect 13445 6496 13509 6500
rect 13525 6556 13589 6560
rect 13525 6500 13529 6556
rect 13529 6500 13585 6556
rect 13585 6500 13589 6556
rect 13525 6496 13589 6500
rect 13605 6556 13669 6560
rect 13605 6500 13609 6556
rect 13609 6500 13665 6556
rect 13665 6500 13669 6556
rect 13605 6496 13669 6500
rect 13685 6556 13749 6560
rect 13685 6500 13689 6556
rect 13689 6500 13745 6556
rect 13745 6500 13749 6556
rect 13685 6496 13749 6500
rect 5949 6012 6013 6016
rect 5949 5956 5953 6012
rect 5953 5956 6009 6012
rect 6009 5956 6013 6012
rect 5949 5952 6013 5956
rect 6029 6012 6093 6016
rect 6029 5956 6033 6012
rect 6033 5956 6089 6012
rect 6089 5956 6093 6012
rect 6029 5952 6093 5956
rect 6109 6012 6173 6016
rect 6109 5956 6113 6012
rect 6113 5956 6169 6012
rect 6169 5956 6173 6012
rect 6109 5952 6173 5956
rect 6189 6012 6253 6016
rect 6189 5956 6193 6012
rect 6193 5956 6249 6012
rect 6249 5956 6253 6012
rect 6189 5952 6253 5956
rect 10946 6012 11010 6016
rect 10946 5956 10950 6012
rect 10950 5956 11006 6012
rect 11006 5956 11010 6012
rect 10946 5952 11010 5956
rect 11026 6012 11090 6016
rect 11026 5956 11030 6012
rect 11030 5956 11086 6012
rect 11086 5956 11090 6012
rect 11026 5952 11090 5956
rect 11106 6012 11170 6016
rect 11106 5956 11110 6012
rect 11110 5956 11166 6012
rect 11166 5956 11170 6012
rect 11106 5952 11170 5956
rect 11186 6012 11250 6016
rect 11186 5956 11190 6012
rect 11190 5956 11246 6012
rect 11246 5956 11250 6012
rect 11186 5952 11250 5956
rect 3450 5468 3514 5472
rect 3450 5412 3454 5468
rect 3454 5412 3510 5468
rect 3510 5412 3514 5468
rect 3450 5408 3514 5412
rect 3530 5468 3594 5472
rect 3530 5412 3534 5468
rect 3534 5412 3590 5468
rect 3590 5412 3594 5468
rect 3530 5408 3594 5412
rect 3610 5468 3674 5472
rect 3610 5412 3614 5468
rect 3614 5412 3670 5468
rect 3670 5412 3674 5468
rect 3610 5408 3674 5412
rect 3690 5468 3754 5472
rect 3690 5412 3694 5468
rect 3694 5412 3750 5468
rect 3750 5412 3754 5468
rect 3690 5408 3754 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 13445 5468 13509 5472
rect 13445 5412 13449 5468
rect 13449 5412 13505 5468
rect 13505 5412 13509 5468
rect 13445 5408 13509 5412
rect 13525 5468 13589 5472
rect 13525 5412 13529 5468
rect 13529 5412 13585 5468
rect 13585 5412 13589 5468
rect 13525 5408 13589 5412
rect 13605 5468 13669 5472
rect 13605 5412 13609 5468
rect 13609 5412 13665 5468
rect 13665 5412 13669 5468
rect 13605 5408 13669 5412
rect 13685 5468 13749 5472
rect 13685 5412 13689 5468
rect 13689 5412 13745 5468
rect 13745 5412 13749 5468
rect 13685 5408 13749 5412
rect 5949 4924 6013 4928
rect 5949 4868 5953 4924
rect 5953 4868 6009 4924
rect 6009 4868 6013 4924
rect 5949 4864 6013 4868
rect 6029 4924 6093 4928
rect 6029 4868 6033 4924
rect 6033 4868 6089 4924
rect 6089 4868 6093 4924
rect 6029 4864 6093 4868
rect 6109 4924 6173 4928
rect 6109 4868 6113 4924
rect 6113 4868 6169 4924
rect 6169 4868 6173 4924
rect 6109 4864 6173 4868
rect 6189 4924 6253 4928
rect 6189 4868 6193 4924
rect 6193 4868 6249 4924
rect 6249 4868 6253 4924
rect 6189 4864 6253 4868
rect 10946 4924 11010 4928
rect 10946 4868 10950 4924
rect 10950 4868 11006 4924
rect 11006 4868 11010 4924
rect 10946 4864 11010 4868
rect 11026 4924 11090 4928
rect 11026 4868 11030 4924
rect 11030 4868 11086 4924
rect 11086 4868 11090 4924
rect 11026 4864 11090 4868
rect 11106 4924 11170 4928
rect 11106 4868 11110 4924
rect 11110 4868 11166 4924
rect 11166 4868 11170 4924
rect 11106 4864 11170 4868
rect 11186 4924 11250 4928
rect 11186 4868 11190 4924
rect 11190 4868 11246 4924
rect 11246 4868 11250 4924
rect 11186 4864 11250 4868
rect 3450 4380 3514 4384
rect 3450 4324 3454 4380
rect 3454 4324 3510 4380
rect 3510 4324 3514 4380
rect 3450 4320 3514 4324
rect 3530 4380 3594 4384
rect 3530 4324 3534 4380
rect 3534 4324 3590 4380
rect 3590 4324 3594 4380
rect 3530 4320 3594 4324
rect 3610 4380 3674 4384
rect 3610 4324 3614 4380
rect 3614 4324 3670 4380
rect 3670 4324 3674 4380
rect 3610 4320 3674 4324
rect 3690 4380 3754 4384
rect 3690 4324 3694 4380
rect 3694 4324 3750 4380
rect 3750 4324 3754 4380
rect 3690 4320 3754 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 13445 4380 13509 4384
rect 13445 4324 13449 4380
rect 13449 4324 13505 4380
rect 13505 4324 13509 4380
rect 13445 4320 13509 4324
rect 13525 4380 13589 4384
rect 13525 4324 13529 4380
rect 13529 4324 13585 4380
rect 13585 4324 13589 4380
rect 13525 4320 13589 4324
rect 13605 4380 13669 4384
rect 13605 4324 13609 4380
rect 13609 4324 13665 4380
rect 13665 4324 13669 4380
rect 13605 4320 13669 4324
rect 13685 4380 13749 4384
rect 13685 4324 13689 4380
rect 13689 4324 13745 4380
rect 13745 4324 13749 4380
rect 13685 4320 13749 4324
rect 5949 3836 6013 3840
rect 5949 3780 5953 3836
rect 5953 3780 6009 3836
rect 6009 3780 6013 3836
rect 5949 3776 6013 3780
rect 6029 3836 6093 3840
rect 6029 3780 6033 3836
rect 6033 3780 6089 3836
rect 6089 3780 6093 3836
rect 6029 3776 6093 3780
rect 6109 3836 6173 3840
rect 6109 3780 6113 3836
rect 6113 3780 6169 3836
rect 6169 3780 6173 3836
rect 6109 3776 6173 3780
rect 6189 3836 6253 3840
rect 6189 3780 6193 3836
rect 6193 3780 6249 3836
rect 6249 3780 6253 3836
rect 6189 3776 6253 3780
rect 10946 3836 11010 3840
rect 10946 3780 10950 3836
rect 10950 3780 11006 3836
rect 11006 3780 11010 3836
rect 10946 3776 11010 3780
rect 11026 3836 11090 3840
rect 11026 3780 11030 3836
rect 11030 3780 11086 3836
rect 11086 3780 11090 3836
rect 11026 3776 11090 3780
rect 11106 3836 11170 3840
rect 11106 3780 11110 3836
rect 11110 3780 11166 3836
rect 11166 3780 11170 3836
rect 11106 3776 11170 3780
rect 11186 3836 11250 3840
rect 11186 3780 11190 3836
rect 11190 3780 11246 3836
rect 11246 3780 11250 3836
rect 11186 3776 11250 3780
rect 3450 3292 3514 3296
rect 3450 3236 3454 3292
rect 3454 3236 3510 3292
rect 3510 3236 3514 3292
rect 3450 3232 3514 3236
rect 3530 3292 3594 3296
rect 3530 3236 3534 3292
rect 3534 3236 3590 3292
rect 3590 3236 3594 3292
rect 3530 3232 3594 3236
rect 3610 3292 3674 3296
rect 3610 3236 3614 3292
rect 3614 3236 3670 3292
rect 3670 3236 3674 3292
rect 3610 3232 3674 3236
rect 3690 3292 3754 3296
rect 3690 3236 3694 3292
rect 3694 3236 3750 3292
rect 3750 3236 3754 3292
rect 3690 3232 3754 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 13445 3292 13509 3296
rect 13445 3236 13449 3292
rect 13449 3236 13505 3292
rect 13505 3236 13509 3292
rect 13445 3232 13509 3236
rect 13525 3292 13589 3296
rect 13525 3236 13529 3292
rect 13529 3236 13585 3292
rect 13585 3236 13589 3292
rect 13525 3232 13589 3236
rect 13605 3292 13669 3296
rect 13605 3236 13609 3292
rect 13609 3236 13665 3292
rect 13665 3236 13669 3292
rect 13605 3232 13669 3236
rect 13685 3292 13749 3296
rect 13685 3236 13689 3292
rect 13689 3236 13745 3292
rect 13745 3236 13749 3292
rect 13685 3232 13749 3236
rect 5949 2748 6013 2752
rect 5949 2692 5953 2748
rect 5953 2692 6009 2748
rect 6009 2692 6013 2748
rect 5949 2688 6013 2692
rect 6029 2748 6093 2752
rect 6029 2692 6033 2748
rect 6033 2692 6089 2748
rect 6089 2692 6093 2748
rect 6029 2688 6093 2692
rect 6109 2748 6173 2752
rect 6109 2692 6113 2748
rect 6113 2692 6169 2748
rect 6169 2692 6173 2748
rect 6109 2688 6173 2692
rect 6189 2748 6253 2752
rect 6189 2692 6193 2748
rect 6193 2692 6249 2748
rect 6249 2692 6253 2748
rect 6189 2688 6253 2692
rect 10946 2748 11010 2752
rect 10946 2692 10950 2748
rect 10950 2692 11006 2748
rect 11006 2692 11010 2748
rect 10946 2688 11010 2692
rect 11026 2748 11090 2752
rect 11026 2692 11030 2748
rect 11030 2692 11086 2748
rect 11086 2692 11090 2748
rect 11026 2688 11090 2692
rect 11106 2748 11170 2752
rect 11106 2692 11110 2748
rect 11110 2692 11166 2748
rect 11166 2692 11170 2748
rect 11106 2688 11170 2692
rect 11186 2748 11250 2752
rect 11186 2692 11190 2748
rect 11190 2692 11246 2748
rect 11246 2692 11250 2748
rect 11186 2688 11250 2692
rect 3450 2204 3514 2208
rect 3450 2148 3454 2204
rect 3454 2148 3510 2204
rect 3510 2148 3514 2204
rect 3450 2144 3514 2148
rect 3530 2204 3594 2208
rect 3530 2148 3534 2204
rect 3534 2148 3590 2204
rect 3590 2148 3594 2204
rect 3530 2144 3594 2148
rect 3610 2204 3674 2208
rect 3610 2148 3614 2204
rect 3614 2148 3670 2204
rect 3670 2148 3674 2204
rect 3610 2144 3674 2148
rect 3690 2204 3754 2208
rect 3690 2148 3694 2204
rect 3694 2148 3750 2204
rect 3750 2148 3754 2204
rect 3690 2144 3754 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 13445 2204 13509 2208
rect 13445 2148 13449 2204
rect 13449 2148 13505 2204
rect 13505 2148 13509 2204
rect 13445 2144 13509 2148
rect 13525 2204 13589 2208
rect 13525 2148 13529 2204
rect 13529 2148 13585 2204
rect 13585 2148 13589 2204
rect 13525 2144 13589 2148
rect 13605 2204 13669 2208
rect 13605 2148 13609 2204
rect 13609 2148 13665 2204
rect 13665 2148 13669 2204
rect 13605 2144 13669 2148
rect 13685 2204 13749 2208
rect 13685 2148 13689 2204
rect 13689 2148 13745 2204
rect 13745 2148 13749 2204
rect 13685 2144 13749 2148
<< metal4 >>
rect 3442 17440 3763 17456
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3763 17440
rect 3442 16352 3763 17376
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3763 16352
rect 3442 15264 3763 16288
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3763 15264
rect 3442 14176 3763 15200
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3763 14176
rect 3442 13088 3763 14112
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3763 13088
rect 3442 12000 3763 13024
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3763 12000
rect 3442 10912 3763 11936
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3763 10912
rect 3442 9824 3763 10848
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3763 9824
rect 3442 8736 3763 9760
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3763 8736
rect 3442 7648 3763 8672
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3763 7648
rect 3442 6560 3763 7584
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3763 6560
rect 3442 5472 3763 6496
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3763 5472
rect 3442 4384 3763 5408
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3763 4384
rect 3442 3296 3763 4320
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3763 3296
rect 3442 2208 3763 3232
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3763 2208
rect 3442 2128 3763 2144
rect 5941 16896 6261 17456
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 15808 6261 16832
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 14720 6261 15744
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 13632 6261 14656
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 12544 6261 13568
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 11456 6261 12480
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 10368 6261 11392
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 9280 6261 10304
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 8192 6261 9216
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 7104 6261 8128
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 6016 6261 7040
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 4928 6261 5952
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 3840 6261 4864
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 2752 6261 3776
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2128 6261 2688
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10938 16896 11259 17456
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11259 16896
rect 10938 15808 11259 16832
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11259 15808
rect 10938 14720 11259 15744
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11259 14720
rect 10938 13632 11259 14656
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11259 13632
rect 10938 12544 11259 13568
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11259 12544
rect 10938 11456 11259 12480
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11259 11456
rect 10938 10368 11259 11392
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11259 10368
rect 10938 9280 11259 10304
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11259 9280
rect 10938 8192 11259 9216
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11259 8192
rect 10938 7104 11259 8128
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11259 7104
rect 10938 6016 11259 7040
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11259 6016
rect 10938 4928 11259 5952
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11259 4928
rect 10938 3840 11259 4864
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11259 3840
rect 10938 2752 11259 3776
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11259 2752
rect 10938 2128 11259 2688
rect 13437 17440 13757 17456
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 16352 13757 17376
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 15264 13757 16288
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 14176 13757 15200
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 13088 13757 14112
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 12000 13757 13024
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 10912 13757 11936
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 9824 13757 10848
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 8736 13757 9760
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 7648 13757 8672
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 6560 13757 7584
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 5472 13757 6496
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 4384 13757 5408
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 3296 13757 4320
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 13437 2208 13757 3232
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2128 13757 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output46
timestamp 1624635492
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2944 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform -1 0 3220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform -1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1624635492
transform -1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1840 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_26
timestamp 1624635492
transform 1 0 3496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform -1 0 3956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform -1 0 4232 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform -1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40
timestamp 1624635492
transform 1 0 4784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34
timestamp 1624635492
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform -1 0 4416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output48
timestamp 1624635492
transform -1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output47
timestamp 1624635492
transform -1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_36
timestamp 1624635492
transform 1 0 4416 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5520 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45
timestamp 1624635492
transform 1 0 5244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output50
timestamp 1624635492
transform -1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output49
timestamp 1624635492
transform -1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56
timestamp 1624635492
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output51
timestamp 1624635492
transform -1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output52
timestamp 1624635492
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform -1 0 7636 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform -1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1624635492
transform -1 0 8372 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform -1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1624635492
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1624635492
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1624635492
transform 1 0 9476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1624635492
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform -1 0 9844 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1624635492
transform 1 0 9752 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 10488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 10028 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform -1 0 10764 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1624635492
transform 1 0 10028 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_97
timestamp 1624635492
transform 1 0 10028 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_111
timestamp 1624635492
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105
timestamp 1624635492
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 11316 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 11316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1624635492
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1624635492
transform 1 0 10856 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_117
timestamp 1624635492
transform 1 0 11868 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 11868 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1624635492
transform 1 0 12144 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp 1624635492
transform 1 0 12604 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1624635492
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_130
timestamp 1624635492
transform 1 0 13064 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 13064 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 13064 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform -1 0 13340 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp 1624635492
transform 1 0 13616 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133
timestamp 1624635492
transform 1 0 13340 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1624635492
transform 1 0 13432 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_139
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1624635492
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1624635492
transform 1 0 13892 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_146
timestamp 1624635492
transform 1 0 14536 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1624635492
transform 1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 15180 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform 1 0 15364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1624635492
transform 1 0 15180 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1624635492
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1624635492
transform -1 0 15732 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1624635492
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1624635492
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1624635492
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1624635492
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1624635492
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1624635492
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1624635492
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1624635492
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1624635492
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1624635492
transform 1 0 15456 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1624635492
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1624635492
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1624635492
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1624635492
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1624635492
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1624635492
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1624635492
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1624635492
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1624635492
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1624635492
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_151
timestamp 1624635492
transform 1 0 14996 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1624635492
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1624635492
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1624635492
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1624635492
transform -1 0 9568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_92
timestamp 1624635492
transform 1 0 9568 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_104
timestamp 1624635492
transform 1 0 10672 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_116
timestamp 1624635492
transform 1 0 11776 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_128
timestamp 1624635492
transform 1 0 12880 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_140
timestamp 1624635492
transform 1 0 13984 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 16008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp 1624635492
transform 1 0 15456 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_7
timestamp 1624635492
transform 1 0 1748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1624635492
transform 1 0 2852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1624635492
transform 1 0 4784 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1624635492
transform 1 0 4416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_35
timestamp 1624635492
transform 1 0 4324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_39
timestamp 1624635492
transform 1 0 4692 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _02_
timestamp 1624635492
transform -1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _04_
timestamp 1624635492
transform -1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1624635492
transform 1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1624635492
transform 1 0 5152 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _41_
timestamp 1624635492
transform -1 0 5704 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp 1624635492
transform 1 0 5060 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_50
timestamp 1624635492
transform 1 0 5704 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _05_
timestamp 1624635492
transform -1 0 7268 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _06_
timestamp 1624635492
transform -1 0 7728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _07_
timestamp 1624635492
transform 1 0 7912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _08_
timestamp 1624635492
transform 1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1624635492
transform 1 0 8556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 1624635492
transform 1 0 6900 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_67
timestamp 1624635492
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_72
timestamp 1624635492
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1624635492
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _10_
timestamp 1624635492
transform -1 0 9384 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _11_
timestamp 1624635492
transform -1 0 9844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _12_
timestamp 1624635492
transform -1 0 10304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _13_
timestamp 1624635492
transform -1 0 10672 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1624635492
transform 1 0 8832 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1624635492
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp 1624635492
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_100
timestamp 1624635492
transform 1 0 10304 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_104
timestamp 1624635492
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _14_
timestamp 1624635492
transform -1 0 11132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _16_
timestamp 1624635492
transform -1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_
timestamp 1624635492
transform -1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _18_
timestamp 1624635492
transform -1 0 12880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1624635492
transform 1 0 11132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1624635492
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1624635492
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1624635492
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1624635492
transform 1 0 12880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1624635492
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_134
timestamp 1624635492
transform 1 0 13432 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_146
timestamp 1624635492
transform 1 0 14536 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1624635492
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1624635492
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624635492
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_33
timestamp 1624635492
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1624635492
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1624635492
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_45
timestamp 1624635492
transform 1 0 5244 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 1624635492
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_62
timestamp 1624635492
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1624635492
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1624635492
transform 1 0 6992 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1624635492
transform 1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1624635492
transform 1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1624635492
transform 1 0 7268 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1624635492
transform 1 0 7912 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1624635492
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1624635492
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1624635492
transform 1 0 9476 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1624635492
transform 1 0 9936 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_90
timestamp 1624635492
transform 1 0 9384 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_94
timestamp 1624635492
transform 1 0 9752 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_99
timestamp 1624635492
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1624635492
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1624635492
transform 1 0 10764 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1624635492
transform 1 0 11592 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_108
timestamp 1624635492
transform 1 0 11040 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1624635492
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1624635492
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1624635492
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1624635492
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1624635492
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1624635492
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp 1624635492
transform 1 0 15456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_151
timestamp 1624635492
transform 1 0 14996 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1624635492
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1624635492
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1624635492
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1624635492
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1624635492
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1624635492
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1624635492
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1624635492
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp 1624635492
transform 1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3312 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_23
timestamp 1624635492
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1624635492
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1624635492
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1624635492
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1624635492
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_106
timestamp 1624635492
transform 1 0 10856 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1624635492
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1624635492
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_151
timestamp 1624635492
transform 1 0 14996 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1624635492
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1624635492
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1624635492
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1624635492
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1624635492
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1624635492
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1624635492
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1624635492
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_156
timestamp 1624635492
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform -1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_7
timestamp 1624635492
transform 1 0 1748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_19
timestamp 1624635492
transform 1 0 2852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1624635492
transform 1 0 3956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1624635492
transform 1 0 5060 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1624635492
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1624635492
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1624635492
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1624635492
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1624635492
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1624635492
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1624635492
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_151
timestamp 1624635492
transform 1 0 14996 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1624635492
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6624 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1624635492
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_54
timestamp 1624635492
transform 1 0 6072 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_69
timestamp 1624635492
transform 1 0 7452 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_81
timestamp 1624635492
transform 1 0 8556 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1624635492
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1624635492
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_111
timestamp 1624635492
transform 1 0 11316 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_119
timestamp 1624635492
transform 1 0 12052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_136
timestamp 1624635492
transform 1 0 13616 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_142
timestamp 1624635492
transform 1 0 14168 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_156
timestamp 1624635492
transform 1 0 15456 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_12
timestamp 1624635492
transform 1 0 2208 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1624635492
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1624635492
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1624635492
transform 1 0 3312 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_28
timestamp 1624635492
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 7360 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1624635492
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1624635492
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1624635492
transform 1 0 6072 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1624635492
transform 1 0 6440 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8832 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7084 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 8280 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_64
timestamp 1624635492
transform 1 0 6992 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1624635492
transform 1 0 7912 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 9568 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_87
timestamp 1624635492
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1624635492
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1624635492
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1624635492
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_101
timestamp 1624635492
transform 1 0 10396 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_111
timestamp 1624635492
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_113
timestamp 1624635492
transform 1 0 11500 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_125
timestamp 1624635492
transform 1 0 12604 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1624635492
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1624635492
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_137
timestamp 1624635492
transform 1 0 13708 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_151
timestamp 1624635492
transform 1 0 14996 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_156
timestamp 1624635492
transform 1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1624635492
transform 1 0 2484 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1624635492
transform 1 0 3128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_26
timestamp 1624635492
transform 1 0 3496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_40
timestamp 1624635492
transform 1 0 4784 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform -1 0 7636 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1624635492
transform 1 0 5888 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1624635492
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9108 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9108 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9936 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_109
timestamp 1624635492
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1624635492
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1624635492
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1624635492
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_151
timestamp 1624635492
transform 1 0 14996 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1624635492
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 7360 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624635492
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1624635492
transform 1 0 6072 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1624635492
transform 1 0 6440 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _01_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 10120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1624635492
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1624635492
transform 1 0 9384 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_94
timestamp 1624635492
transform 1 0 9752 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_98
timestamp 1624635492
transform 1 0 10120 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_110
timestamp 1624635492
transform 1 0 11224 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_122
timestamp 1624635492
transform 1 0 12328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_134
timestamp 1624635492
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1624635492
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_156
timestamp 1624635492
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1624635492
transform -1 0 1656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 1840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_8
timestamp 1624635492
transform 1 0 1840 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_20
timestamp 1624635492
transform 1 0 2944 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1624635492
transform 1 0 4048 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8556 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1624635492
transform 1 0 5152 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_56
timestamp 1624635492
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8556 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_97
timestamp 1624635492
transform 1 0 10028 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_109
timestamp 1624635492
transform 1 0 11132 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1624635492
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1624635492
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1624635492
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_151
timestamp 1624635492
transform 1 0 14996 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624635492
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1624635492
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_54
timestamp 1624635492
transform 1 0 6072 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_62
timestamp 1624635492
transform 1 0 6808 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform -1 0 7728 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_72
timestamp 1624635492
transform 1 0 7728 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1624635492
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1624635492
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1624635492
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1624635492
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1624635492
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output45
timestamp 1624635492
transform 1 0 15364 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_152
timestamp 1624635492
transform 1 0 15088 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2760 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1624635492
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_15
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4416 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1624635492
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_39
timestamp 1624635492
transform 1 0 4692 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_25
timestamp 1624635492
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 5152 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_43
timestamp 1624635492
transform 1 0 5060 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1624635492
transform 1 0 5428 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_55
timestamp 1624635492
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_52
timestamp 1624635492
transform 1 0 5888 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1624635492
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1624635492
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_64
timestamp 1624635492
transform 1 0 6992 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp 1624635492
transform 1 0 8096 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1624635492
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1624635492
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1624635492
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1624635492
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1624635492
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1624635492
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1624635492
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1624635492
transform -1 0 15640 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 16008 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1624635492
transform 1 0 15180 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_151
timestamp 1624635492
transform 1 0 14996 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1624635492
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1624635492
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1624635492
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1624635492
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1624635492
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1624635492
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1624635492
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1624635492
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1624635492
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1624635492
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1624635492
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1624635492
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_151
timestamp 1624635492
transform 1 0 14996 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1624635492
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1624635492
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1624635492
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1624635492
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1624635492
transform 1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_87
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1624635492
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1624635492
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1624635492
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1624635492
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1624635492
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_156
timestamp 1624635492
transform 1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform -1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_7
timestamp 1624635492
transform 1 0 1748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_19
timestamp 1624635492
transform 1 0 2852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1624635492
transform 1 0 3864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1624635492
transform 1 0 4508 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_27
timestamp 1624635492
transform 1 0 3588 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_33
timestamp 1624635492
transform 1 0 4140 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_40
timestamp 1624635492
transform 1 0 4784 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1624635492
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_49
timestamp 1624635492
transform 1 0 5612 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1624635492
transform 1 0 7176 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1624635492
transform -1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_71
timestamp 1624635492
transform 1 0 7636 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_83
timestamp 1624635492
transform 1 0 8740 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_95
timestamp 1624635492
transform 1 0 9844 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_107
timestamp 1624635492
transform 1 0 10948 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1624635492
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1624635492
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1624635492
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_151
timestamp 1624635492
transform 1 0 14996 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1624635492
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1624635492
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1624635492
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1624635492
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1624635492
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1624635492
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1624635492
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1624635492
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1624635492
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1624635492
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 15640 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1624635492
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1624635492
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1624635492
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1624635492
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1624635492
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1624635492
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1624635492
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1624635492
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1624635492
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1624635492
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_139
timestamp 1624635492
transform 1 0 13892 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1624635492
transform -1 0 15732 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_147
timestamp 1624635492
transform 1 0 14628 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 2116 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform -1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1624635492
transform -1 0 1932 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform -1 0 1656 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 2300 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 3220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 2852 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 2484 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_13
timestamp 1624635492
transform 1 0 2300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1624635492
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_25
timestamp 1624635492
transform 1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 4232 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1624635492
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform -1 0 4600 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform -1 0 5152 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform -1 0 5520 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 5980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 6900 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1624635492
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1624635492
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_48
timestamp 1624635492
transform 1 0 5520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 7268 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 7636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 8096 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform -1 0 8464 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1624635492
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1624635492
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_71
timestamp 1624635492
transform 1 0 7636 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1624635492
transform 1 0 8464 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1624635492
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 9568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9108 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_96
timestamp 1624635492
transform 1 0 9936 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1624635492
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 9936 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 9936 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1624635492
transform -1 0 10212 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_102
timestamp 1624635492
transform 1 0 10488 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_99
timestamp 1624635492
transform 1 0 10212 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1624635492
transform -1 0 10764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1624635492
transform -1 0 10488 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 1624635492
transform 1 0 11316 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1624635492
transform 1 0 10764 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1624635492
transform -1 0 11592 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1624635492
transform -1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1624635492
transform -1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_120
timestamp 1624635492
transform 1 0 12144 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_117
timestamp 1624635492
transform 1 0 11868 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 12144 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1624635492
transform -1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1624635492
transform -1 0 12144 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 11776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform -1 0 12696 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_134
timestamp 1624635492
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_128
timestamp 1624635492
transform 1 0 12880 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 13156 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 13156 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1624635492
transform -1 0 12972 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1624635492
transform -1 0 13800 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1624635492
transform -1 0 13432 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 14536 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 13984 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1624635492
transform -1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_131
timestamp 1624635492
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 14904 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 14720 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1624635492
transform -1 0 15180 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1624635492
transform -1 0 15088 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1624635492
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform 1 0 15364 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1624635492
transform -1 0 15456 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1624635492
transform -1 0 15364 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1624635492
transform -1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 16400 12384 17200 12504 6 ccff_tail
port 2 nsew signal tristate
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_in[10]
port 4 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[11]
port 5 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_in[12]
port 6 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_in[13]
port 7 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_in[14]
port 8 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_in[15]
port 9 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_in[16]
port 10 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_in[17]
port 11 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_in[18]
port 12 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_in[19]
port 13 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[1]
port 14 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[2]
port 15 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[3]
port 16 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[4]
port 17 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[5]
port 18 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[6]
port 19 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[7]
port 20 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[8]
port 21 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_in[9]
port 22 nsew signal input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 23 nsew signal tristate
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_out[10]
port 24 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[11]
port 25 nsew signal tristate
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_out[12]
port 26 nsew signal tristate
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_out[13]
port 27 nsew signal tristate
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_out[14]
port 28 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_out[15]
port 29 nsew signal tristate
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_out[16]
port 30 nsew signal tristate
rlabel metal2 s 7470 0 7526 800 6 chany_bottom_out[17]
port 31 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 chany_bottom_out[18]
port 32 nsew signal tristate
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_out[19]
port 33 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 34 nsew signal tristate
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 35 nsew signal tristate
rlabel metal2 s 1490 0 1546 800 6 chany_bottom_out[3]
port 36 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 37 nsew signal tristate
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_out[5]
port 38 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[6]
port 39 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[7]
port 40 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_out[8]
port 41 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 chany_bottom_out[9]
port 42 nsew signal tristate
rlabel metal2 s 8942 19200 8998 20000 6 chany_top_in[0]
port 43 nsew signal input
rlabel metal2 s 13174 19200 13230 20000 6 chany_top_in[10]
port 44 nsew signal input
rlabel metal2 s 13542 19200 13598 20000 6 chany_top_in[11]
port 45 nsew signal input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[12]
port 46 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[13]
port 47 nsew signal input
rlabel metal2 s 14830 19200 14886 20000 6 chany_top_in[14]
port 48 nsew signal input
rlabel metal2 s 15290 19200 15346 20000 6 chany_top_in[15]
port 49 nsew signal input
rlabel metal2 s 15658 19200 15714 20000 6 chany_top_in[16]
port 50 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[17]
port 51 nsew signal input
rlabel metal2 s 16486 19200 16542 20000 6 chany_top_in[18]
port 52 nsew signal input
rlabel metal2 s 16946 19200 17002 20000 6 chany_top_in[19]
port 53 nsew signal input
rlabel metal2 s 9402 19200 9458 20000 6 chany_top_in[1]
port 54 nsew signal input
rlabel metal2 s 9770 19200 9826 20000 6 chany_top_in[2]
port 55 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[3]
port 56 nsew signal input
rlabel metal2 s 10690 19200 10746 20000 6 chany_top_in[4]
port 57 nsew signal input
rlabel metal2 s 11058 19200 11114 20000 6 chany_top_in[5]
port 58 nsew signal input
rlabel metal2 s 11518 19200 11574 20000 6 chany_top_in[6]
port 59 nsew signal input
rlabel metal2 s 11886 19200 11942 20000 6 chany_top_in[7]
port 60 nsew signal input
rlabel metal2 s 12346 19200 12402 20000 6 chany_top_in[8]
port 61 nsew signal input
rlabel metal2 s 12714 19200 12770 20000 6 chany_top_in[9]
port 62 nsew signal input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 63 nsew signal tristate
rlabel metal2 s 4802 19200 4858 20000 6 chany_top_out[10]
port 64 nsew signal tristate
rlabel metal2 s 5170 19200 5226 20000 6 chany_top_out[11]
port 65 nsew signal tristate
rlabel metal2 s 5630 19200 5686 20000 6 chany_top_out[12]
port 66 nsew signal tristate
rlabel metal2 s 5998 19200 6054 20000 6 chany_top_out[13]
port 67 nsew signal tristate
rlabel metal2 s 6458 19200 6514 20000 6 chany_top_out[14]
port 68 nsew signal tristate
rlabel metal2 s 6826 19200 6882 20000 6 chany_top_out[15]
port 69 nsew signal tristate
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[16]
port 70 nsew signal tristate
rlabel metal2 s 7746 19200 7802 20000 6 chany_top_out[17]
port 71 nsew signal tristate
rlabel metal2 s 8114 19200 8170 20000 6 chany_top_out[18]
port 72 nsew signal tristate
rlabel metal2 s 8574 19200 8630 20000 6 chany_top_out[19]
port 73 nsew signal tristate
rlabel metal2 s 1030 19200 1086 20000 6 chany_top_out[1]
port 74 nsew signal tristate
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 75 nsew signal tristate
rlabel metal2 s 1858 19200 1914 20000 6 chany_top_out[3]
port 76 nsew signal tristate
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 77 nsew signal tristate
rlabel metal2 s 2686 19200 2742 20000 6 chany_top_out[5]
port 78 nsew signal tristate
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 79 nsew signal tristate
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[7]
port 80 nsew signal tristate
rlabel metal2 s 3974 19200 4030 20000 6 chany_top_out[8]
port 81 nsew signal tristate
rlabel metal2 s 4342 19200 4398 20000 6 chany_top_out[9]
port 82 nsew signal tristate
rlabel metal3 s 0 8304 800 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew signal tristate
rlabel metal3 s 0 4904 800 5024 6 left_grid_pin_0_
port 86 nsew signal tristate
rlabel metal3 s 16400 7352 17200 7472 6 prog_clk_0_E_in
port 87 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 right_width_0_height_0__pin_0_
port 88 nsew signal input
rlabel metal3 s 16400 2456 17200 2576 6 right_width_0_height_0__pin_1_lower
port 89 nsew signal tristate
rlabel metal3 s 16400 17416 17200 17536 6 right_width_0_height_0__pin_1_upper
port 90 nsew signal tristate
rlabel metal4 s 13437 2128 13757 17456 6 VPWR
port 91 nsew power bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VPWR
port 92 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 17456 6 VPWR
port 93 nsew power bidirectional
rlabel metal4 s 10939 2128 11259 17456 6 VGND
port 94 nsew ground bidirectional
rlabel metal4 s 5941 2128 6261 17456 6 VGND
port 95 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
