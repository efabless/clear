* NGSPICE file created from sb_0__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt sb_0__1_ bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk_0_E_in right_bottom_grid_pin_34_ right_bottom_grid_pin_35_
+ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_
+ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ top_left_grid_pin_1_ VPWR VGND
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_20.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l1_in_1_ input5/X input17/X mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__124__A _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_1
X_062_ VGND VGND VPWR VPWR _062_/HI _062_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input55_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__119__A _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_2__A1 input68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_114_ _114_/A VGND VGND VPWR VPWR _114_/X sky130_fd_sc_hd__clkbuf_1
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l1_in_0_ _104_/A _095_/A mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input18_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput75 _077_/X VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__clkbuf_2
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_1
Xoutput97 _099_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput86 _069_/X VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_0_ _100_/A _091_/A mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_10.mux_l2_in_0__A0 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_26.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ VGND VGND VPWR VPWR _061_/HI _061_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input48_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_113_ _113_/A VGND VGND VPWR VPWR _113_/X sky130_fd_sc_hd__clkbuf_1
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput76 _078_/X VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput98 _100_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput87 _070_/X VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input30_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_1__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_mem_bottom_track_1.prog_clk clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_10.mux_l3_in_0_ mux_right_track_10.mux_l2_in_1_/X mux_right_track_10.mux_l2_in_0_/X
+ mux_right_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_060_ VGND VGND VPWR VPWR _060_/HI _060_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
X_112_ _112_/A VGND VGND VPWR VPWR _112_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input60_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.mux_l2_in_1_ _062_/HI _116_/A mux_right_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput77 _079_/X VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput99 _101_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput88 _071_/X VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input23_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_6.mux_l1_in_1__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_0_FTB00 prog_clk_0_E_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_111_ _111_/A VGND VGND VPWR VPWR _111_/X sky130_fd_sc_hd__clkbuf_1
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input53_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.mux_l2_in_0_ input64/X mux_right_track_10.mux_l1_in_0_/X mux_right_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput78 _080_/X VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput89 _072_/X VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input16_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_1_ _046_/HI _115_/A mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ _047_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input8_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l1_in_0__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_2_ _119_/A _109_/A mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _114_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_110_ _110_/A VGND VGND VPWR VPWR _110_/X sky130_fd_sc_hd__clkbuf_1
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input46_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__buf_1
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_12.mux_l2_in_1__A1 _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput79 _081_/X VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__clkbuf_2
Xmux_right_track_10.mux_l1_in_0_ input45/X _096_/A mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ input63/X mux_right_track_8.mux_l1_in_0_/X mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_22.mux_l2_in_0_ mux_right_track_22.mux_l1_in_1_/X mux_right_track_22.mux_l1_in_0_/X
+ mux_right_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_22.mux_l1_in_0__A1 _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_1_ input9/X input21/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_22.mux_l1_in_1_ _036_/HI _124_/A mux_right_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input39_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _071_/A sky130_fd_sc_hd__buf_1
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_30.mux_l1_in_0__A1 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input21_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l1_in_0_ _095_/A input60/X mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__089__A _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_0_ input14/X input71/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input69_A right_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_22.mux_l1_in_0_ _085_/A _104_/A mux_right_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_18.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_34.mux_l2_in_0_ _042_/HI mux_right_track_34.mux_l1_in_0_/X mux_right_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _070_/A sky130_fd_sc_hd__buf_1
Xmux_bottom_track_25.mux_l2_in_1_ _056_/HI input8/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input51_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_1_ _060_/HI mux_bottom_track_9.mux_l1_in_2_/X mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l1_in_2_ input1/X input10/X mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input14_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__buf_1
XANTENNA_input6_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_30.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_34.mux_l1_in_0_ input34/X input68/X mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_1_ input20/X input3/X mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input44_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l1_in_1_ input22/X input15/X mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_28.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l2_in_1_ _048_/HI _124_/A mux_top_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_0_ _105_/A _096_/A mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input37_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_36.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l1_in_0_ _103_/A _093_/A mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input67_A right_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__100__A _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_3_ _044_/HI _112_/A mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_34.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l1_in_1_ _115_/A input13/X mux_top_track_16.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_36.mux_l1_in_0__A0 input23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input12_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_28.mux_l1_in_0__A1 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input4_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l1_in_2_ input69/X input67/X mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ input6/X input18/X mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l1_in_1_ _065_/HI _120_/A mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_1_ input65/X input63/X mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_22.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__125__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input65_A right_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 bottom_left_grid_pin_1_ VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_1
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_16.mux_l1_in_0_ input67/X _100_/A mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_0_ _092_/A input54/X mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_28.mux_l2_in_0_ _039_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _068_/A sky130_fd_sc_hd__clkbuf_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input28_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_30.mux_l2_in_0_ _040_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_2
X_059_ VGND VGND VPWR VPWR _059_/HI _059_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 right_bottom_grid_pin_41_ VGND VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_1_ _059_/HI mux_bottom_track_5.mux_l1_in_2_/X mux_bottom_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input10_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input2_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input58_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 ccff_head VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_5.mux_l1_in_2_ input1/X input11/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_28.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ VGND VGND VPWR VPWR _058_/HI _058_/LO sky130_fd_sc_hd__conb_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput60 chany_top_in[7] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
Xinput71 top_left_grid_pin_1_ VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input40_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l1_in_0_ input25/X input65/X mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_30.mux_l1_in_0_ input40/X input66/X mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 chanx_right_in[0] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_1
Xmux_bottom_track_5.mux_l1_in_1_ input4/X input16/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input70_A right_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_26.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_12.mux_l2_in_0__A0 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_057_ VGND VGND VPWR VPWR _057_/HI _057_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput50 chany_top_in[16] VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_2
Xinput61 chany_top_in[8] VGND VGND VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_E_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input33_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ _109_/A VGND VGND VPWR VPWR _109_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ output72/A VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_1
Xinput4 chanx_right_in[10] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
Xmux_bottom_track_5.mux_l1_in_0_ _101_/A _092_/A mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_1_ _058_/HI input7/X mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input63_A right_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_125_ _125_/A VGND VGND VPWR VPWR _125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_056_ VGND VGND VPWR VPWR _056_/HI _056_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput51 chany_top_in[17] VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__clkbuf_2
Xinput62 chany_top_in[9] VGND VGND VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_2
Xinput40 chany_bottom_in[7] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_1_0_mem_bottom_track_1.prog_clk clkbuf_3_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input26_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A VGND VGND VPWR VPWR _108_/X sky130_fd_sc_hd__clkbuf_1
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_20.mux_l1_in_1__A1 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 chanx_right_in[11] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_1
Xmux_top_track_24.mux_l2_in_1_ _050_/HI _125_/A mux_top_track_24.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_33.mux_l1_in_0_ input19/X _097_/A mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input56_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_6.mux_l1_in_3__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_124_ _124_/A VGND VGND VPWR VPWR _124_/X sky130_fd_sc_hd__clkbuf_1
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.mux_l3_in_0_ mux_right_track_12.mux_l2_in_1_/X mux_right_track_12.mux_l2_in_0_/X
+ mux_right_track_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput52 chany_top_in[18] VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__clkbuf_2
Xinput63 right_bottom_grid_pin_34_ VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_2
Xinput41 chany_bottom_in[8] VGND VGND VPWR VPWR _115_/A sky130_fd_sc_hd__clkbuf_2
Xinput30 chany_bottom_in[16] VGND VGND VPWR VPWR _123_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input19_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.mux_l2_in_1_ _063_/HI _117_/A mux_right_track_12.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_1_ _061_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_2_ _109_/A input69/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__092__A _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput6 chanx_right_in[12] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l2_in_0_ _116_/A mux_top_track_24.mux_l1_in_0_/X mux_top_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input49_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_123_ _123_/A VGND VGND VPWR VPWR _123_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
Xinput31 chany_bottom_in[17] VGND VGND VPWR VPWR _124_/A sky130_fd_sc_hd__clkbuf_2
Xinput20 chanx_right_in[7] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
Xinput53 chany_top_in[19] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 right_bottom_grid_pin_35_ VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
Xinput42 chany_bottom_in[9] VGND VGND VPWR VPWR _116_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_12.mux_l2_in_0_ input65/X mux_right_track_12.mux_l1_in_0_/X mux_right_track_12.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input31_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_14.mux_l2_in_1__A1 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ input67/X input65/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l2_in_1_ _049_/HI _120_/A mux_top_track_2.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l2_in_1_ _037_/HI input33/X mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 chanx_right_in[13] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _118_/A sky130_fd_sc_hd__clkbuf_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput130 _113_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__clkbuf_2
X_122_ _122_/A VGND VGND VPWR VPWR _122_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input61_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_0_ input7/X input19/X mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput43 chany_top_in[0] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__buf_1
Xinput54 chany_top_in[1] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_1
Xinput32 chany_bottom_in[18] VGND VGND VPWR VPWR _125_/A sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_right_in[8] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_1
Xinput10 chanx_right_in[16] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__buf_1
Xinput65 right_bottom_grid_pin_36_ VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input24_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _066_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_12.mux_l1_in_0_ input49/X _097_/A mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_0_ input63/X _089_/A mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_24.mux_l2_in_0_ _125_/A mux_right_track_24.mux_l1_in_0_/X mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput8 chanx_right_in[14] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_2.mux_l1_in_1_ _111_/A input10/X mux_top_track_2.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput131 _114_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__clkbuf_2
Xoutput120 _122_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__clkbuf_2
X_121_ _121_/A VGND VGND VPWR VPWR _121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input54_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xinput44 chany_top_in[10] VGND VGND VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_2
Xinput55 chany_top_in[2] VGND VGND VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_2
Xinput33 chany_bottom_in[19] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput66 right_bottom_grid_pin_37_ VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__clkbuf_2
Xinput22 chanx_right_in[9] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_1
Xinput11 chanx_right_in[17] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_1
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_1_ _054_/HI mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l1_in_2_ input1/X input13/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input9_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 chanx_right_in[15] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_1
Xclkbuf_3_0_0_mem_bottom_track_1.prog_clk clkbuf_3_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_18.mux_l1_in_1__A1 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_0_ input22/X input15/X mux_top_track_2.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_24.mux_l1_in_0_ input63/X _105_/A mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput121 _123_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__clkbuf_2
Xoutput132 _115_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__clkbuf_2
Xoutput110 _093_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A mux_right_track_34.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_120_ _120_/A VGND VGND VPWR VPWR _120_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_36.mux_l2_in_0_ _043_/HI mux_right_track_36.mux_l1_in_0_/X mux_right_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input47_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_30.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput45 chany_top_in[11] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_1
Xinput56 chany_top_in[3] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_1
Xinput67 right_bottom_grid_pin_38_ VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__clkbuf_2
Xinput23 chany_bottom_in[0] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__buf_1
Xinput34 chany_bottom_in[1] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__buf_1
Xinput12 chanx_right_in[18] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_1
XFILLER_20_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_1_ input6/X input18/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__101__A _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ input2/X VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput122 _124_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__clkbuf_2
Xoutput111 _094_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__clkbuf_2
Xoutput100 _102_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__clkbuf_2
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 chanx_right_in[19] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_1
Xinput46 chany_top_in[12] VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_2
Xinput57 chany_top_in[4] VGND VGND VPWR VPWR _091_/A sky130_fd_sc_hd__clkbuf_2
Xinput68 right_bottom_grid_pin_39_ VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_2
Xinput35 chany_bottom_in[2] VGND VGND VPWR VPWR _109_/A sky130_fd_sc_hd__clkbuf_2
Xinput24 chany_bottom_in[10] VGND VGND VPWR VPWR _117_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_1
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_36.mux_l1_in_0_ input23/X input69/X mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__104__A _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l1_in_0_ _099_/A _089_/A mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__112__A _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput123 _125_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput101 _103_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__clkbuf_2
Xoutput112 _095_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xinput14 chanx_right_in[1] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__buf_1
Xinput36 chany_bottom_in[3] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__buf_1
Xinput25 chany_bottom_in[11] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xinput47 chany_top_in[13] VGND VGND VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_2
Xinput58 chany_top_in[5] VGND VGND VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_2
Xinput69 right_bottom_grid_pin_40_ VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input52_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__120__A _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input15_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input7_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput124 _107_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput113 _106_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput102 _104_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_6.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput48 chany_top_in[14] VGND VGND VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_2
Xinput59 chany_top_in[6] VGND VGND VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_right_in[2] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_1
Xinput37 chany_bottom_in[4] VGND VGND VPWR VPWR _111_/A sky130_fd_sc_hd__clkbuf_2
Xinput26 chany_bottom_in[12] VGND VGND VPWR VPWR _119_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__123__A _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input45_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l1_in_3_ _045_/HI _113_/A mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l2_in_1_ _051_/HI _117_/A mux_top_track_32.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput114 _116_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput125 _108_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput103 _105_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput49 chany_top_in[15] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
Xinput16 chanx_right_in[3] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_1
Xinput38 chany_bottom_in[5] VGND VGND VPWR VPWR _112_/A sky130_fd_sc_hd__clkbuf_2
Xinput27 chany_bottom_in[13] VGND VGND VPWR VPWR _120_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input38_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l2_in_1_ mux_right_track_6.mux_l1_in_3_/X mux_right_track_6.mux_l1_in_2_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l1_in_3__A1 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l1_in_2_ _085_/A input68/X mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input20_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_32.mux_l2_in_0_ input8/X mux_top_track_32.mux_l1_in_0_/X mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input68_A right_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput115 _117_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput126 _109_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput104 _087_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 chany_bottom_in[6] VGND VGND VPWR VPWR _113_/A sky130_fd_sc_hd__clkbuf_2
Xinput28 chany_bottom_in[14] VGND VGND VPWR VPWR _121_/A sky130_fd_sc_hd__clkbuf_2
Xinput17 chanx_right_in[4] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_1
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_18.mux_l2_in_0_ mux_right_track_18.mux_l1_in_1_/X mux_right_track_18.mux_l1_in_0_/X
+ mux_right_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_20.mux_l2_in_0_ mux_right_track_20.mux_l1_in_1_/X mux_right_track_20.mux_l1_in_0_/X
+ mux_right_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input50_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.mux_l1_in_1_ _033_/HI _121_/A mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l1_in_1_ input66/X input64/X mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l2_in_1_ _053_/HI mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l1_in_1_ _035_/HI _123_/A mux_right_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input13_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input5_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_2_ _123_/A _113_/A mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput116 _118_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput127 _110_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput105 _088_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_right_track_6.mux_l1_in_2__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_right_in[5] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
Xinput29 chany_bottom_in[15] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_32.mux_l1_in_0_ input20/X input3/X mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_10.mux_l2_in_1__A1 _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input43_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_20.mux_l1_in_0__A1 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.mux_l1_in_0_ input68/X _101_/A mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_36.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l1_in_0_ _093_/A input56/X mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l1_in_0_ input69/X _103_/A mux_right_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_32.mux_l2_in_0_ _041_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_1_ input12/X input5/X mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _110_/A sky130_fd_sc_hd__clkbuf_1
Xoutput117 _119_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput128 _111_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput106 _089_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_2__A1 input68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 chanx_right_in[6] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input36_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l1_in_0_ input17/X input71/X mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput107 _090_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput118 _120_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput129 _112_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_0_ input36/X input67/X mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input66_A right_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__093__A _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input11_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput119 _121_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput108 _091_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput90 _073_/X VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input3_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input59_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l1_in_1__A1 _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_18.mux_l1_in_0__A0 input68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput109 _092_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput80 _082_/X VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__clkbuf_2
XANTENNA_output72_A output72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput91 _074_/X VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A0 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input71_A top_left_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_3_ _034_/HI _111_/A mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ _067_/A VGND VGND VPWR VPWR _067_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input34_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_119_ _119_/A VGND VGND VPWR VPWR _119_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_14.mux_l3_in_0_ mux_right_track_14.mux_l2_in_1_/X mux_right_track_14.mux_l2_in_0_/X
+ mux_right_track_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput81 _083_/X VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__clkbuf_2
Xmux_right_track_14.mux_l2_in_1_ _064_/HI _119_/A mux_right_track_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xoutput92 _075_/X VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A mux_right_track_30.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input64_A right_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_2_ _085_/A input68/X mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_066_ _066_/A VGND VGND VPWR VPWR _066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_34.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input27_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_118_ _118_/A VGND VGND VPWR VPWR _118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l1_in_1_/S VGND VGND VPWR VPWR output72/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput82 _084_/X VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__clkbuf_2
Xoutput93 _086_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__clkbuf_2
Xmux_right_track_14.mux_l2_in_0_ input66/X mux_right_track_14.mux_l1_in_0_/X mux_right_track_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2__A0 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input1_A bottom_left_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A1 _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input57_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_1_ input66/X input64/X mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ _052_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _122_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A mux_right_track_36.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_34.mux_l1_in_0__A1 input68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ VGND VGND VPWR VPWR _065_/HI _065_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_mem_bottom_track_1.prog_clk clkbuf_3_5_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l1_in_2_ _121_/A _112_/A mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_117_ _117_/A VGND VGND VPWR VPWR _117_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput83 _085_/X VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput94 _096_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput72 output72/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__clkbuf_2
XFILLER_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l2_in_1__A1 _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_8.mux_l1_in_2__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _067_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_14.mux_l1_in_0_ input53/X _099_/A mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_2.mux_l1_in_0_ _091_/A input43/X mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_26.mux_l2_in_0_ _038_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_064_ VGND VGND VPWR VPWR _064_/HI _064_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_1_ _055_/HI input9/X mux_bottom_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_1_ input11/X input4/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ _116_/A VGND VGND VPWR VPWR _116_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input32_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_32.mux_l2_in_1__A1 _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ _057_/HI input12/X mux_bottom_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput95 _097_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput73 _066_/X VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput84 _067_/X VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ VGND VGND VPWR VPWR _063_/HI _063_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input62_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.mux_l1_in_0_ input16/X input71/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l1_in_2__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_26.mux_l1_in_0_ input29/X input64/X mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
X_115_ _115_/A VGND VGND VPWR VPWR _115_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__121__A _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ input21/X input14/X mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__116__A _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S output72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput74 _076_/X VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput96 _098_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput85 _068_/X VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

