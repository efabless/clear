magic
tech sky130A
magscale 1 2
timestamp 1682557368
<< viali >>
rect 14565 54281 14599 54315
rect 16405 54281 16439 54315
rect 24501 54281 24535 54315
rect 24685 54281 24719 54315
rect 10977 54213 11011 54247
rect 14105 54213 14139 54247
rect 18889 54213 18923 54247
rect 21465 54213 21499 54247
rect 23305 54213 23339 54247
rect 3433 54145 3467 54179
rect 6009 54145 6043 54179
rect 8585 54145 8619 54179
rect 9965 54145 9999 54179
rect 11713 54145 11747 54179
rect 12541 54145 12575 54179
rect 14841 54145 14875 54179
rect 15853 54145 15887 54179
rect 16129 54145 16163 54179
rect 16865 54145 16899 54179
rect 17877 54145 17911 54179
rect 18521 54145 18555 54179
rect 19717 54145 19751 54179
rect 20453 54145 20487 54179
rect 21189 54145 21223 54179
rect 22293 54145 22327 54179
rect 22753 54145 22787 54179
rect 24041 54145 24075 54179
rect 25329 54145 25363 54179
rect 2973 54077 3007 54111
rect 5549 54077 5583 54111
rect 8125 54077 8159 54111
rect 12817 54077 12851 54111
rect 17693 54009 17727 54043
rect 11897 53941 11931 53975
rect 15025 53941 15059 53975
rect 15669 53941 15703 53975
rect 17049 53941 17083 53975
rect 18429 53941 18463 53975
rect 19533 53941 19567 53975
rect 20269 53941 20303 53975
rect 21005 53941 21039 53975
rect 22109 53941 22143 53975
rect 22937 53941 22971 53975
rect 23857 53941 23891 53975
rect 25145 53941 25179 53975
rect 16405 53737 16439 53771
rect 18889 53737 18923 53771
rect 9781 53669 9815 53703
rect 21833 53669 21867 53703
rect 23121 53669 23155 53703
rect 2973 53601 3007 53635
rect 6285 53601 6319 53635
rect 8125 53601 8159 53635
rect 11069 53601 11103 53635
rect 12725 53601 12759 53635
rect 24409 53601 24443 53635
rect 3433 53533 3467 53567
rect 4629 53533 4663 53567
rect 6745 53533 6779 53567
rect 8585 53533 8619 53567
rect 9137 53533 9171 53567
rect 11805 53533 11839 53567
rect 12449 53533 12483 53567
rect 14565 53533 14599 53567
rect 14841 53533 14875 53567
rect 15761 53533 15795 53567
rect 16129 53533 16163 53567
rect 16681 53533 16715 53567
rect 17417 53533 17451 53567
rect 18337 53533 18371 53567
rect 18705 53533 18739 53567
rect 19441 53533 19475 53567
rect 20361 53533 20395 53567
rect 20729 53533 20763 53567
rect 21097 53533 21131 53567
rect 22017 53533 22051 53567
rect 22661 53533 22695 53567
rect 23305 53533 23339 53567
rect 23949 53533 23983 53567
rect 25237 53533 25271 53567
rect 3985 53397 4019 53431
rect 14381 53397 14415 53431
rect 15669 53397 15703 53431
rect 16865 53397 16899 53431
rect 17601 53397 17635 53431
rect 18245 53397 18279 53431
rect 19625 53397 19659 53431
rect 20269 53397 20303 53431
rect 21281 53397 21315 53431
rect 22477 53397 22511 53431
rect 23857 53397 23891 53431
rect 25145 53397 25179 53431
rect 17325 53193 17359 53227
rect 19533 53193 19567 53227
rect 19717 53193 19751 53227
rect 21005 53193 21039 53227
rect 21189 53193 21223 53227
rect 21833 53193 21867 53227
rect 22293 53193 22327 53227
rect 22569 53193 22603 53227
rect 23029 53193 23063 53227
rect 13829 53125 13863 53159
rect 2329 53057 2363 53091
rect 4077 53057 4111 53091
rect 6009 53057 6043 53091
rect 7205 53057 7239 53091
rect 9137 53057 9171 53091
rect 9781 53057 9815 53091
rect 11897 53057 11931 53091
rect 14473 53057 14507 53091
rect 14933 53057 14967 53091
rect 15945 53057 15979 53091
rect 16405 53057 16439 53091
rect 19073 53057 19107 53091
rect 19349 53057 19383 53091
rect 20545 53057 20579 53091
rect 20821 53057 20855 53091
rect 23489 53057 23523 53091
rect 24133 53057 24167 53091
rect 24409 53057 24443 53091
rect 24777 53057 24811 53091
rect 25329 53057 25363 53091
rect 3709 52989 3743 53023
rect 5549 52989 5583 53023
rect 8861 52989 8895 53023
rect 10333 52989 10367 53023
rect 12357 52989 12391 53023
rect 14013 52921 14047 52955
rect 14657 52921 14691 52955
rect 1685 52853 1719 52887
rect 6561 52853 6595 52887
rect 16129 52853 16163 52887
rect 18889 52853 18923 52887
rect 20361 52853 20395 52887
rect 23305 52853 23339 52887
rect 23949 52853 23983 52887
rect 25145 52853 25179 52887
rect 9229 52649 9263 52683
rect 12633 52649 12667 52683
rect 14105 52649 14139 52683
rect 24593 52649 24627 52683
rect 25145 52581 25179 52615
rect 2973 52513 3007 52547
rect 6285 52513 6319 52547
rect 7757 52513 7791 52547
rect 11253 52513 11287 52547
rect 3341 52445 3375 52479
rect 3985 52445 4019 52479
rect 6745 52445 6779 52479
rect 8585 52445 8619 52479
rect 10793 52445 10827 52479
rect 12817 52445 12851 52479
rect 13645 52445 13679 52479
rect 24777 52445 24811 52479
rect 25329 52445 25363 52479
rect 9321 52377 9355 52411
rect 13461 52377 13495 52411
rect 4629 52309 4663 52343
rect 7205 52105 7239 52139
rect 11897 52105 11931 52139
rect 12541 52105 12575 52139
rect 13277 52105 13311 52139
rect 25237 52105 25271 52139
rect 3249 52037 3283 52071
rect 4813 52037 4847 52071
rect 7481 52037 7515 52071
rect 9873 52037 9907 52071
rect 1593 51969 1627 52003
rect 4077 51969 4111 52003
rect 6009 51969 6043 52003
rect 6561 51969 6595 52003
rect 9045 51969 9079 52003
rect 10885 51969 10919 52003
rect 11713 51969 11747 52003
rect 12357 51969 12391 52003
rect 8493 51901 8527 51935
rect 2237 51833 2271 51867
rect 25421 51765 25455 51799
rect 10241 51561 10275 51595
rect 2881 51425 2915 51459
rect 5549 51425 5583 51459
rect 7297 51425 7331 51459
rect 3433 51357 3467 51391
rect 4629 51357 4663 51391
rect 6653 51357 6687 51391
rect 8493 51357 8527 51391
rect 10425 51357 10459 51391
rect 25329 51357 25363 51391
rect 3985 51221 4019 51255
rect 25145 51221 25179 51255
rect 1777 51017 1811 51051
rect 7665 51017 7699 51051
rect 2789 50949 2823 50983
rect 4353 50949 4387 50983
rect 6837 50949 6871 50983
rect 9413 50949 9447 50983
rect 9597 50949 9631 50983
rect 1593 50881 1627 50915
rect 3709 50881 3743 50915
rect 5457 50881 5491 50915
rect 7021 50881 7055 50915
rect 7757 50881 7791 50915
rect 24777 50881 24811 50915
rect 25329 50881 25363 50915
rect 25145 50677 25179 50711
rect 9229 50473 9263 50507
rect 2237 50337 2271 50371
rect 7205 50337 7239 50371
rect 24869 50337 24903 50371
rect 3433 50269 3467 50303
rect 3985 50269 4019 50303
rect 7481 50269 7515 50303
rect 9413 50269 9447 50303
rect 24685 50269 24719 50303
rect 25329 50269 25363 50303
rect 4629 50133 4663 50167
rect 25145 50133 25179 50167
rect 11897 49929 11931 49963
rect 2145 49861 2179 49895
rect 4261 49861 4295 49895
rect 6377 49861 6411 49895
rect 9505 49861 9539 49895
rect 3341 49793 3375 49827
rect 3985 49793 4019 49827
rect 9321 49793 9355 49827
rect 11713 49793 11747 49827
rect 6009 49725 6043 49759
rect 25053 49725 25087 49759
rect 25329 49725 25363 49759
rect 12817 49385 12851 49419
rect 1777 49249 1811 49283
rect 2973 49181 3007 49215
rect 13001 49181 13035 49215
rect 24869 49181 24903 49215
rect 25329 49181 25363 49215
rect 3341 49045 3375 49079
rect 25145 49045 25179 49079
rect 25053 48705 25087 48739
rect 25329 48637 25363 48671
rect 18337 48229 18371 48263
rect 17325 48161 17359 48195
rect 17509 48161 17543 48195
rect 17601 48093 17635 48127
rect 19441 48093 19475 48127
rect 17969 47957 18003 47991
rect 20085 47957 20119 47991
rect 25237 47957 25271 47991
rect 25421 47957 25455 47991
rect 9229 47753 9263 47787
rect 11897 47753 11931 47787
rect 17233 47753 17267 47787
rect 17325 47753 17359 47787
rect 19533 47685 19567 47719
rect 9413 47617 9447 47651
rect 11713 47617 11747 47651
rect 20269 47617 20303 47651
rect 17417 47549 17451 47583
rect 19809 47549 19843 47583
rect 25053 47549 25087 47583
rect 25329 47549 25363 47583
rect 16865 47413 16899 47447
rect 18061 47413 18095 47447
rect 20913 47413 20947 47447
rect 7389 47209 7423 47243
rect 17785 47209 17819 47243
rect 19349 47209 19383 47243
rect 20913 47209 20947 47243
rect 18153 47141 18187 47175
rect 19625 47141 19659 47175
rect 22017 47141 22051 47175
rect 10057 47073 10091 47107
rect 15669 47073 15703 47107
rect 18797 47073 18831 47107
rect 20085 47073 20119 47107
rect 20177 47073 20211 47107
rect 21465 47073 21499 47107
rect 23765 47073 23799 47107
rect 7573 47005 7607 47039
rect 12265 47005 12299 47039
rect 17417 47005 17451 47039
rect 19993 47005 20027 47039
rect 20637 47005 20671 47039
rect 21649 47005 21683 47039
rect 24041 47005 24075 47039
rect 10333 46937 10367 46971
rect 17141 46937 17175 46971
rect 18521 46937 18555 46971
rect 21557 46937 21591 46971
rect 24501 46937 24535 46971
rect 11805 46869 11839 46903
rect 12909 46869 12943 46903
rect 14197 46869 14231 46903
rect 18613 46869 18647 46903
rect 25421 46869 25455 46903
rect 9045 46665 9079 46699
rect 10609 46665 10643 46699
rect 11897 46665 11931 46699
rect 16313 46665 16347 46699
rect 19073 46665 19107 46699
rect 22661 46665 22695 46699
rect 8033 46597 8067 46631
rect 22109 46597 22143 46631
rect 8217 46529 8251 46563
rect 8861 46529 8895 46563
rect 10793 46529 10827 46563
rect 18613 46529 18647 46563
rect 22753 46529 22787 46563
rect 25053 46529 25087 46563
rect 13829 46461 13863 46495
rect 14105 46461 14139 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 18337 46461 18371 46495
rect 20545 46461 20579 46495
rect 20821 46461 20855 46495
rect 22569 46461 22603 46495
rect 25329 46461 25363 46495
rect 7665 46325 7699 46359
rect 12357 46325 12391 46359
rect 16865 46325 16899 46359
rect 23121 46325 23155 46359
rect 11437 46121 11471 46155
rect 14197 46121 14231 46155
rect 16681 46121 16715 46155
rect 17785 46121 17819 46155
rect 7757 46053 7791 46087
rect 9137 46053 9171 46087
rect 10885 45985 10919 46019
rect 11897 45985 11931 46019
rect 16221 45985 16255 46019
rect 20729 45985 20763 46019
rect 20913 45985 20947 46019
rect 17325 45917 17359 45951
rect 18429 45917 18463 45951
rect 24041 45917 24075 45951
rect 24593 45917 24627 45951
rect 7941 45849 7975 45883
rect 9321 45849 9355 45883
rect 10977 45849 11011 45883
rect 12173 45849 12207 45883
rect 15945 45849 15979 45883
rect 20637 45849 20671 45883
rect 21281 45849 21315 45883
rect 23765 45849 23799 45883
rect 8401 45781 8435 45815
rect 9689 45781 9723 45815
rect 11069 45781 11103 45815
rect 13645 45781 13679 45815
rect 14473 45781 14507 45815
rect 20269 45781 20303 45815
rect 22293 45781 22327 45815
rect 25237 45781 25271 45815
rect 11253 45577 11287 45611
rect 14565 45577 14599 45611
rect 18153 45577 18187 45611
rect 8677 45509 8711 45543
rect 9321 45509 9355 45543
rect 11713 45509 11747 45543
rect 16865 45509 16899 45543
rect 20729 45509 20763 45543
rect 23489 45509 23523 45543
rect 11897 45441 11931 45475
rect 13737 45441 13771 45475
rect 15209 45441 15243 45475
rect 17509 45441 17543 45475
rect 18797 45441 18831 45475
rect 23765 45441 23799 45475
rect 9045 45373 9079 45407
rect 11161 45373 11195 45407
rect 13829 45373 13863 45407
rect 13921 45373 13955 45407
rect 21005 45373 21039 45407
rect 24225 45373 24259 45407
rect 24501 45373 24535 45407
rect 24777 45373 24811 45407
rect 10793 45305 10827 45339
rect 13369 45305 13403 45339
rect 6469 45237 6503 45271
rect 12265 45237 12299 45271
rect 19257 45237 19291 45271
rect 22017 45237 22051 45271
rect 6101 45033 6135 45067
rect 6653 45033 6687 45067
rect 8217 45033 8251 45067
rect 10425 45033 10459 45067
rect 12081 45033 12115 45067
rect 19441 45033 19475 45067
rect 25237 45033 25271 45067
rect 7297 44965 7331 44999
rect 9137 44965 9171 44999
rect 11069 44965 11103 44999
rect 18245 44965 18279 44999
rect 22201 44897 22235 44931
rect 5917 44829 5951 44863
rect 8033 44829 8067 44863
rect 13369 44829 13403 44863
rect 15301 44829 15335 44863
rect 18889 44829 18923 44863
rect 21189 44829 21223 44863
rect 24593 44829 24627 44863
rect 6745 44761 6779 44795
rect 7481 44761 7515 44795
rect 9321 44761 9355 44795
rect 9689 44761 9723 44795
rect 10057 44761 10091 44795
rect 10517 44761 10551 44795
rect 11253 44761 11287 44795
rect 11713 44761 11747 44795
rect 12173 44761 12207 44795
rect 15577 44761 15611 44795
rect 20913 44761 20947 44795
rect 22477 44761 22511 44795
rect 12725 44693 12759 44727
rect 17049 44693 17083 44727
rect 21833 44693 21867 44727
rect 23949 44693 23983 44727
rect 9137 44489 9171 44523
rect 9689 44489 9723 44523
rect 11897 44489 11931 44523
rect 12265 44489 12299 44523
rect 21373 44489 21407 44523
rect 22477 44489 22511 44523
rect 22569 44489 22603 44523
rect 6561 44421 6595 44455
rect 10885 44421 10919 44455
rect 6193 44353 6227 44387
rect 6745 44353 6779 44387
rect 8769 44353 8803 44387
rect 9229 44353 9263 44387
rect 11069 44353 11103 44387
rect 16037 44353 16071 44387
rect 19073 44353 19107 44387
rect 20729 44353 20763 44387
rect 23305 44353 23339 44387
rect 12357 44285 12391 44319
rect 12449 44285 12483 44319
rect 13185 44285 13219 44319
rect 13461 44285 13495 44319
rect 16313 44285 16347 44319
rect 16865 44285 16899 44319
rect 17141 44285 17175 44319
rect 22753 44285 22787 44319
rect 24501 44285 24535 44319
rect 24777 44285 24811 44319
rect 11621 44217 11655 44251
rect 7205 44149 7239 44183
rect 14933 44149 14967 44183
rect 15393 44149 15427 44183
rect 18613 44149 18647 44183
rect 19717 44149 19751 44183
rect 22109 44149 22143 44183
rect 23949 44149 23983 44183
rect 8033 43945 8067 43979
rect 8585 43945 8619 43979
rect 9965 43945 9999 43979
rect 15393 43945 15427 43979
rect 23489 43945 23523 43979
rect 10241 43877 10275 43911
rect 11989 43877 12023 43911
rect 9321 43809 9355 43843
rect 9505 43809 9539 43843
rect 12633 43809 12667 43843
rect 15945 43809 15979 43843
rect 17693 43809 17727 43843
rect 17785 43809 17819 43843
rect 18521 43809 18555 43843
rect 21189 43809 21223 43843
rect 22109 43809 22143 43843
rect 23121 43809 23155 43843
rect 8401 43741 8435 43775
rect 14289 43741 14323 43775
rect 15761 43741 15795 43775
rect 21465 43741 21499 43775
rect 22293 43741 22327 43775
rect 24593 43741 24627 43775
rect 9597 43673 9631 43707
rect 12449 43673 12483 43707
rect 17601 43673 17635 43707
rect 23765 43673 23799 43707
rect 24133 43673 24167 43707
rect 12357 43605 12391 43639
rect 14933 43605 14967 43639
rect 15853 43605 15887 43639
rect 17233 43605 17267 43639
rect 18245 43605 18279 43639
rect 19717 43605 19751 43639
rect 22201 43605 22235 43639
rect 22661 43605 22695 43639
rect 25237 43605 25271 43639
rect 8125 43401 8159 43435
rect 15393 43401 15427 43435
rect 17233 43401 17267 43435
rect 22293 43401 22327 43435
rect 13001 43333 13035 43367
rect 24961 43333 24995 43367
rect 1685 43265 1719 43299
rect 2145 43265 2179 43299
rect 7941 43265 7975 43299
rect 10425 43265 10459 43299
rect 16037 43265 16071 43299
rect 17325 43265 17359 43299
rect 19901 43265 19935 43299
rect 20361 43265 20395 43299
rect 22385 43265 22419 43299
rect 10149 43197 10183 43231
rect 11161 43197 11195 43231
rect 12725 43197 12759 43231
rect 15485 43197 15519 43231
rect 15577 43197 15611 43231
rect 17141 43197 17175 43231
rect 19625 43197 19659 43231
rect 22201 43197 22235 43231
rect 25237 43197 25271 43231
rect 1869 43129 1903 43163
rect 14473 43129 14507 43163
rect 16221 43129 16255 43163
rect 17693 43129 17727 43163
rect 22753 43129 22787 43163
rect 8677 43061 8711 43095
rect 15025 43061 15059 43095
rect 18153 43061 18187 43095
rect 21005 43061 21039 43095
rect 21373 43061 21407 43095
rect 21649 43061 21683 43095
rect 23121 43061 23155 43095
rect 23489 43061 23523 43095
rect 15190 42857 15224 42891
rect 22556 42857 22590 42891
rect 24593 42857 24627 42891
rect 4721 42721 4755 42755
rect 5733 42721 5767 42755
rect 9689 42721 9723 42755
rect 11069 42721 11103 42755
rect 12817 42721 12851 42755
rect 16681 42721 16715 42755
rect 17785 42721 17819 42755
rect 19717 42721 19751 42755
rect 19901 42721 19935 42755
rect 21189 42721 21223 42755
rect 21281 42721 21315 42755
rect 22293 42721 22327 42755
rect 8585 42653 8619 42687
rect 14933 42653 14967 42687
rect 17601 42653 17635 42687
rect 18337 42653 18371 42687
rect 21373 42653 21407 42687
rect 25237 42653 25271 42687
rect 4905 42585 4939 42619
rect 5917 42585 5951 42619
rect 10241 42585 10275 42619
rect 10517 42585 10551 42619
rect 11345 42585 11379 42619
rect 17509 42585 17543 42619
rect 18245 42585 18279 42619
rect 5273 42517 5307 42551
rect 6377 42517 6411 42551
rect 7941 42517 7975 42551
rect 9137 42517 9171 42551
rect 9505 42517 9539 42551
rect 9597 42517 9631 42551
rect 13369 42517 13403 42551
rect 13921 42517 13955 42551
rect 17141 42517 17175 42551
rect 19993 42517 20027 42551
rect 20361 42517 20395 42551
rect 21741 42517 21775 42551
rect 24041 42517 24075 42551
rect 4997 42313 5031 42347
rect 9597 42313 9631 42347
rect 11713 42313 11747 42347
rect 13369 42313 13403 42347
rect 13737 42313 13771 42347
rect 17141 42313 17175 42347
rect 17601 42313 17635 42347
rect 18429 42313 18463 42347
rect 25145 42313 25179 42347
rect 3433 42245 3467 42279
rect 4169 42245 4203 42279
rect 15117 42245 15151 42279
rect 24409 42245 24443 42279
rect 3617 42177 3651 42211
rect 4353 42177 4387 42211
rect 5089 42177 5123 42211
rect 7849 42177 7883 42211
rect 10057 42177 10091 42211
rect 12081 42177 12115 42211
rect 14841 42177 14875 42211
rect 16129 42177 16163 42211
rect 17509 42177 17543 42211
rect 20821 42177 20855 42211
rect 21465 42177 21499 42211
rect 22569 42177 22603 42211
rect 25329 42177 25363 42211
rect 3157 42109 3191 42143
rect 8125 42109 8159 42143
rect 12173 42109 12207 42143
rect 12265 42109 12299 42143
rect 13185 42109 13219 42143
rect 13277 42109 13311 42143
rect 16865 42109 16899 42143
rect 17693 42109 17727 42143
rect 18705 42109 18739 42143
rect 18981 42109 19015 42143
rect 22201 42109 22235 42143
rect 24685 42109 24719 42143
rect 21281 42041 21315 42075
rect 5549 41973 5583 42007
rect 10701 41973 10735 42007
rect 14197 41973 14231 42007
rect 15485 41973 15519 42007
rect 18153 41973 18187 42007
rect 20453 41973 20487 42007
rect 20913 41973 20947 42007
rect 22937 41973 22971 42007
rect 4077 41769 4111 41803
rect 8033 41769 8067 41803
rect 9413 41769 9447 41803
rect 11529 41769 11563 41803
rect 18705 41769 18739 41803
rect 4537 41701 4571 41735
rect 8309 41701 8343 41735
rect 24041 41701 24075 41735
rect 6285 41633 6319 41667
rect 14565 41633 14599 41667
rect 16037 41633 16071 41667
rect 16957 41633 16991 41667
rect 17049 41633 17083 41667
rect 19533 41633 19567 41667
rect 22201 41633 22235 41667
rect 23397 41633 23431 41667
rect 25053 41633 25087 41667
rect 25145 41633 25179 41667
rect 11161 41565 11195 41599
rect 12909 41565 12943 41599
rect 14289 41565 14323 41599
rect 17693 41565 17727 41599
rect 20821 41565 20855 41599
rect 23213 41565 23247 41599
rect 4721 41497 4755 41531
rect 5089 41497 5123 41531
rect 6561 41497 6595 41531
rect 10885 41497 10919 41531
rect 12081 41497 12115 41531
rect 18981 41497 19015 41531
rect 20361 41497 20395 41531
rect 21465 41497 21499 41531
rect 23305 41497 23339 41531
rect 13369 41429 13403 41463
rect 16497 41429 16531 41463
rect 16865 41429 16899 41463
rect 18337 41429 18371 41463
rect 21005 41429 21039 41463
rect 22845 41429 22879 41463
rect 24225 41429 24259 41463
rect 24593 41429 24627 41463
rect 24961 41429 24995 41463
rect 10885 41225 10919 41259
rect 11345 41225 11379 41259
rect 13277 41225 13311 41259
rect 15761 41225 15795 41259
rect 17141 41225 17175 41259
rect 18521 41225 18555 41259
rect 19901 41225 19935 41259
rect 20637 41225 20671 41259
rect 22661 41225 22695 41259
rect 22753 41225 22787 41259
rect 23121 41225 23155 41259
rect 10425 41157 10459 41191
rect 1593 41089 1627 41123
rect 2053 41089 2087 41123
rect 9689 41089 9723 41123
rect 12081 41089 12115 41123
rect 12817 41089 12851 41123
rect 15025 41089 15059 41123
rect 15853 41089 15887 41123
rect 17233 41089 17267 41123
rect 18613 41089 18647 41123
rect 19809 41089 19843 41123
rect 21005 41089 21039 41123
rect 24501 41089 24535 41123
rect 24777 41089 24811 41123
rect 8125 41021 8159 41055
rect 8401 41021 8435 41055
rect 8769 41021 8803 41055
rect 12173 41021 12207 41055
rect 12265 41021 12299 41055
rect 14749 41021 14783 41055
rect 15577 41021 15611 41055
rect 17049 41021 17083 41055
rect 18337 41021 18371 41055
rect 19993 41021 20027 41055
rect 21097 41021 21131 41055
rect 21281 41021 21315 41055
rect 22569 41021 22603 41055
rect 23765 41021 23799 41055
rect 8861 40953 8895 40987
rect 11713 40953 11747 40987
rect 17969 40953 18003 40987
rect 1777 40885 1811 40919
rect 6653 40885 6687 40919
rect 9137 40885 9171 40919
rect 11069 40885 11103 40919
rect 16221 40885 16255 40919
rect 17601 40885 17635 40919
rect 18981 40885 19015 40919
rect 19441 40885 19475 40919
rect 21833 40885 21867 40919
rect 22109 40885 22143 40919
rect 23489 40885 23523 40919
rect 8401 40681 8435 40715
rect 13921 40681 13955 40715
rect 15853 40681 15887 40715
rect 21925 40681 21959 40715
rect 23857 40613 23891 40647
rect 9321 40545 9355 40579
rect 10977 40545 11011 40579
rect 11713 40545 11747 40579
rect 12909 40545 12943 40579
rect 13093 40545 13127 40579
rect 15209 40545 15243 40579
rect 16313 40545 16347 40579
rect 16405 40545 16439 40579
rect 17141 40545 17175 40579
rect 18613 40545 18647 40579
rect 18889 40545 18923 40579
rect 21281 40545 21315 40579
rect 22661 40545 22695 40579
rect 7757 40477 7791 40511
rect 11989 40477 12023 40511
rect 13185 40477 13219 40511
rect 21189 40477 21223 40511
rect 22109 40477 22143 40511
rect 22937 40477 22971 40511
rect 24041 40477 24075 40511
rect 24593 40477 24627 40511
rect 9597 40409 9631 40443
rect 10793 40409 10827 40443
rect 11897 40409 11931 40443
rect 14473 40409 14507 40443
rect 16221 40409 16255 40443
rect 20361 40409 20395 40443
rect 22845 40409 22879 40443
rect 8769 40341 8803 40375
rect 9505 40341 9539 40375
rect 9965 40341 9999 40375
rect 10425 40341 10459 40375
rect 10885 40341 10919 40375
rect 12357 40341 12391 40375
rect 13553 40341 13587 40375
rect 20729 40341 20763 40375
rect 21097 40341 21131 40375
rect 23305 40341 23339 40375
rect 25237 40341 25271 40375
rect 13461 40137 13495 40171
rect 15301 40137 15335 40171
rect 16865 40137 16899 40171
rect 19533 40137 19567 40171
rect 19993 40137 20027 40171
rect 22385 40137 22419 40171
rect 22753 40137 22787 40171
rect 8861 40069 8895 40103
rect 11989 40069 12023 40103
rect 13829 40069 13863 40103
rect 14933 40069 14967 40103
rect 15761 40069 15795 40103
rect 17233 40069 17267 40103
rect 18061 40069 18095 40103
rect 19625 40069 19659 40103
rect 10885 40001 10919 40035
rect 11713 40001 11747 40035
rect 17325 40001 17359 40035
rect 21189 40001 21223 40035
rect 21465 40001 21499 40035
rect 25329 40001 25363 40035
rect 10609 39933 10643 39967
rect 14749 39933 14783 39967
rect 14841 39933 14875 39967
rect 17509 39933 17543 39967
rect 19349 39933 19383 39967
rect 22109 39933 22143 39967
rect 22293 39933 22327 39967
rect 23581 39933 23615 39967
rect 25053 39933 25087 39967
rect 21557 39865 21591 39899
rect 11253 39797 11287 39831
rect 14197 39797 14231 39831
rect 16313 39797 16347 39831
rect 20269 39797 20303 39831
rect 23121 39797 23155 39831
rect 7205 39593 7239 39627
rect 7573 39593 7607 39627
rect 9137 39593 9171 39627
rect 10241 39593 10275 39627
rect 11529 39593 11563 39627
rect 17141 39593 17175 39627
rect 25329 39593 25363 39627
rect 11897 39525 11931 39559
rect 15117 39525 15151 39559
rect 18705 39525 18739 39559
rect 9689 39457 9723 39491
rect 10977 39457 11011 39491
rect 12909 39457 12943 39491
rect 15761 39457 15795 39491
rect 16589 39457 16623 39491
rect 20269 39457 20303 39491
rect 20453 39457 20487 39491
rect 24041 39457 24075 39491
rect 5457 39389 5491 39423
rect 11161 39389 11195 39423
rect 12725 39389 12759 39423
rect 17785 39389 17819 39423
rect 20545 39389 20579 39423
rect 24685 39389 24719 39423
rect 5733 39321 5767 39355
rect 12633 39321 12667 39355
rect 16773 39321 16807 39355
rect 19441 39321 19475 39355
rect 23765 39321 23799 39355
rect 8585 39253 8619 39287
rect 9505 39253 9539 39287
rect 9597 39253 9631 39287
rect 10517 39253 10551 39287
rect 11069 39253 11103 39287
rect 12265 39253 12299 39287
rect 13277 39253 13311 39287
rect 15485 39253 15519 39287
rect 15577 39253 15611 39287
rect 16681 39253 16715 39287
rect 18429 39253 18463 39287
rect 20913 39253 20947 39287
rect 21649 39253 21683 39287
rect 22293 39253 22327 39287
rect 5365 39049 5399 39083
rect 6561 39049 6595 39083
rect 8033 39049 8067 39083
rect 8677 39049 8711 39083
rect 8769 39049 8803 39083
rect 9137 39049 9171 39083
rect 10425 39049 10459 39083
rect 17417 39049 17451 39083
rect 19257 39049 19291 39083
rect 20361 39049 20395 39083
rect 23581 39049 23615 39083
rect 10793 38981 10827 39015
rect 13921 38981 13955 39015
rect 15393 38981 15427 39015
rect 17785 38981 17819 39015
rect 22385 38981 22419 39015
rect 23489 38981 23523 39015
rect 25329 38981 25363 39015
rect 6009 38913 6043 38947
rect 6929 38913 6963 38947
rect 10885 38913 10919 38947
rect 14197 38913 14231 38947
rect 15485 38913 15519 38947
rect 16037 38913 16071 38947
rect 17877 38913 17911 38947
rect 18429 38913 18463 38947
rect 20453 38913 20487 38947
rect 21465 38913 21499 38947
rect 7021 38845 7055 38879
rect 7113 38845 7147 38879
rect 8585 38845 8619 38879
rect 9965 38845 9999 38879
rect 10977 38845 11011 38879
rect 11713 38845 11747 38879
rect 15577 38845 15611 38879
rect 17969 38845 18003 38879
rect 19073 38845 19107 38879
rect 19165 38845 19199 38879
rect 20177 38845 20211 38879
rect 22477 38845 22511 38879
rect 22661 38845 22695 38879
rect 23397 38845 23431 38879
rect 24593 38845 24627 38879
rect 12449 38777 12483 38811
rect 17049 38777 17083 38811
rect 19625 38777 19659 38811
rect 14473 38709 14507 38743
rect 15025 38709 15059 38743
rect 16221 38709 16255 38743
rect 20821 38709 20855 38743
rect 21281 38709 21315 38743
rect 22017 38709 22051 38743
rect 23949 38709 23983 38743
rect 10517 38505 10551 38539
rect 11713 38505 11747 38539
rect 18153 38505 18187 38539
rect 19441 38505 19475 38539
rect 24041 38505 24075 38539
rect 24593 38505 24627 38539
rect 12725 38437 12759 38471
rect 14749 38437 14783 38471
rect 21189 38437 21223 38471
rect 5641 38369 5675 38403
rect 7389 38369 7423 38403
rect 9873 38369 9907 38403
rect 11069 38369 11103 38403
rect 13277 38369 13311 38403
rect 13829 38369 13863 38403
rect 15669 38369 15703 38403
rect 16313 38369 16347 38403
rect 16497 38369 16531 38403
rect 17509 38369 17543 38403
rect 17693 38369 17727 38403
rect 18429 38369 18463 38403
rect 19993 38369 20027 38403
rect 21925 38369 21959 38403
rect 22109 38369 22143 38403
rect 23213 38369 23247 38403
rect 23305 38369 23339 38403
rect 1593 38301 1627 38335
rect 2053 38301 2087 38335
rect 7849 38301 7883 38335
rect 9505 38301 9539 38335
rect 10149 38301 10183 38335
rect 11345 38301 11379 38335
rect 17785 38301 17819 38335
rect 18981 38301 19015 38335
rect 19901 38301 19935 38335
rect 21373 38301 21407 38335
rect 22201 38301 22235 38335
rect 25237 38301 25271 38335
rect 5917 38233 5951 38267
rect 12449 38233 12483 38267
rect 13185 38233 13219 38267
rect 16589 38233 16623 38267
rect 19809 38233 19843 38267
rect 20913 38233 20947 38267
rect 1777 38165 1811 38199
rect 8493 38165 8527 38199
rect 9321 38165 9355 38199
rect 10057 38165 10091 38199
rect 11253 38165 11287 38199
rect 13093 38165 13127 38199
rect 15025 38165 15059 38199
rect 15393 38165 15427 38199
rect 15485 38165 15519 38199
rect 16957 38165 16991 38199
rect 18705 38165 18739 38199
rect 20545 38165 20579 38199
rect 22569 38165 22603 38199
rect 23397 38165 23431 38199
rect 23765 38165 23799 38199
rect 6009 37961 6043 37995
rect 8861 37961 8895 37995
rect 9965 37961 9999 37995
rect 10609 37961 10643 37995
rect 12081 37961 12115 37995
rect 16129 37961 16163 37995
rect 16865 37961 16899 37995
rect 19073 37961 19107 37995
rect 19533 37961 19567 37995
rect 20637 37961 20671 37995
rect 21005 37961 21039 37995
rect 21281 37961 21315 37995
rect 24409 37961 24443 37995
rect 8309 37893 8343 37927
rect 12173 37893 12207 37927
rect 18337 37893 18371 37927
rect 20545 37893 20579 37927
rect 4261 37825 4295 37859
rect 9873 37825 9907 37859
rect 13553 37825 13587 37859
rect 15301 37825 15335 37859
rect 19441 37825 19475 37859
rect 21465 37825 21499 37859
rect 22201 37825 22235 37859
rect 25329 37825 25363 37859
rect 4537 37757 4571 37791
rect 6561 37757 6595 37791
rect 8585 37757 8619 37791
rect 10057 37757 10091 37791
rect 12265 37757 12299 37791
rect 14013 37757 14047 37791
rect 14657 37757 14691 37791
rect 15393 37757 15427 37791
rect 15577 37757 15611 37791
rect 18613 37757 18647 37791
rect 19625 37757 19659 37791
rect 20453 37757 20487 37791
rect 22661 37757 22695 37791
rect 22937 37757 22971 37791
rect 24685 37757 24719 37791
rect 11253 37689 11287 37723
rect 12909 37689 12943 37723
rect 9505 37621 9539 37655
rect 11713 37621 11747 37655
rect 14933 37621 14967 37655
rect 22017 37621 22051 37655
rect 25145 37621 25179 37655
rect 8217 37417 8251 37451
rect 14473 37417 14507 37451
rect 16129 37417 16163 37451
rect 20821 37417 20855 37451
rect 21097 37417 21131 37451
rect 23949 37417 23983 37451
rect 24225 37417 24259 37451
rect 15853 37349 15887 37383
rect 7573 37281 7607 37315
rect 9229 37281 9263 37315
rect 11069 37281 11103 37315
rect 13185 37281 13219 37315
rect 14105 37281 14139 37315
rect 15301 37281 15335 37315
rect 16681 37281 16715 37315
rect 18613 37281 18647 37315
rect 20729 37281 20763 37315
rect 7757 37213 7791 37247
rect 10057 37213 10091 37247
rect 12541 37213 12575 37247
rect 13277 37213 13311 37247
rect 13369 37213 13403 37247
rect 15117 37213 15151 37247
rect 18429 37213 18463 37247
rect 20361 37213 20395 37247
rect 21465 37213 21499 37247
rect 22845 37213 22879 37247
rect 24593 37213 24627 37247
rect 10977 37145 11011 37179
rect 15209 37145 15243 37179
rect 16497 37145 16531 37179
rect 19533 37145 19567 37179
rect 22293 37145 22327 37179
rect 7849 37077 7883 37111
rect 10517 37077 10551 37111
rect 10885 37077 10919 37111
rect 11897 37077 11931 37111
rect 13737 37077 13771 37111
rect 14749 37077 14783 37111
rect 16589 37077 16623 37111
rect 17325 37077 17359 37111
rect 18061 37077 18095 37111
rect 18521 37077 18555 37111
rect 23489 37077 23523 37111
rect 25237 37077 25271 37111
rect 7481 36873 7515 36907
rect 11529 36873 11563 36907
rect 15945 36873 15979 36907
rect 16405 36873 16439 36907
rect 17141 36873 17175 36907
rect 17233 36873 17267 36907
rect 17601 36873 17635 36907
rect 20637 36873 20671 36907
rect 21465 36873 21499 36907
rect 22293 36873 22327 36907
rect 22753 36873 22787 36907
rect 23581 36873 23615 36907
rect 8953 36805 8987 36839
rect 9505 36805 9539 36839
rect 11161 36805 11195 36839
rect 15117 36805 15151 36839
rect 20729 36805 20763 36839
rect 21281 36805 21315 36839
rect 23029 36805 23063 36839
rect 25053 36805 25087 36839
rect 9229 36737 9263 36771
rect 13001 36737 13035 36771
rect 13645 36737 13679 36771
rect 15025 36737 15059 36771
rect 19349 36737 19383 36771
rect 22385 36737 22419 36771
rect 10333 36669 10367 36703
rect 11989 36669 12023 36703
rect 13093 36669 13127 36703
rect 13185 36669 13219 36703
rect 15209 36669 15243 36703
rect 17049 36669 17083 36703
rect 19441 36669 19475 36703
rect 19533 36669 19567 36703
rect 20821 36669 20855 36703
rect 22109 36669 22143 36703
rect 25329 36669 25363 36703
rect 18981 36601 19015 36635
rect 12173 36533 12207 36567
rect 12265 36533 12299 36567
rect 12633 36533 12667 36567
rect 14657 36533 14691 36567
rect 15761 36533 15795 36567
rect 20269 36533 20303 36567
rect 23213 36533 23247 36567
rect 9505 36329 9539 36363
rect 13185 36329 13219 36363
rect 15025 36329 15059 36363
rect 16957 36329 16991 36363
rect 8401 36193 8435 36227
rect 10057 36193 10091 36227
rect 12541 36193 12575 36227
rect 14473 36193 14507 36227
rect 19901 36193 19935 36227
rect 19993 36193 20027 36227
rect 21281 36193 21315 36227
rect 21373 36193 21407 36227
rect 22293 36193 22327 36227
rect 25145 36193 25179 36227
rect 1593 36125 1627 36159
rect 2053 36125 2087 36159
rect 6653 36125 6687 36159
rect 9965 36125 9999 36159
rect 11989 36125 12023 36159
rect 12817 36125 12851 36159
rect 17509 36125 17543 36159
rect 21189 36125 21223 36159
rect 25053 36125 25087 36159
rect 6929 36057 6963 36091
rect 9873 36057 9907 36091
rect 14657 36057 14691 36091
rect 15485 36057 15519 36091
rect 19809 36057 19843 36091
rect 22569 36057 22603 36091
rect 24961 36057 24995 36091
rect 1777 35989 1811 36023
rect 11345 35989 11379 36023
rect 12725 35989 12759 36023
rect 13921 35989 13955 36023
rect 14565 35989 14599 36023
rect 18153 35989 18187 36023
rect 19441 35989 19475 36023
rect 20821 35989 20855 36023
rect 24041 35989 24075 36023
rect 24593 35989 24627 36023
rect 7389 35785 7423 35819
rect 11713 35785 11747 35819
rect 13829 35785 13863 35819
rect 6469 35717 6503 35751
rect 18153 35717 18187 35751
rect 4261 35649 4295 35683
rect 8033 35649 8067 35683
rect 8493 35649 8527 35683
rect 17877 35649 17911 35683
rect 4537 35581 4571 35615
rect 6009 35581 6043 35615
rect 8769 35581 8803 35615
rect 13185 35581 13219 35615
rect 13461 35581 13495 35615
rect 22661 35581 22695 35615
rect 24685 35581 24719 35615
rect 24961 35581 24995 35615
rect 25329 35581 25363 35615
rect 7021 35445 7055 35479
rect 10241 35445 10275 35479
rect 19625 35445 19659 35479
rect 23213 35445 23247 35479
rect 25421 35445 25455 35479
rect 5549 35241 5583 35275
rect 7849 35241 7883 35275
rect 8953 35241 8987 35275
rect 9321 35241 9355 35275
rect 13093 35241 13127 35275
rect 15485 35241 15519 35275
rect 23949 35241 23983 35275
rect 25237 35241 25271 35275
rect 7297 35105 7331 35139
rect 8401 35105 8435 35139
rect 9781 35105 9815 35139
rect 9965 35105 9999 35139
rect 12357 35105 12391 35139
rect 17233 35105 17267 35139
rect 22201 35105 22235 35139
rect 23397 35105 23431 35139
rect 8309 35037 8343 35071
rect 13737 35037 13771 35071
rect 18245 35037 18279 35071
rect 19441 35037 19475 35071
rect 22385 35037 22419 35071
rect 23581 35037 23615 35071
rect 24593 35037 24627 35071
rect 7021 34969 7055 35003
rect 8217 34969 8251 35003
rect 12081 34969 12115 35003
rect 16957 34969 16991 35003
rect 18889 34969 18923 35003
rect 19717 34969 19751 35003
rect 23489 34969 23523 35003
rect 9689 34901 9723 34935
rect 10609 34901 10643 34935
rect 12725 34901 12759 34935
rect 14105 34901 14139 34935
rect 21189 34901 21223 34935
rect 22293 34901 22327 34935
rect 22753 34901 22787 34935
rect 4905 34697 4939 34731
rect 5549 34697 5583 34731
rect 6009 34697 6043 34731
rect 8861 34697 8895 34731
rect 10977 34697 11011 34731
rect 11253 34697 11287 34731
rect 13921 34697 13955 34731
rect 14381 34697 14415 34731
rect 17233 34697 17267 34731
rect 18337 34697 18371 34731
rect 18705 34697 18739 34731
rect 20637 34697 20671 34731
rect 22477 34697 22511 34731
rect 23213 34697 23247 34731
rect 23949 34697 23983 34731
rect 24593 34697 24627 34731
rect 11989 34629 12023 34663
rect 21833 34629 21867 34663
rect 5641 34561 5675 34595
rect 10609 34561 10643 34595
rect 11713 34561 11747 34595
rect 14289 34561 14323 34595
rect 17877 34561 17911 34595
rect 19349 34561 19383 34595
rect 19533 34561 19567 34595
rect 20177 34561 20211 34595
rect 20269 34561 20303 34595
rect 22569 34561 22603 34595
rect 23765 34561 23799 34595
rect 24409 34561 24443 34595
rect 25329 34561 25363 34595
rect 5457 34493 5491 34527
rect 6561 34493 6595 34527
rect 6837 34493 6871 34527
rect 8309 34493 8343 34527
rect 10333 34493 10367 34527
rect 11161 34493 11195 34527
rect 13461 34493 13495 34527
rect 14473 34493 14507 34527
rect 18797 34493 18831 34527
rect 18889 34493 18923 34527
rect 20085 34493 20119 34527
rect 20913 34493 20947 34527
rect 22293 34493 22327 34527
rect 22937 34425 22971 34459
rect 25145 34357 25179 34391
rect 7113 34153 7147 34187
rect 7941 34153 7975 34187
rect 9137 34153 9171 34187
rect 10425 34153 10459 34187
rect 11069 34153 11103 34187
rect 14289 34153 14323 34187
rect 17325 34153 17359 34187
rect 20361 34153 20395 34187
rect 23857 34153 23891 34187
rect 24501 34153 24535 34187
rect 5825 34017 5859 34051
rect 9689 34017 9723 34051
rect 11529 34017 11563 34051
rect 11621 34017 11655 34051
rect 13553 34017 13587 34051
rect 14841 34017 14875 34051
rect 19809 34017 19843 34051
rect 21465 34017 21499 34051
rect 6469 33949 6503 33983
rect 8585 33949 8619 33983
rect 10609 33949 10643 33983
rect 15577 33949 15611 33983
rect 21281 33949 21315 33983
rect 22017 33949 22051 33983
rect 24041 33949 24075 33983
rect 24869 33949 24903 33983
rect 25329 33949 25363 33983
rect 9597 33881 9631 33915
rect 13461 33881 13495 33915
rect 15853 33881 15887 33915
rect 19993 33881 20027 33915
rect 21189 33881 21223 33915
rect 9505 33813 9539 33847
rect 11437 33813 11471 33847
rect 13001 33813 13035 33847
rect 13369 33813 13403 33847
rect 14657 33813 14691 33847
rect 14749 33813 14783 33847
rect 19349 33813 19383 33847
rect 19901 33813 19935 33847
rect 20821 33813 20855 33847
rect 22661 33813 22695 33847
rect 23121 33813 23155 33847
rect 25145 33813 25179 33847
rect 7665 33609 7699 33643
rect 8309 33609 8343 33643
rect 8769 33609 8803 33643
rect 10517 33609 10551 33643
rect 11713 33609 11747 33643
rect 12173 33609 12207 33643
rect 15117 33609 15151 33643
rect 16037 33609 16071 33643
rect 22385 33609 22419 33643
rect 25237 33609 25271 33643
rect 15945 33541 15979 33575
rect 19533 33541 19567 33575
rect 20453 33541 20487 33575
rect 1593 33473 1627 33507
rect 2053 33473 2087 33507
rect 8401 33473 8435 33507
rect 10149 33473 10183 33507
rect 10977 33473 11011 33507
rect 12081 33473 12115 33507
rect 14473 33473 14507 33507
rect 21097 33473 21131 33507
rect 8217 33405 8251 33439
rect 9873 33405 9907 33439
rect 10057 33405 10091 33439
rect 12265 33405 12299 33439
rect 16129 33405 16163 33439
rect 19809 33405 19843 33439
rect 22477 33405 22511 33439
rect 22569 33405 22603 33439
rect 23489 33405 23523 33439
rect 23765 33405 23799 33439
rect 13921 33337 13955 33371
rect 23029 33337 23063 33371
rect 1777 33269 1811 33303
rect 9045 33269 9079 33303
rect 14105 33269 14139 33303
rect 15577 33269 15611 33303
rect 18061 33269 18095 33303
rect 22017 33269 22051 33303
rect 7573 33065 7607 33099
rect 7941 33065 7975 33099
rect 16405 33065 16439 33099
rect 17785 33065 17819 33099
rect 23489 33065 23523 33099
rect 23857 33065 23891 33099
rect 25145 33065 25179 33099
rect 20637 32997 20671 33031
rect 23029 32997 23063 33031
rect 6101 32929 6135 32963
rect 8401 32929 8435 32963
rect 16957 32929 16991 32963
rect 19993 32929 20027 32963
rect 21373 32929 21407 32963
rect 5825 32861 5859 32895
rect 9137 32861 9171 32895
rect 16037 32861 16071 32895
rect 17141 32861 17175 32895
rect 20453 32861 20487 32895
rect 21465 32861 21499 32895
rect 22385 32861 22419 32895
rect 23213 32861 23247 32895
rect 24041 32861 24075 32895
rect 24869 32861 24903 32895
rect 25329 32861 25363 32895
rect 15761 32793 15795 32827
rect 21557 32793 21591 32827
rect 24501 32793 24535 32827
rect 9781 32725 9815 32759
rect 14289 32725 14323 32759
rect 17049 32725 17083 32759
rect 17509 32725 17543 32759
rect 21925 32725 21959 32759
rect 22569 32725 22603 32759
rect 24685 32725 24719 32759
rect 12081 32521 12115 32555
rect 12633 32521 12667 32555
rect 13093 32521 13127 32555
rect 14473 32521 14507 32555
rect 18061 32521 18095 32555
rect 20453 32521 20487 32555
rect 21465 32521 21499 32555
rect 22477 32521 22511 32555
rect 24133 32521 24167 32555
rect 8309 32453 8343 32487
rect 10241 32453 10275 32487
rect 14381 32453 14415 32487
rect 17969 32453 18003 32487
rect 20361 32453 20395 32487
rect 12725 32385 12759 32419
rect 15945 32385 15979 32419
rect 19165 32385 19199 32419
rect 21281 32385 21315 32419
rect 23489 32385 23523 32419
rect 24685 32385 24719 32419
rect 7573 32317 7607 32351
rect 8033 32317 8067 32351
rect 12541 32317 12575 32351
rect 14197 32317 14231 32351
rect 18153 32317 18187 32351
rect 19257 32317 19291 32351
rect 19441 32317 19475 32351
rect 20545 32317 20579 32351
rect 22201 32317 22235 32351
rect 22385 32317 22419 32351
rect 25237 32317 25271 32351
rect 9781 32249 9815 32283
rect 14841 32181 14875 32215
rect 15301 32181 15335 32215
rect 17601 32181 17635 32215
rect 18797 32181 18831 32215
rect 19993 32181 20027 32215
rect 22845 32181 22879 32215
rect 6653 31977 6687 32011
rect 8769 31977 8803 32011
rect 11621 31977 11655 32011
rect 14289 31977 14323 32011
rect 15485 31977 15519 32011
rect 19441 31977 19475 32011
rect 19809 31977 19843 32011
rect 20637 31977 20671 32011
rect 21649 31977 21683 32011
rect 22556 31977 22590 32011
rect 24041 31977 24075 32011
rect 13829 31909 13863 31943
rect 21925 31909 21959 31943
rect 8401 31841 8435 31875
rect 9873 31841 9907 31875
rect 12817 31841 12851 31875
rect 14841 31841 14875 31875
rect 16957 31841 16991 31875
rect 18337 31841 18371 31875
rect 19625 31841 19659 31875
rect 21097 31841 21131 31875
rect 21189 31841 21223 31875
rect 22293 31841 22327 31875
rect 11897 31773 11931 31807
rect 13645 31773 13679 31807
rect 14749 31773 14783 31807
rect 17233 31773 17267 31807
rect 17693 31773 17727 31807
rect 24593 31773 24627 31807
rect 8125 31705 8159 31739
rect 10149 31705 10183 31739
rect 9137 31637 9171 31671
rect 14657 31637 14691 31671
rect 21281 31637 21315 31671
rect 25237 31637 25271 31671
rect 7849 31433 7883 31467
rect 16313 31433 16347 31467
rect 18337 31433 18371 31467
rect 19901 31433 19935 31467
rect 21097 31433 21131 31467
rect 21189 31433 21223 31467
rect 16037 31365 16071 31399
rect 19993 31365 20027 31399
rect 22293 31365 22327 31399
rect 23121 31365 23155 31399
rect 24961 31365 24995 31399
rect 3801 31297 3835 31331
rect 10517 31297 10551 31331
rect 12633 31297 12667 31331
rect 15209 31297 15243 31331
rect 15301 31297 15335 31331
rect 17233 31297 17267 31331
rect 18705 31297 18739 31331
rect 18797 31297 18831 31331
rect 22385 31297 22419 31331
rect 25237 31297 25271 31331
rect 3985 31229 4019 31263
rect 4905 31229 4939 31263
rect 7205 31229 7239 31263
rect 7665 31229 7699 31263
rect 7757 31229 7791 31263
rect 12909 31229 12943 31263
rect 15485 31229 15519 31263
rect 17325 31229 17359 31263
rect 17417 31229 17451 31263
rect 18889 31229 18923 31263
rect 20085 31229 20119 31263
rect 21281 31229 21315 31263
rect 22109 31229 22143 31263
rect 23489 31229 23523 31263
rect 6929 31161 6963 31195
rect 8217 31161 8251 31195
rect 14841 31161 14875 31195
rect 16865 31161 16899 31195
rect 11161 31093 11195 31127
rect 14381 31093 14415 31127
rect 15853 31093 15887 31127
rect 19533 31093 19567 31127
rect 20729 31093 20763 31127
rect 22753 31093 22787 31127
rect 8309 30889 8343 30923
rect 12633 30889 12667 30923
rect 17141 30889 17175 30923
rect 21557 30889 21591 30923
rect 15853 30821 15887 30855
rect 20269 30821 20303 30855
rect 7665 30753 7699 30787
rect 11161 30753 11195 30787
rect 11437 30753 11471 30787
rect 13185 30753 13219 30787
rect 13645 30753 13679 30787
rect 14657 30753 14691 30787
rect 16497 30753 16531 30787
rect 19717 30753 19751 30787
rect 23121 30753 23155 30787
rect 7941 30685 7975 30719
rect 14381 30685 14415 30719
rect 18889 30685 18923 30719
rect 20729 30685 20763 30719
rect 23213 30685 23247 30719
rect 24593 30685 24627 30719
rect 15393 30617 15427 30651
rect 18613 30617 18647 30651
rect 19809 30617 19843 30651
rect 21189 30617 21223 30651
rect 7849 30549 7883 30583
rect 9689 30549 9723 30583
rect 11897 30549 11931 30583
rect 13001 30549 13035 30583
rect 13093 30549 13127 30583
rect 15485 30549 15519 30583
rect 16221 30549 16255 30583
rect 16313 30549 16347 30583
rect 19901 30549 19935 30583
rect 20913 30549 20947 30583
rect 21925 30549 21959 30583
rect 23305 30549 23339 30583
rect 23673 30549 23707 30583
rect 24777 30549 24811 30583
rect 16773 30345 16807 30379
rect 9597 30277 9631 30311
rect 10793 30277 10827 30311
rect 12909 30277 12943 30311
rect 17049 30277 17083 30311
rect 19809 30277 19843 30311
rect 25329 30277 25363 30311
rect 9505 30209 9539 30243
rect 13001 30209 13035 30243
rect 17693 30209 17727 30243
rect 17785 30209 17819 30243
rect 18705 30209 18739 30243
rect 20453 30209 20487 30243
rect 22753 30209 22787 30243
rect 23213 30209 23247 30243
rect 23673 30209 23707 30243
rect 24501 30209 24535 30243
rect 9413 30141 9447 30175
rect 10609 30141 10643 30175
rect 10701 30141 10735 30175
rect 12725 30141 12759 30175
rect 17509 30141 17543 30175
rect 20913 30141 20947 30175
rect 9965 30073 9999 30107
rect 11161 30073 11195 30107
rect 11621 30073 11655 30107
rect 18153 30073 18187 30107
rect 23029 30073 23063 30107
rect 8677 30005 8711 30039
rect 8861 30005 8895 30039
rect 11805 30005 11839 30039
rect 12357 30005 12391 30039
rect 13369 30005 13403 30039
rect 19349 30005 19383 30039
rect 23857 30005 23891 30039
rect 8033 29801 8067 29835
rect 11897 29801 11931 29835
rect 15209 29801 15243 29835
rect 16957 29801 16991 29835
rect 22017 29801 22051 29835
rect 25421 29801 25455 29835
rect 20913 29733 20947 29767
rect 22477 29733 22511 29767
rect 24593 29733 24627 29767
rect 4077 29665 4111 29699
rect 11253 29665 11287 29699
rect 11529 29665 11563 29699
rect 18429 29665 18463 29699
rect 18705 29665 18739 29699
rect 19625 29665 19659 29699
rect 19809 29665 19843 29699
rect 21465 29665 21499 29699
rect 22937 29665 22971 29699
rect 23121 29665 23155 29699
rect 19901 29597 19935 29631
rect 21557 29597 21591 29631
rect 22845 29597 22879 29631
rect 23581 29597 23615 29631
rect 24041 29597 24075 29631
rect 24777 29597 24811 29631
rect 4261 29529 4295 29563
rect 5917 29529 5951 29563
rect 16497 29529 16531 29563
rect 9781 29461 9815 29495
rect 18981 29461 19015 29495
rect 20269 29461 20303 29495
rect 21649 29461 21683 29495
rect 23857 29461 23891 29495
rect 25053 29461 25087 29495
rect 3571 29257 3605 29291
rect 8401 29257 8435 29291
rect 8769 29257 8803 29291
rect 12725 29257 12759 29291
rect 13829 29257 13863 29291
rect 13921 29257 13955 29291
rect 15853 29257 15887 29291
rect 17969 29257 18003 29291
rect 18705 29257 18739 29291
rect 19165 29257 19199 29291
rect 21465 29257 21499 29291
rect 15761 29189 15795 29223
rect 17877 29189 17911 29223
rect 24593 29189 24627 29223
rect 24777 29189 24811 29223
rect 3500 29121 3534 29155
rect 7665 29121 7699 29155
rect 10333 29121 10367 29155
rect 12357 29121 12391 29155
rect 19073 29121 19107 29155
rect 19901 29121 19935 29155
rect 22017 29121 22051 29155
rect 23305 29121 23339 29155
rect 23949 29121 23983 29155
rect 8861 29053 8895 29087
rect 8953 29053 8987 29087
rect 12173 29053 12207 29087
rect 12265 29053 12299 29087
rect 14105 29053 14139 29087
rect 15945 29053 15979 29087
rect 18061 29053 18095 29087
rect 19349 29053 19383 29087
rect 22661 29053 22695 29087
rect 8033 28985 8067 29019
rect 11621 28985 11655 29019
rect 13461 28985 13495 29019
rect 15393 28985 15427 29019
rect 16773 28985 16807 29019
rect 23121 28985 23155 29019
rect 23765 28985 23799 29019
rect 24317 28985 24351 29019
rect 7021 28917 7055 28951
rect 9689 28917 9723 28951
rect 17509 28917 17543 28951
rect 20545 28917 20579 28951
rect 18889 28713 18923 28747
rect 4261 28577 4295 28611
rect 5733 28577 5767 28611
rect 11805 28577 11839 28611
rect 12817 28577 12851 28611
rect 14749 28577 14783 28611
rect 14841 28577 14875 28611
rect 16589 28577 16623 28611
rect 16681 28577 16715 28611
rect 18061 28577 18095 28611
rect 18245 28577 18279 28611
rect 18981 28577 19015 28611
rect 20913 28577 20947 28611
rect 8585 28509 8619 28543
rect 9781 28509 9815 28543
rect 12725 28509 12759 28543
rect 13553 28509 13587 28543
rect 16773 28509 16807 28543
rect 17969 28509 18003 28543
rect 18613 28509 18647 28543
rect 21189 28509 21223 28543
rect 22293 28509 22327 28543
rect 24685 28509 24719 28543
rect 4445 28441 4479 28475
rect 8309 28441 8343 28475
rect 9137 28441 9171 28475
rect 14657 28441 14691 28475
rect 21465 28441 21499 28475
rect 22569 28441 22603 28475
rect 24869 28441 24903 28475
rect 6837 28373 6871 28407
rect 12265 28373 12299 28407
rect 12633 28373 12667 28407
rect 13369 28373 13403 28407
rect 14289 28373 14323 28407
rect 15301 28373 15335 28407
rect 15577 28373 15611 28407
rect 17141 28373 17175 28407
rect 17601 28373 17635 28407
rect 19441 28373 19475 28407
rect 24041 28373 24075 28407
rect 8585 28169 8619 28203
rect 17049 28169 17083 28203
rect 18981 28169 19015 28203
rect 19717 28169 19751 28203
rect 22109 28169 22143 28203
rect 7113 28101 7147 28135
rect 10517 28101 10551 28135
rect 11713 28101 11747 28135
rect 13093 28101 13127 28135
rect 17785 28101 17819 28135
rect 18613 28101 18647 28135
rect 24777 28101 24811 28135
rect 12357 28033 12391 28067
rect 15669 28033 15703 28067
rect 17877 28033 17911 28067
rect 19809 28033 19843 28067
rect 21465 28033 21499 28067
rect 6837 27965 6871 27999
rect 9045 27965 9079 27999
rect 10793 27965 10827 27999
rect 12817 27965 12851 27999
rect 17693 27965 17727 27999
rect 19625 27965 19659 27999
rect 21189 27965 21223 27999
rect 23581 27965 23615 27999
rect 23857 27965 23891 27999
rect 17141 27897 17175 27931
rect 24593 27897 24627 27931
rect 14565 27829 14599 27863
rect 15025 27829 15059 27863
rect 18245 27829 18279 27863
rect 19073 27829 19107 27863
rect 20177 27829 20211 27863
rect 9584 27625 9618 27659
rect 11069 27625 11103 27659
rect 13001 27557 13035 27591
rect 16957 27557 16991 27591
rect 18889 27557 18923 27591
rect 20453 27557 20487 27591
rect 2789 27489 2823 27523
rect 3249 27489 3283 27523
rect 3985 27489 4019 27523
rect 11713 27489 11747 27523
rect 11897 27489 11931 27523
rect 13553 27489 13587 27523
rect 15209 27489 15243 27523
rect 17969 27489 18003 27523
rect 18061 27489 18095 27523
rect 19625 27489 19659 27523
rect 21649 27489 21683 27523
rect 23121 27489 23155 27523
rect 3433 27421 3467 27455
rect 7481 27421 7515 27455
rect 9321 27421 9355 27455
rect 13369 27421 13403 27455
rect 18705 27421 18739 27455
rect 19809 27421 19843 27455
rect 21097 27421 21131 27455
rect 23397 27421 23431 27455
rect 24593 27421 24627 27455
rect 4169 27353 4203 27387
rect 5825 27353 5859 27387
rect 14289 27353 14323 27387
rect 15485 27353 15519 27387
rect 6837 27285 6871 27319
rect 11989 27285 12023 27319
rect 12357 27285 12391 27319
rect 13461 27285 13495 27319
rect 14197 27285 14231 27319
rect 14657 27285 14691 27319
rect 17509 27285 17543 27319
rect 17877 27285 17911 27319
rect 19717 27285 19751 27319
rect 20177 27285 20211 27319
rect 20913 27285 20947 27319
rect 23857 27285 23891 27319
rect 25237 27285 25271 27319
rect 3479 27081 3513 27115
rect 6561 27081 6595 27115
rect 10057 27081 10091 27115
rect 15761 27081 15795 27115
rect 18337 27081 18371 27115
rect 21373 27081 21407 27115
rect 23857 27081 23891 27115
rect 8033 27013 8067 27047
rect 11069 27013 11103 27047
rect 15669 27013 15703 27047
rect 24317 27013 24351 27047
rect 3376 26945 3410 26979
rect 4537 26945 4571 26979
rect 8309 26945 8343 26979
rect 9597 26945 9631 26979
rect 9689 26945 9723 26979
rect 10517 26945 10551 26979
rect 16313 26945 16347 26979
rect 17233 26945 17267 26979
rect 18429 26945 18463 26979
rect 20453 26945 20487 26979
rect 20545 26945 20579 26979
rect 21649 26945 21683 26979
rect 22293 26945 22327 26979
rect 22385 26945 22419 26979
rect 23213 26945 23247 26979
rect 24961 26945 24995 26979
rect 4077 26877 4111 26911
rect 9505 26877 9539 26911
rect 11161 26877 11195 26911
rect 11713 26877 11747 26911
rect 13093 26877 13127 26911
rect 13369 26877 13403 26911
rect 15945 26877 15979 26911
rect 17325 26877 17359 26911
rect 17417 26877 17451 26911
rect 18153 26877 18187 26911
rect 19533 26877 19567 26911
rect 20269 26877 20303 26911
rect 22109 26877 22143 26911
rect 25237 26877 25271 26911
rect 20913 26809 20947 26843
rect 4445 26741 4479 26775
rect 9045 26741 9079 26775
rect 14841 26741 14875 26775
rect 15301 26741 15335 26775
rect 16865 26741 16899 26775
rect 18797 26741 18831 26775
rect 21189 26741 21223 26775
rect 22753 26741 22787 26775
rect 3801 26537 3835 26571
rect 8585 26537 8619 26571
rect 16221 26537 16255 26571
rect 16773 26537 16807 26571
rect 20361 26537 20395 26571
rect 11621 26469 11655 26503
rect 14381 26469 14415 26503
rect 7113 26401 7147 26435
rect 11069 26401 11103 26435
rect 11161 26401 11195 26435
rect 13185 26401 13219 26435
rect 13277 26401 13311 26435
rect 14933 26401 14967 26435
rect 16865 26401 16899 26435
rect 17785 26401 17819 26435
rect 23029 26401 23063 26435
rect 23121 26401 23155 26435
rect 4905 26333 4939 26367
rect 6837 26333 6871 26367
rect 11253 26333 11287 26367
rect 15577 26333 15611 26367
rect 19993 26333 20027 26367
rect 22109 26333 22143 26367
rect 22937 26333 22971 26367
rect 23949 26333 23983 26367
rect 24777 26333 24811 26367
rect 10149 26265 10183 26299
rect 10333 26265 10367 26299
rect 14841 26265 14875 26299
rect 17049 26265 17083 26299
rect 21833 26265 21867 26299
rect 23765 26265 23799 26299
rect 24593 26265 24627 26299
rect 5549 26197 5583 26231
rect 13369 26197 13403 26231
rect 13737 26197 13771 26231
rect 14749 26197 14783 26231
rect 16589 26197 16623 26231
rect 17877 26197 17911 26231
rect 22569 26197 22603 26231
rect 3295 25993 3329 26027
rect 13001 25993 13035 26027
rect 14565 25993 14599 26027
rect 16681 25993 16715 26027
rect 18337 25993 18371 26027
rect 19625 25993 19659 26027
rect 21925 25993 21959 26027
rect 5273 25925 5307 25959
rect 12909 25925 12943 25959
rect 18245 25925 18279 25959
rect 20453 25925 20487 25959
rect 22477 25925 22511 25959
rect 24501 25925 24535 25959
rect 3224 25857 3258 25891
rect 5549 25857 5583 25891
rect 8217 25857 8251 25891
rect 11069 25857 11103 25891
rect 16313 25857 16347 25891
rect 19533 25857 19567 25891
rect 21465 25857 21499 25891
rect 7757 25789 7791 25823
rect 8493 25789 8527 25823
rect 9965 25789 9999 25823
rect 12173 25789 12207 25823
rect 12725 25789 12759 25823
rect 16037 25789 16071 25823
rect 18521 25789 18555 25823
rect 19349 25789 19383 25823
rect 23029 25789 23063 25823
rect 24777 25789 24811 25823
rect 10425 25721 10459 25755
rect 21281 25721 21315 25755
rect 3801 25653 3835 25687
rect 5825 25653 5859 25687
rect 13369 25653 13403 25687
rect 17877 25653 17911 25687
rect 19993 25653 20027 25687
rect 22385 25653 22419 25687
rect 3341 25449 3375 25483
rect 4445 25449 4479 25483
rect 11805 25449 11839 25483
rect 12909 25449 12943 25483
rect 15761 25449 15795 25483
rect 9873 25381 9907 25415
rect 18245 25381 18279 25415
rect 6193 25313 6227 25347
rect 7941 25313 7975 25347
rect 9229 25313 9263 25347
rect 10701 25313 10735 25347
rect 10885 25313 10919 25347
rect 12357 25313 12391 25347
rect 14565 25313 14599 25347
rect 17325 25313 17359 25347
rect 17509 25313 17543 25347
rect 20085 25313 20119 25347
rect 20821 25313 20855 25347
rect 22661 25313 22695 25347
rect 22845 25313 22879 25347
rect 2605 25245 2639 25279
rect 3433 25245 3467 25279
rect 7297 25245 7331 25279
rect 8217 25245 8251 25279
rect 9413 25245 9447 25279
rect 12541 25245 12575 25279
rect 14841 25245 14875 25279
rect 16405 25245 16439 25279
rect 18061 25245 18095 25279
rect 19901 25245 19935 25279
rect 22569 25245 22603 25279
rect 23857 25245 23891 25279
rect 24869 25245 24903 25279
rect 5917 25177 5951 25211
rect 6653 25177 6687 25211
rect 8125 25177 8159 25211
rect 10977 25177 11011 25211
rect 14749 25177 14783 25211
rect 17233 25177 17267 25211
rect 19809 25177 19843 25211
rect 20913 25177 20947 25211
rect 2973 25109 3007 25143
rect 8585 25109 8619 25143
rect 9505 25109 9539 25143
rect 10241 25109 10275 25143
rect 11345 25109 11379 25143
rect 12449 25109 12483 25143
rect 15209 25109 15243 25143
rect 16865 25109 16899 25143
rect 19441 25109 19475 25143
rect 21005 25109 21039 25143
rect 21373 25109 21407 25143
rect 22201 25109 22235 25143
rect 23949 25109 23983 25143
rect 24685 25109 24719 25143
rect 7665 24905 7699 24939
rect 8953 24905 8987 24939
rect 16773 24905 16807 24939
rect 19901 24905 19935 24939
rect 21097 24905 21131 24939
rect 9689 24837 9723 24871
rect 4353 24769 4387 24803
rect 9413 24769 9447 24803
rect 12357 24769 12391 24803
rect 13185 24769 13219 24803
rect 15853 24769 15887 24803
rect 15945 24769 15979 24803
rect 19993 24769 20027 24803
rect 21005 24769 21039 24803
rect 23397 24769 23431 24803
rect 23949 24769 23983 24803
rect 2881 24701 2915 24735
rect 3525 24701 3559 24735
rect 3709 24701 3743 24735
rect 15761 24701 15795 24735
rect 17233 24701 17267 24735
rect 18705 24701 18739 24735
rect 18981 24701 19015 24735
rect 20177 24701 20211 24735
rect 20913 24701 20947 24735
rect 22937 24701 22971 24735
rect 24685 24701 24719 24735
rect 19533 24633 19567 24667
rect 4169 24565 4203 24599
rect 6377 24565 6411 24599
rect 11161 24565 11195 24599
rect 11713 24565 11747 24599
rect 12909 24565 12943 24599
rect 13645 24565 13679 24599
rect 16313 24565 16347 24599
rect 21465 24565 21499 24599
rect 5365 24361 5399 24395
rect 10885 24361 10919 24395
rect 21649 24293 21683 24327
rect 7113 24225 7147 24259
rect 10241 24225 10275 24259
rect 10333 24225 10367 24259
rect 17141 24225 17175 24259
rect 20177 24225 20211 24259
rect 2237 24157 2271 24191
rect 4261 24157 4295 24191
rect 8217 24157 8251 24191
rect 11437 24157 11471 24191
rect 18245 24157 18279 24191
rect 19901 24157 19935 24191
rect 24041 24157 24075 24191
rect 6837 24089 6871 24123
rect 7573 24089 7607 24123
rect 11713 24089 11747 24123
rect 16865 24089 16899 24123
rect 17601 24089 17635 24123
rect 22845 24089 22879 24123
rect 24961 24089 24995 24123
rect 25329 24089 25363 24123
rect 2053 24021 2087 24055
rect 4905 24021 4939 24055
rect 9781 24021 9815 24055
rect 10149 24021 10183 24055
rect 13185 24021 13219 24055
rect 15393 24021 15427 24055
rect 24685 24021 24719 24055
rect 4215 23817 4249 23851
rect 9413 23817 9447 23851
rect 9965 23817 9999 23851
rect 10701 23817 10735 23851
rect 12173 23817 12207 23851
rect 16313 23817 16347 23851
rect 17233 23817 17267 23851
rect 17325 23817 17359 23851
rect 21465 23817 21499 23851
rect 22385 23817 22419 23851
rect 15945 23749 15979 23783
rect 18061 23749 18095 23783
rect 22293 23749 22327 23783
rect 23213 23749 23247 23783
rect 4112 23681 4146 23715
rect 10793 23681 10827 23715
rect 12081 23681 12115 23715
rect 13829 23681 13863 23715
rect 15301 23681 15335 23715
rect 19349 23681 19383 23715
rect 10609 23613 10643 23647
rect 11897 23613 11931 23647
rect 15761 23613 15795 23647
rect 15853 23613 15887 23647
rect 17417 23613 17451 23647
rect 19625 23613 19659 23647
rect 21097 23613 21131 23647
rect 22937 23613 22971 23647
rect 24685 23613 24719 23647
rect 11161 23545 11195 23579
rect 12541 23545 12575 23579
rect 7297 23477 7331 23511
rect 13185 23477 13219 23511
rect 16865 23477 16899 23511
rect 4445 23273 4479 23307
rect 15393 23273 15427 23307
rect 20085 23273 20119 23307
rect 13185 23205 13219 23239
rect 15025 23205 15059 23239
rect 2789 23137 2823 23171
rect 3249 23137 3283 23171
rect 6101 23137 6135 23171
rect 6653 23137 6687 23171
rect 8125 23137 8159 23171
rect 8401 23137 8435 23171
rect 10241 23137 10275 23171
rect 11437 23137 11471 23171
rect 12633 23137 12667 23171
rect 14381 23137 14415 23171
rect 14565 23137 14599 23171
rect 21649 23137 21683 23171
rect 21741 23137 21775 23171
rect 3433 23069 3467 23103
rect 14657 23069 14691 23103
rect 19441 23069 19475 23103
rect 23121 23069 23155 23103
rect 24041 23069 24075 23103
rect 24593 23069 24627 23103
rect 5917 23001 5951 23035
rect 9965 23001 9999 23035
rect 10793 23001 10827 23035
rect 12541 23001 12575 23035
rect 21005 23001 21039 23035
rect 21833 23001 21867 23035
rect 5457 22933 5491 22967
rect 5825 22933 5859 22967
rect 8677 22933 8711 22967
rect 9597 22933 9631 22967
rect 10057 22933 10091 22967
rect 12081 22933 12115 22967
rect 12449 22933 12483 22967
rect 16773 22933 16807 22967
rect 20361 22933 20395 22967
rect 22201 22933 22235 22967
rect 25237 22933 25271 22967
rect 4629 22729 4663 22763
rect 7297 22729 7331 22763
rect 7665 22729 7699 22763
rect 10517 22729 10551 22763
rect 19441 22729 19475 22763
rect 8585 22661 8619 22695
rect 13093 22661 13127 22695
rect 15301 22661 15335 22695
rect 19993 22661 20027 22695
rect 20821 22661 20855 22695
rect 24409 22661 24443 22695
rect 3893 22593 3927 22627
rect 5089 22593 5123 22627
rect 7757 22593 7791 22627
rect 9413 22593 9447 22627
rect 15393 22593 15427 22627
rect 16865 22593 16899 22627
rect 17693 22593 17727 22627
rect 22109 22593 22143 22627
rect 7849 22525 7883 22559
rect 12817 22525 12851 22559
rect 15209 22525 15243 22559
rect 17969 22525 18003 22559
rect 23857 22525 23891 22559
rect 24133 22525 24167 22559
rect 9781 22457 9815 22491
rect 4077 22389 4111 22423
rect 4997 22389 5031 22423
rect 11897 22389 11931 22423
rect 12541 22389 12575 22423
rect 14565 22389 14599 22423
rect 15761 22389 15795 22423
rect 17049 22389 17083 22423
rect 4616 22185 4650 22219
rect 19349 22185 19383 22219
rect 24593 22185 24627 22219
rect 14289 22117 14323 22151
rect 15301 22117 15335 22151
rect 15853 22117 15887 22151
rect 4353 22049 4387 22083
rect 7113 22049 7147 22083
rect 11529 22049 11563 22083
rect 13461 22049 13495 22083
rect 14841 22049 14875 22083
rect 16589 22049 16623 22083
rect 18061 22049 18095 22083
rect 18245 22049 18279 22083
rect 20729 22049 20763 22083
rect 21281 22049 21315 22083
rect 14749 21981 14783 22015
rect 15669 21981 15703 22015
rect 16773 21981 16807 22015
rect 19901 21981 19935 22015
rect 25237 21981 25271 22015
rect 10793 21913 10827 21947
rect 13277 21913 13311 21947
rect 15577 21913 15611 21947
rect 17969 21913 18003 21947
rect 21557 21913 21591 21947
rect 23673 21913 23707 21947
rect 23857 21913 23891 21947
rect 6101 21845 6135 21879
rect 6561 21845 6595 21879
rect 6929 21845 6963 21879
rect 7021 21845 7055 21879
rect 12449 21845 12483 21879
rect 12909 21845 12943 21879
rect 13369 21845 13403 21879
rect 14657 21845 14691 21879
rect 16681 21845 16715 21879
rect 17141 21845 17175 21879
rect 17601 21845 17635 21879
rect 19533 21845 19567 21879
rect 23029 21845 23063 21879
rect 24133 21845 24167 21879
rect 6377 21641 6411 21675
rect 7481 21641 7515 21675
rect 8677 21641 8711 21675
rect 9045 21641 9079 21675
rect 15853 21641 15887 21675
rect 18337 21641 18371 21675
rect 21465 21641 21499 21675
rect 22385 21641 22419 21675
rect 22477 21641 22511 21675
rect 25237 21641 25271 21675
rect 12173 21573 12207 21607
rect 13093 21573 13127 21607
rect 15945 21573 15979 21607
rect 23489 21573 23523 21607
rect 1961 21505 1995 21539
rect 4261 21505 4295 21539
rect 7849 21505 7883 21539
rect 7941 21505 7975 21539
rect 10793 21505 10827 21539
rect 13001 21505 13035 21539
rect 14657 21505 14691 21539
rect 17417 21505 17451 21539
rect 20085 21505 20119 21539
rect 20545 21505 20579 21539
rect 23213 21505 23247 21539
rect 2881 21437 2915 21471
rect 4077 21437 4111 21471
rect 8125 21437 8159 21471
rect 9137 21437 9171 21471
rect 9229 21437 9263 21471
rect 10885 21437 10919 21471
rect 10977 21437 11011 21471
rect 12909 21437 12943 21471
rect 14749 21437 14783 21471
rect 14841 21437 14875 21471
rect 15761 21437 15795 21471
rect 16773 21437 16807 21471
rect 17969 21437 18003 21471
rect 19809 21437 19843 21471
rect 21189 21437 21223 21471
rect 22569 21437 22603 21471
rect 16313 21369 16347 21403
rect 1777 21301 1811 21335
rect 10149 21301 10183 21335
rect 10425 21301 10459 21335
rect 11621 21301 11655 21335
rect 11805 21301 11839 21335
rect 12449 21301 12483 21335
rect 13461 21301 13495 21335
rect 13829 21301 13863 21335
rect 14013 21301 14047 21335
rect 14289 21301 14323 21335
rect 16865 21301 16899 21335
rect 17601 21301 17635 21335
rect 22017 21301 22051 21335
rect 24961 21301 24995 21335
rect 7113 21097 7147 21131
rect 8493 21097 8527 21131
rect 8953 21097 8987 21131
rect 16037 21097 16071 21131
rect 18889 21097 18923 21131
rect 22109 21097 22143 21131
rect 18429 21029 18463 21063
rect 2053 20961 2087 20995
rect 5365 20961 5399 20995
rect 9413 20961 9447 20995
rect 9689 20961 9723 20995
rect 14289 20961 14323 20995
rect 17877 20961 17911 20995
rect 17969 20961 18003 20995
rect 18797 20961 18831 20995
rect 21833 20961 21867 20995
rect 23397 20961 23431 20995
rect 1777 20893 1811 20927
rect 7573 20893 7607 20927
rect 11529 20893 11563 20927
rect 13001 20893 13035 20927
rect 16497 20893 16531 20927
rect 24041 20893 24075 20927
rect 5641 20825 5675 20859
rect 14565 20825 14599 20859
rect 18061 20825 18095 20859
rect 19441 20825 19475 20859
rect 21557 20825 21591 20859
rect 8217 20757 8251 20791
rect 8769 20757 8803 20791
rect 11161 20757 11195 20791
rect 11713 20757 11747 20791
rect 12817 20757 12851 20791
rect 17141 20757 17175 20791
rect 20085 20757 20119 20791
rect 3709 20553 3743 20587
rect 4353 20553 4387 20587
rect 8861 20553 8895 20587
rect 10425 20553 10459 20587
rect 10793 20553 10827 20587
rect 12173 20553 12207 20587
rect 15117 20553 15151 20587
rect 19533 20553 19567 20587
rect 21465 20553 21499 20587
rect 18429 20485 18463 20519
rect 19441 20485 19475 20519
rect 3893 20417 3927 20451
rect 4537 20417 4571 20451
rect 8309 20417 8343 20451
rect 9229 20417 9263 20451
rect 12081 20417 12115 20451
rect 16037 20417 16071 20451
rect 17049 20417 17083 20451
rect 17693 20417 17727 20451
rect 20821 20417 20855 20451
rect 22293 20417 22327 20451
rect 23305 20417 23339 20451
rect 25145 20417 25179 20451
rect 8033 20349 8067 20383
rect 9321 20349 9355 20383
rect 9505 20349 9539 20383
rect 10885 20349 10919 20383
rect 10977 20349 11011 20383
rect 12265 20349 12299 20383
rect 14473 20349 14507 20383
rect 15209 20349 15243 20383
rect 15301 20349 15335 20383
rect 19349 20349 19383 20383
rect 24777 20349 24811 20383
rect 12817 20281 12851 20315
rect 16221 20281 16255 20315
rect 18613 20281 18647 20315
rect 6561 20213 6595 20247
rect 9965 20213 9999 20247
rect 11713 20213 11747 20247
rect 14749 20213 14783 20247
rect 16865 20213 16899 20247
rect 17785 20213 17819 20247
rect 19901 20213 19935 20247
rect 6101 20009 6135 20043
rect 7849 20009 7883 20043
rect 10057 20009 10091 20043
rect 14289 20009 14323 20043
rect 16957 20009 16991 20043
rect 24409 20009 24443 20043
rect 16405 19941 16439 19975
rect 18061 19941 18095 19975
rect 8401 19873 8435 19907
rect 10609 19873 10643 19907
rect 11897 19873 11931 19907
rect 16037 19873 16071 19907
rect 23397 19873 23431 19907
rect 6745 19805 6779 19839
rect 10425 19805 10459 19839
rect 11713 19805 11747 19839
rect 16773 19805 16807 19839
rect 18245 19805 18279 19839
rect 18889 19805 18923 19839
rect 22017 19805 22051 19839
rect 23857 19805 23891 19839
rect 24593 19805 24627 19839
rect 8217 19737 8251 19771
rect 15761 19737 15795 19771
rect 20913 19737 20947 19771
rect 22201 19737 22235 19771
rect 8309 19669 8343 19703
rect 9597 19669 9631 19703
rect 10517 19669 10551 19703
rect 11345 19669 11379 19703
rect 11805 19669 11839 19703
rect 12633 19669 12667 19703
rect 13461 19669 13495 19703
rect 18705 19669 18739 19703
rect 21005 19669 21039 19703
rect 6653 19465 6687 19499
rect 10057 19465 10091 19499
rect 10517 19465 10551 19499
rect 13553 19465 13587 19499
rect 13921 19465 13955 19499
rect 18429 19465 18463 19499
rect 19165 19465 19199 19499
rect 2237 19397 2271 19431
rect 9597 19397 9631 19431
rect 12173 19397 12207 19431
rect 14013 19397 14047 19431
rect 15577 19397 15611 19431
rect 16129 19397 16163 19431
rect 21189 19397 21223 19431
rect 24961 19397 24995 19431
rect 7113 19329 7147 19363
rect 7573 19329 7607 19363
rect 10425 19329 10459 19363
rect 12081 19329 12115 19363
rect 12909 19329 12943 19363
rect 14841 19329 14875 19363
rect 18245 19329 18279 19363
rect 24225 19329 24259 19363
rect 6101 19261 6135 19295
rect 7849 19261 7883 19295
rect 10609 19261 10643 19295
rect 11069 19261 11103 19295
rect 11253 19261 11287 19295
rect 12357 19261 12391 19295
rect 14197 19261 14231 19295
rect 16313 19261 16347 19295
rect 20637 19261 20671 19295
rect 20913 19261 20947 19295
rect 22017 19261 22051 19295
rect 22293 19261 22327 19295
rect 2053 19193 2087 19227
rect 7021 19125 7055 19159
rect 11713 19125 11747 19159
rect 23765 19125 23799 19159
rect 6009 18921 6043 18955
rect 9137 18921 9171 18955
rect 10241 18921 10275 18955
rect 11437 18921 11471 18955
rect 15301 18921 15335 18955
rect 16681 18921 16715 18955
rect 21741 18921 21775 18955
rect 22293 18921 22327 18955
rect 12633 18853 12667 18887
rect 17785 18853 17819 18887
rect 21557 18853 21591 18887
rect 2053 18785 2087 18819
rect 6653 18785 6687 18819
rect 10793 18785 10827 18819
rect 11989 18785 12023 18819
rect 13185 18785 13219 18819
rect 17141 18785 17175 18819
rect 17325 18785 17359 18819
rect 18061 18785 18095 18819
rect 19625 18785 19659 18819
rect 24041 18785 24075 18819
rect 1685 18717 1719 18751
rect 6469 18717 6503 18751
rect 7941 18717 7975 18751
rect 9781 18717 9815 18751
rect 10609 18717 10643 18751
rect 13093 18717 13127 18751
rect 14933 18717 14967 18751
rect 16037 18717 16071 18751
rect 17417 18717 17451 18751
rect 18337 18717 18371 18751
rect 18705 18717 18739 18751
rect 20637 18717 20671 18751
rect 24593 18717 24627 18751
rect 6377 18649 6411 18683
rect 11805 18649 11839 18683
rect 14289 18649 14323 18683
rect 18889 18649 18923 18683
rect 23765 18649 23799 18683
rect 25237 18649 25271 18683
rect 7205 18581 7239 18615
rect 8585 18581 8619 18615
rect 10701 18581 10735 18615
rect 11897 18581 11931 18615
rect 13001 18581 13035 18615
rect 15945 18581 15979 18615
rect 19717 18581 19751 18615
rect 19809 18581 19843 18615
rect 20177 18581 20211 18615
rect 21281 18581 21315 18615
rect 9137 18377 9171 18411
rect 11161 18377 11195 18411
rect 13461 18377 13495 18411
rect 14473 18377 14507 18411
rect 14749 18377 14783 18411
rect 20085 18377 20119 18411
rect 22385 18377 22419 18411
rect 12173 18309 12207 18343
rect 20453 18309 20487 18343
rect 25145 18309 25179 18343
rect 12081 18241 12115 18275
rect 13829 18241 13863 18275
rect 18061 18241 18095 18275
rect 22293 18241 22327 18275
rect 23305 18241 23339 18275
rect 23949 18241 23983 18275
rect 6561 18173 6595 18207
rect 6837 18173 6871 18207
rect 8585 18173 8619 18207
rect 10609 18173 10643 18207
rect 10885 18173 10919 18207
rect 12265 18173 12299 18207
rect 13185 18173 13219 18207
rect 13921 18173 13955 18207
rect 14105 18173 14139 18207
rect 18337 18173 18371 18207
rect 21189 18173 21223 18207
rect 22201 18173 22235 18207
rect 23489 18105 23523 18139
rect 11713 18037 11747 18071
rect 19809 18037 19843 18071
rect 22753 18037 22787 18071
rect 6837 17833 6871 17867
rect 7297 17833 7331 17867
rect 13001 17833 13035 17867
rect 17509 17833 17543 17867
rect 23581 17833 23615 17867
rect 10517 17765 10551 17799
rect 14289 17765 14323 17799
rect 24133 17765 24167 17799
rect 5089 17697 5123 17731
rect 7757 17697 7791 17731
rect 7849 17697 7883 17731
rect 13553 17697 13587 17731
rect 14749 17697 14783 17731
rect 14841 17697 14875 17731
rect 21373 17697 21407 17731
rect 21833 17697 21867 17731
rect 9229 17629 9263 17663
rect 11805 17629 11839 17663
rect 12081 17629 12115 17663
rect 15485 17629 15519 17663
rect 16865 17629 16899 17663
rect 18153 17629 18187 17663
rect 18889 17629 18923 17663
rect 19257 17629 19291 17663
rect 24593 17629 24627 17663
rect 5365 17561 5399 17595
rect 8769 17561 8803 17595
rect 10057 17561 10091 17595
rect 11069 17561 11103 17595
rect 12725 17561 12759 17595
rect 13461 17561 13495 17595
rect 16313 17561 16347 17595
rect 21097 17561 21131 17595
rect 22109 17561 22143 17595
rect 7665 17493 7699 17527
rect 8401 17493 8435 17527
rect 8585 17493 8619 17527
rect 10333 17493 10367 17527
rect 13369 17493 13403 17527
rect 14657 17493 14691 17527
rect 15669 17493 15703 17527
rect 16221 17493 16255 17527
rect 19625 17493 19659 17527
rect 25237 17493 25271 17527
rect 5365 17289 5399 17323
rect 7481 17289 7515 17323
rect 9137 17289 9171 17323
rect 9505 17289 9539 17323
rect 12265 17289 12299 17323
rect 12817 17289 12851 17323
rect 13185 17289 13219 17323
rect 14013 17289 14047 17323
rect 16865 17289 16899 17323
rect 21465 17289 21499 17323
rect 22661 17289 22695 17323
rect 2421 17221 2455 17255
rect 8309 17221 8343 17255
rect 13277 17221 13311 17255
rect 14381 17221 14415 17255
rect 15117 17221 15151 17255
rect 18337 17221 18371 17255
rect 25145 17221 25179 17255
rect 6009 17153 6043 17187
rect 6837 17153 6871 17187
rect 9597 17153 9631 17187
rect 10793 17153 10827 17187
rect 12541 17153 12575 17187
rect 15209 17153 15243 17187
rect 15945 17153 15979 17187
rect 20177 17153 20211 17187
rect 20821 17153 20855 17187
rect 22017 17153 22051 17187
rect 23213 17153 23247 17187
rect 23949 17153 23983 17187
rect 8401 17085 8435 17119
rect 8585 17085 8619 17119
rect 9689 17085 9723 17119
rect 10885 17085 10919 17119
rect 10977 17085 11011 17119
rect 13461 17085 13495 17119
rect 14473 17085 14507 17119
rect 14565 17085 14599 17119
rect 15669 17085 15703 17119
rect 15853 17085 15887 17119
rect 18613 17085 18647 17119
rect 10425 17017 10459 17051
rect 11621 17017 11655 17051
rect 20361 17017 20395 17051
rect 23397 17017 23431 17051
rect 2329 16949 2363 16983
rect 6561 16949 6595 16983
rect 7941 16949 7975 16983
rect 11713 16949 11747 16983
rect 16313 16949 16347 16983
rect 6193 16745 6227 16779
rect 8309 16745 8343 16779
rect 16405 16745 16439 16779
rect 18705 16745 18739 16779
rect 8677 16677 8711 16711
rect 7941 16609 7975 16643
rect 9321 16609 9355 16643
rect 10793 16609 10827 16643
rect 10885 16609 10919 16643
rect 13001 16609 13035 16643
rect 13829 16609 13863 16643
rect 21281 16609 21315 16643
rect 23213 16609 23247 16643
rect 23489 16609 23523 16643
rect 1777 16541 1811 16575
rect 9413 16541 9447 16575
rect 9505 16541 9539 16575
rect 13277 16541 13311 16575
rect 18061 16541 18095 16575
rect 21097 16541 21131 16575
rect 2513 16473 2547 16507
rect 7665 16473 7699 16507
rect 10701 16473 10735 16507
rect 9873 16405 9907 16439
rect 10333 16405 10367 16439
rect 11529 16405 11563 16439
rect 19349 16405 19383 16439
rect 20085 16405 20119 16439
rect 21741 16405 21775 16439
rect 7389 16201 7423 16235
rect 7757 16201 7791 16235
rect 7849 16201 7883 16235
rect 10333 16201 10367 16235
rect 10701 16201 10735 16235
rect 19901 16201 19935 16235
rect 19993 16201 20027 16235
rect 22293 16201 22327 16235
rect 9321 16133 9355 16167
rect 15669 16133 15703 16167
rect 9229 16065 9263 16099
rect 10057 16065 10091 16099
rect 12357 16065 12391 16099
rect 20821 16065 20855 16099
rect 22385 16065 22419 16099
rect 23213 16065 23247 16099
rect 24133 16065 24167 16099
rect 8033 15997 8067 16031
rect 9413 15997 9447 16031
rect 10793 15997 10827 16031
rect 10885 15997 10919 16031
rect 18153 15997 18187 16031
rect 19165 15997 19199 16031
rect 19809 15997 19843 16031
rect 22201 15997 22235 16031
rect 24777 15997 24811 16031
rect 8861 15929 8895 15963
rect 20361 15929 20395 15963
rect 11713 15861 11747 15895
rect 18705 15861 18739 15895
rect 21465 15861 21499 15895
rect 22753 15861 22787 15895
rect 7941 15657 7975 15691
rect 9597 15657 9631 15691
rect 13203 15657 13237 15691
rect 17693 15657 17727 15691
rect 20177 15657 20211 15691
rect 10241 15521 10275 15555
rect 13461 15521 13495 15555
rect 15393 15521 15427 15555
rect 15945 15521 15979 15555
rect 18245 15521 18279 15555
rect 19625 15521 19659 15555
rect 20821 15521 20855 15555
rect 20913 15521 20947 15555
rect 22293 15521 22327 15555
rect 7481 15453 7515 15487
rect 8585 15453 8619 15487
rect 10057 15453 10091 15487
rect 15209 15453 15243 15487
rect 18521 15453 18555 15487
rect 19809 15453 19843 15487
rect 22017 15453 22051 15487
rect 22753 15453 22787 15487
rect 14289 15385 14323 15419
rect 15117 15385 15151 15419
rect 16221 15385 16255 15419
rect 19717 15385 19751 15419
rect 23857 15385 23891 15419
rect 6837 15317 6871 15351
rect 9229 15317 9263 15351
rect 9965 15317 9999 15351
rect 11253 15317 11287 15351
rect 11713 15317 11747 15351
rect 13737 15317 13771 15351
rect 14473 15317 14507 15351
rect 14749 15317 14783 15351
rect 18429 15317 18463 15351
rect 18889 15317 18923 15351
rect 21005 15317 21039 15351
rect 21373 15317 21407 15351
rect 21833 15317 21867 15351
rect 8769 15113 8803 15147
rect 13645 15113 13679 15147
rect 14105 15113 14139 15147
rect 16313 15113 16347 15147
rect 17509 15113 17543 15147
rect 18153 15113 18187 15147
rect 20821 15113 20855 15147
rect 7021 15045 7055 15079
rect 10885 15045 10919 15079
rect 13369 15045 13403 15079
rect 15025 15045 15059 15079
rect 17049 15045 17083 15079
rect 11713 14977 11747 15011
rect 14013 14977 14047 15011
rect 15669 14977 15703 15011
rect 19073 14977 19107 15011
rect 21465 14977 21499 15011
rect 22753 14977 22787 15011
rect 23949 14977 23983 15011
rect 6745 14909 6779 14943
rect 11161 14909 11195 14943
rect 14197 14909 14231 14943
rect 17969 14909 18003 14943
rect 18061 14909 18095 14943
rect 19349 14909 19383 14943
rect 21833 14909 21867 14943
rect 24685 14909 24719 14943
rect 14841 14841 14875 14875
rect 16865 14841 16899 14875
rect 22937 14841 22971 14875
rect 8493 14773 8527 14807
rect 9413 14773 9447 14807
rect 12357 14773 12391 14807
rect 18521 14773 18555 14807
rect 21281 14773 21315 14807
rect 6837 14569 6871 14603
rect 11989 14569 12023 14603
rect 13001 14569 13035 14603
rect 15577 14569 15611 14603
rect 20453 14569 20487 14603
rect 12725 14501 12759 14535
rect 18981 14501 19015 14535
rect 8585 14433 8619 14467
rect 9873 14433 9907 14467
rect 12541 14433 12575 14467
rect 13461 14433 13495 14467
rect 13553 14433 13587 14467
rect 14565 14433 14599 14467
rect 17325 14433 17359 14467
rect 21373 14433 21407 14467
rect 14749 14365 14783 14399
rect 17785 14365 17819 14399
rect 19625 14365 19659 14399
rect 21097 14365 21131 14399
rect 23397 14365 23431 14399
rect 8309 14297 8343 14331
rect 10149 14297 10183 14331
rect 13369 14297 13403 14331
rect 17049 14297 17083 14331
rect 18429 14297 18463 14331
rect 23581 14297 23615 14331
rect 8953 14229 8987 14263
rect 11621 14229 11655 14263
rect 14657 14229 14691 14263
rect 15117 14229 15151 14263
rect 19441 14229 19475 14263
rect 22845 14229 22879 14263
rect 10241 14025 10275 14059
rect 11805 14025 11839 14059
rect 13001 14025 13035 14059
rect 13369 14025 13403 14059
rect 19441 14025 19475 14059
rect 20545 14025 20579 14059
rect 21005 14025 21039 14059
rect 9965 13957 9999 13991
rect 12265 13957 12299 13991
rect 15761 13957 15795 13991
rect 16221 13957 16255 13991
rect 17877 13957 17911 13991
rect 18337 13957 18371 13991
rect 20637 13957 20671 13991
rect 23305 13957 23339 13991
rect 25145 13957 25179 13991
rect 2789 13889 2823 13923
rect 7941 13889 7975 13923
rect 12173 13889 12207 13923
rect 13461 13889 13495 13923
rect 14381 13889 14415 13923
rect 18797 13889 18831 13923
rect 22845 13889 22879 13923
rect 23949 13889 23983 13923
rect 1777 13821 1811 13855
rect 8217 13821 8251 13855
rect 12357 13821 12391 13855
rect 13553 13821 13587 13855
rect 14197 13821 14231 13855
rect 15301 13821 15335 13855
rect 15945 13821 15979 13855
rect 17141 13821 17175 13855
rect 18061 13821 18095 13855
rect 20453 13821 20487 13855
rect 22201 13821 22235 13855
rect 14749 13685 14783 13719
rect 9781 13481 9815 13515
rect 12265 13481 12299 13515
rect 14197 13481 14231 13515
rect 15209 13481 15243 13515
rect 22293 13481 22327 13515
rect 13369 13413 13403 13447
rect 12725 13345 12759 13379
rect 12909 13345 12943 13379
rect 13645 13345 13679 13379
rect 14381 13345 14415 13379
rect 19257 13345 19291 13379
rect 9137 13277 9171 13311
rect 13001 13277 13035 13311
rect 13921 13277 13955 13311
rect 16957 13277 16991 13311
rect 17417 13277 17451 13311
rect 18613 13277 18647 13311
rect 18797 13277 18831 13311
rect 21833 13277 21867 13311
rect 22661 13277 22695 13311
rect 16681 13209 16715 13243
rect 18061 13209 18095 13243
rect 20177 13209 20211 13243
rect 20361 13209 20395 13243
rect 21097 13209 21131 13243
rect 23857 13209 23891 13243
rect 20637 13141 20671 13175
rect 11253 12937 11287 12971
rect 12173 12937 12207 12971
rect 14013 12937 14047 12971
rect 14381 12937 14415 12971
rect 17233 12937 17267 12971
rect 18153 12937 18187 12971
rect 22293 12937 22327 12971
rect 12633 12869 12667 12903
rect 14473 12869 14507 12903
rect 15577 12869 15611 12903
rect 16037 12869 16071 12903
rect 20177 12869 20211 12903
rect 20729 12869 20763 12903
rect 21373 12869 21407 12903
rect 13369 12801 13403 12835
rect 17141 12801 17175 12835
rect 21005 12801 21039 12835
rect 22385 12801 22419 12835
rect 23213 12801 23247 12835
rect 23949 12801 23983 12835
rect 14657 12733 14691 12767
rect 17049 12733 17083 12767
rect 19625 12733 19659 12767
rect 19901 12733 19935 12767
rect 22109 12733 22143 12767
rect 24777 12733 24811 12767
rect 12817 12665 12851 12699
rect 15761 12665 15795 12699
rect 23397 12665 23431 12699
rect 13461 12597 13495 12631
rect 17601 12597 17635 12631
rect 22753 12597 22787 12631
rect 16037 12393 16071 12427
rect 19901 12325 19935 12359
rect 23397 12325 23431 12359
rect 9413 12257 9447 12291
rect 9689 12257 9723 12291
rect 14289 12257 14323 12291
rect 17969 12257 18003 12291
rect 18061 12257 18095 12291
rect 18797 12257 18831 12291
rect 21649 12257 21683 12291
rect 22293 12257 22327 12291
rect 11621 12189 11655 12223
rect 13737 12189 13771 12223
rect 23213 12189 23247 12223
rect 23857 12189 23891 12223
rect 13093 12121 13127 12155
rect 14565 12121 14599 12155
rect 18153 12121 18187 12155
rect 21373 12121 21407 12155
rect 11161 12053 11195 12087
rect 12265 12053 12299 12087
rect 18521 12053 18555 12087
rect 24041 12053 24075 12087
rect 10701 11849 10735 11883
rect 16865 11849 16899 11883
rect 17233 11849 17267 11883
rect 21005 11849 21039 11883
rect 15301 11781 15335 11815
rect 15853 11781 15887 11815
rect 16313 11781 16347 11815
rect 21281 11781 21315 11815
rect 22109 11781 22143 11815
rect 23213 11781 23247 11815
rect 25145 11781 25179 11815
rect 10793 11713 10827 11747
rect 18153 11713 18187 11747
rect 20361 11713 20395 11747
rect 22753 11713 22787 11747
rect 23949 11713 23983 11747
rect 10609 11645 10643 11679
rect 12173 11645 12207 11679
rect 12449 11645 12483 11679
rect 14473 11645 14507 11679
rect 17325 11645 17359 11679
rect 17417 11645 17451 11679
rect 18429 11645 18463 11679
rect 16037 11577 16071 11611
rect 22293 11577 22327 11611
rect 22937 11577 22971 11611
rect 11161 11509 11195 11543
rect 13921 11509 13955 11543
rect 19901 11509 19935 11543
rect 12909 11305 12943 11339
rect 13921 11305 13955 11339
rect 15209 11305 15243 11339
rect 18981 11305 19015 11339
rect 19441 11305 19475 11339
rect 14841 11237 14875 11271
rect 10701 11169 10735 11203
rect 12449 11169 12483 11203
rect 15761 11169 15795 11203
rect 13553 11101 13587 11135
rect 14473 11101 14507 11135
rect 15577 11101 15611 11135
rect 18429 11101 18463 11135
rect 20085 11101 20119 11135
rect 20637 11101 20671 11135
rect 21373 11101 21407 11135
rect 21833 11101 21867 11135
rect 10977 11033 11011 11067
rect 14289 11033 14323 11067
rect 15669 11033 15703 11067
rect 18613 11033 18647 11067
rect 20821 11033 20855 11067
rect 21557 11033 21591 11067
rect 16405 10965 16439 10999
rect 11529 10761 11563 10795
rect 12633 10761 12667 10795
rect 15669 10761 15703 10795
rect 19533 10761 19567 10795
rect 20637 10761 20671 10795
rect 11989 10693 12023 10727
rect 15301 10693 15335 10727
rect 19625 10693 19659 10727
rect 21097 10693 21131 10727
rect 16129 10625 16163 10659
rect 18613 10625 18647 10659
rect 20453 10625 20487 10659
rect 22017 10625 22051 10659
rect 23305 10625 23339 10659
rect 23949 10625 23983 10659
rect 14565 10557 14599 10591
rect 15117 10557 15151 10591
rect 15209 10557 15243 10591
rect 19441 10557 19475 10591
rect 24777 10557 24811 10591
rect 16313 10489 16347 10523
rect 22201 10489 22235 10523
rect 12081 10421 12115 10455
rect 18797 10421 18831 10455
rect 19993 10421 20027 10455
rect 23489 10421 23523 10455
rect 16865 10013 16899 10047
rect 22017 10013 22051 10047
rect 22845 10013 22879 10047
rect 23857 10013 23891 10047
rect 17049 9945 17083 9979
rect 24777 9945 24811 9979
rect 22201 9877 22235 9911
rect 24685 9877 24719 9911
rect 22845 9673 22879 9707
rect 14565 9605 14599 9639
rect 22661 9537 22695 9571
rect 23305 9537 23339 9571
rect 23949 9537 23983 9571
rect 24777 9469 24811 9503
rect 14657 9333 14691 9367
rect 23489 9333 23523 9367
rect 16589 8925 16623 8959
rect 19533 8925 19567 8959
rect 23765 8925 23799 8959
rect 24869 8925 24903 8959
rect 19717 8857 19751 8891
rect 7849 8789 7883 8823
rect 16681 8789 16715 8823
rect 23949 8789 23983 8823
rect 24685 8789 24719 8823
rect 7757 8585 7791 8619
rect 8125 8585 8159 8619
rect 20913 8517 20947 8551
rect 25145 8517 25179 8551
rect 7665 8449 7699 8483
rect 22109 8449 22143 8483
rect 23949 8449 23983 8483
rect 7573 8381 7607 8415
rect 21557 8381 21591 8415
rect 22661 8381 22695 8415
rect 20729 8313 20763 8347
rect 3985 7905 4019 7939
rect 23305 7905 23339 7939
rect 6285 7837 6319 7871
rect 21557 7837 21591 7871
rect 22661 7837 22695 7871
rect 24869 7837 24903 7871
rect 4261 7769 4295 7803
rect 6009 7769 6043 7803
rect 19533 7769 19567 7803
rect 19717 7769 19751 7803
rect 21741 7701 21775 7735
rect 24685 7701 24719 7735
rect 4629 7497 4663 7531
rect 18429 7429 18463 7463
rect 25145 7429 25179 7463
rect 3985 7361 4019 7395
rect 20637 7361 20671 7395
rect 23305 7361 23339 7395
rect 23949 7361 23983 7395
rect 23029 7293 23063 7327
rect 18521 7157 18555 7191
rect 20453 7157 20487 7191
rect 23397 6817 23431 6851
rect 19625 6749 19659 6783
rect 20821 6749 20855 6783
rect 24041 6749 24075 6783
rect 24777 6749 24811 6783
rect 21925 6681 21959 6715
rect 19809 6613 19843 6647
rect 24593 6613 24627 6647
rect 3709 6409 3743 6443
rect 19533 6409 19567 6443
rect 19441 6341 19475 6375
rect 3065 6273 3099 6307
rect 21465 6273 21499 6307
rect 22109 6273 22143 6307
rect 23949 6273 23983 6307
rect 21005 6205 21039 6239
rect 22569 6205 22603 6239
rect 24777 6205 24811 6239
rect 22477 5729 22511 5763
rect 20361 5661 20395 5695
rect 22017 5661 22051 5695
rect 24777 5661 24811 5695
rect 21373 5593 21407 5627
rect 24593 5593 24627 5627
rect 2513 5321 2547 5355
rect 1777 5185 1811 5219
rect 3157 5185 3191 5219
rect 19257 5185 19291 5219
rect 21005 5185 21039 5219
rect 22017 5185 22051 5219
rect 24133 5185 24167 5219
rect 18889 5117 18923 5151
rect 19993 5117 20027 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 1961 5049 1995 5083
rect 1501 4981 1535 5015
rect 3985 4777 4019 4811
rect 2881 4709 2915 4743
rect 1961 4641 1995 4675
rect 18429 4641 18463 4675
rect 23489 4641 23523 4675
rect 2697 4573 2731 4607
rect 3249 4573 3283 4607
rect 4169 4573 4203 4607
rect 18889 4573 18923 4607
rect 19625 4573 19659 4607
rect 21281 4573 21315 4607
rect 23213 4573 23247 4607
rect 1777 4505 1811 4539
rect 20361 4505 20395 4539
rect 22201 4505 22235 4539
rect 2237 4437 2271 4471
rect 1593 4097 1627 4131
rect 3341 4097 3375 4131
rect 11989 4097 12023 4131
rect 13553 4097 13587 4131
rect 16129 4097 16163 4131
rect 16313 4097 16347 4131
rect 16865 4097 16899 4131
rect 18797 4097 18831 4131
rect 22201 4097 22235 4131
rect 23857 4097 23891 4131
rect 3617 4029 3651 4063
rect 4077 4029 4111 4063
rect 11345 4029 11379 4063
rect 11713 4029 11747 4063
rect 14013 4029 14047 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 3985 3961 4019 3995
rect 9965 3961 9999 3995
rect 2237 3893 2271 3927
rect 4353 3893 4387 3927
rect 6377 3893 6411 3927
rect 9505 3893 9539 3927
rect 9781 3893 9815 3927
rect 11069 3893 11103 3927
rect 6745 3689 6779 3723
rect 8217 3689 8251 3723
rect 9229 3689 9263 3723
rect 10057 3689 10091 3723
rect 4169 3621 4203 3655
rect 5273 3621 5307 3655
rect 6101 3621 6135 3655
rect 7573 3553 7607 3587
rect 11253 3553 11287 3587
rect 17325 3553 17359 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 2421 3485 2455 3519
rect 2881 3485 2915 3519
rect 3157 3485 3191 3519
rect 3985 3485 4019 3519
rect 5089 3485 5123 3519
rect 5917 3485 5951 3519
rect 6561 3485 6595 3519
rect 8033 3485 8067 3519
rect 9413 3485 9447 3519
rect 9873 3485 9907 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 13737 3485 13771 3519
rect 16405 3485 16439 3519
rect 16865 3485 16899 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 4537 3417 4571 3451
rect 12725 3417 12759 3451
rect 15209 3417 15243 3451
rect 1409 3349 1443 3383
rect 1777 3349 1811 3383
rect 3341 3349 3375 3383
rect 4813 3349 4847 3383
rect 7205 3349 7239 3383
rect 7757 3349 7791 3383
rect 8677 3349 8711 3383
rect 10701 3349 10735 3383
rect 3525 3145 3559 3179
rect 5181 3145 5215 3179
rect 5917 3145 5951 3179
rect 7757 3145 7791 3179
rect 8401 3145 8435 3179
rect 11897 3145 11931 3179
rect 4261 3077 4295 3111
rect 21557 3077 21591 3111
rect 22937 3077 22971 3111
rect 1777 3009 1811 3043
rect 2881 3009 2915 3043
rect 4077 3009 4111 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5733 3009 5767 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 8585 3009 8619 3043
rect 9873 3009 9907 3043
rect 11161 3009 11195 3043
rect 11713 3009 11747 3043
rect 13737 3009 13771 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 22017 3009 22051 3043
rect 23857 3009 23891 3043
rect 2421 2941 2455 2975
rect 9597 2941 9631 2975
rect 10885 2941 10919 2975
rect 13369 2941 13403 2975
rect 14749 2941 14783 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 24317 2941 24351 2975
rect 6469 2805 6503 2839
rect 7021 2805 7055 2839
rect 1593 2601 1627 2635
rect 4077 2601 4111 2635
rect 9781 2601 9815 2635
rect 18521 2601 18555 2635
rect 24685 2601 24719 2635
rect 3341 2465 3375 2499
rect 5273 2465 5307 2499
rect 10885 2465 10919 2499
rect 14105 2465 14139 2499
rect 15209 2465 15243 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 2237 2397 2271 2431
rect 2697 2397 2731 2431
rect 4261 2397 4295 2431
rect 5549 2397 5583 2431
rect 5825 2397 5859 2431
rect 6469 2397 6503 2431
rect 6929 2397 6963 2431
rect 7665 2397 7699 2431
rect 7941 2397 7975 2431
rect 9137 2397 9171 2431
rect 9597 2397 9631 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 12357 2397 12391 2431
rect 14657 2397 14691 2431
rect 17049 2397 17083 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 24041 2397 24075 2431
rect 6101 2329 6135 2363
rect 6653 2329 6687 2363
rect 9321 2329 9355 2363
rect 13553 2329 13587 2363
rect 24777 2329 24811 2363
rect 25145 2329 25179 2363
rect 7113 2261 7147 2295
rect 11897 2261 11931 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 14553 54315 14611 54321
rect 14553 54281 14565 54315
rect 14599 54312 14611 54315
rect 14734 54312 14740 54324
rect 14599 54284 14740 54312
rect 14599 54281 14611 54284
rect 14553 54275 14611 54281
rect 14734 54272 14740 54284
rect 14792 54272 14798 54324
rect 16206 54272 16212 54324
rect 16264 54312 16270 54324
rect 16393 54315 16451 54321
rect 16393 54312 16405 54315
rect 16264 54284 16405 54312
rect 16264 54272 16270 54284
rect 16393 54281 16405 54284
rect 16439 54312 16451 54315
rect 16439 54284 16574 54312
rect 16439 54281 16451 54284
rect 16393 54275 16451 54281
rect 10965 54247 11023 54253
rect 8588 54216 10088 54244
rect 3421 54179 3479 54185
rect 3421 54145 3433 54179
rect 3467 54176 3479 54179
rect 5626 54176 5632 54188
rect 3467 54148 5632 54176
rect 3467 54145 3479 54148
rect 3421 54139 3479 54145
rect 5626 54136 5632 54148
rect 5684 54136 5690 54188
rect 5994 54136 6000 54188
rect 6052 54136 6058 54188
rect 7834 54176 7840 54188
rect 6886 54148 7840 54176
rect 2961 54111 3019 54117
rect 2961 54077 2973 54111
rect 3007 54108 3019 54111
rect 3970 54108 3976 54120
rect 3007 54080 3976 54108
rect 3007 54077 3019 54080
rect 2961 54071 3019 54077
rect 3970 54068 3976 54080
rect 4028 54068 4034 54120
rect 5537 54111 5595 54117
rect 5537 54077 5549 54111
rect 5583 54108 5595 54111
rect 6886 54108 6914 54148
rect 7834 54136 7840 54148
rect 7892 54136 7898 54188
rect 8588 54185 8616 54216
rect 8573 54179 8631 54185
rect 8573 54145 8585 54179
rect 8619 54145 8631 54179
rect 8573 54139 8631 54145
rect 9950 54136 9956 54188
rect 10008 54136 10014 54188
rect 10060 54176 10088 54216
rect 10965 54213 10977 54247
rect 11011 54244 11023 54247
rect 11422 54244 11428 54256
rect 11011 54216 11428 54244
rect 11011 54213 11023 54216
rect 10965 54207 11023 54213
rect 11422 54204 11428 54216
rect 11480 54204 11486 54256
rect 12894 54244 12900 54256
rect 11716 54216 12900 54244
rect 11514 54176 11520 54188
rect 10060 54148 11520 54176
rect 11514 54136 11520 54148
rect 11572 54136 11578 54188
rect 11716 54185 11744 54216
rect 12894 54204 12900 54216
rect 12952 54244 12958 54256
rect 14093 54247 14151 54253
rect 14093 54244 14105 54247
rect 12952 54216 14105 54244
rect 12952 54204 12958 54216
rect 14093 54213 14105 54216
rect 14139 54213 14151 54247
rect 14093 54207 14151 54213
rect 11701 54179 11759 54185
rect 11701 54145 11713 54179
rect 11747 54145 11759 54179
rect 11701 54139 11759 54145
rect 12526 54136 12532 54188
rect 12584 54136 12590 54188
rect 14752 54176 14780 54272
rect 14829 54179 14887 54185
rect 14829 54176 14841 54179
rect 14752 54148 14841 54176
rect 14829 54145 14841 54148
rect 14875 54145 14887 54179
rect 14829 54139 14887 54145
rect 15194 54136 15200 54188
rect 15252 54176 15258 54188
rect 15841 54179 15899 54185
rect 15841 54176 15853 54179
rect 15252 54148 15853 54176
rect 15252 54136 15258 54148
rect 15841 54145 15853 54148
rect 15887 54176 15899 54179
rect 16117 54179 16175 54185
rect 16117 54176 16129 54179
rect 15887 54148 16129 54176
rect 15887 54145 15899 54148
rect 15841 54139 15899 54145
rect 16117 54145 16129 54148
rect 16163 54145 16175 54179
rect 16546 54176 16574 54284
rect 24486 54272 24492 54324
rect 24544 54272 24550 54324
rect 24670 54272 24676 54324
rect 24728 54272 24734 54324
rect 18877 54247 18935 54253
rect 18877 54244 18889 54247
rect 17880 54216 18889 54244
rect 16853 54179 16911 54185
rect 16853 54176 16865 54179
rect 16546 54148 16865 54176
rect 16117 54139 16175 54145
rect 16853 54145 16865 54148
rect 16899 54145 16911 54179
rect 16853 54139 16911 54145
rect 16942 54136 16948 54188
rect 17000 54176 17006 54188
rect 17880 54185 17908 54216
rect 18877 54213 18889 54216
rect 18923 54213 18935 54247
rect 18877 54207 18935 54213
rect 19518 54204 19524 54256
rect 19576 54244 19582 54256
rect 21453 54247 21511 54253
rect 21453 54244 21465 54247
rect 19576 54216 21465 54244
rect 19576 54204 19582 54216
rect 17865 54179 17923 54185
rect 17865 54176 17877 54179
rect 17000 54148 17877 54176
rect 17000 54136 17006 54148
rect 17865 54145 17877 54148
rect 17911 54145 17923 54179
rect 17865 54139 17923 54145
rect 17954 54136 17960 54188
rect 18012 54176 18018 54188
rect 18506 54176 18512 54188
rect 18012 54148 18512 54176
rect 18012 54136 18018 54148
rect 18506 54136 18512 54148
rect 18564 54136 18570 54188
rect 18598 54136 18604 54188
rect 18656 54176 18662 54188
rect 19702 54176 19708 54188
rect 18656 54148 19708 54176
rect 18656 54136 18662 54148
rect 19702 54136 19708 54148
rect 19760 54136 19766 54188
rect 20456 54185 20484 54216
rect 21453 54213 21465 54216
rect 21499 54213 21511 54247
rect 23293 54247 23351 54253
rect 23293 54244 23305 54247
rect 21453 54207 21511 54213
rect 22296 54216 23305 54244
rect 20441 54179 20499 54185
rect 20441 54145 20453 54179
rect 20487 54145 20499 54179
rect 20441 54139 20499 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 21174 54176 21180 54188
rect 20772 54148 21180 54176
rect 20772 54136 20778 54148
rect 21174 54136 21180 54148
rect 21232 54136 21238 54188
rect 21358 54136 21364 54188
rect 21416 54176 21422 54188
rect 22296 54185 22324 54216
rect 23293 54213 23305 54216
rect 23339 54213 23351 54247
rect 23293 54207 23351 54213
rect 22281 54179 22339 54185
rect 22281 54176 22293 54179
rect 21416 54148 22293 54176
rect 21416 54136 21422 54148
rect 22281 54145 22293 54148
rect 22327 54145 22339 54179
rect 22281 54139 22339 54145
rect 22462 54136 22468 54188
rect 22520 54176 22526 54188
rect 22741 54179 22799 54185
rect 22741 54176 22753 54179
rect 22520 54148 22753 54176
rect 22520 54136 22526 54148
rect 22741 54145 22753 54148
rect 22787 54145 22799 54179
rect 22741 54139 22799 54145
rect 24029 54179 24087 54185
rect 24029 54145 24041 54179
rect 24075 54176 24087 54179
rect 24688 54176 24716 54272
rect 24075 54148 24716 54176
rect 24075 54145 24087 54148
rect 24029 54139 24087 54145
rect 25314 54136 25320 54188
rect 25372 54136 25378 54188
rect 5583 54080 6914 54108
rect 8113 54111 8171 54117
rect 5583 54077 5595 54080
rect 5537 54071 5595 54077
rect 8113 54077 8125 54111
rect 8159 54108 8171 54111
rect 9858 54108 9864 54120
rect 8159 54080 9864 54108
rect 8159 54077 8171 54080
rect 8113 54071 8171 54077
rect 9858 54068 9864 54080
rect 9916 54068 9922 54120
rect 12618 54068 12624 54120
rect 12676 54108 12682 54120
rect 12805 54111 12863 54117
rect 12805 54108 12817 54111
rect 12676 54080 12817 54108
rect 12676 54068 12682 54080
rect 12805 54077 12817 54080
rect 12851 54077 12863 54111
rect 12805 54071 12863 54077
rect 16758 54000 16764 54052
rect 16816 54040 16822 54052
rect 17681 54043 17739 54049
rect 17681 54040 17693 54043
rect 16816 54012 17693 54040
rect 16816 54000 16822 54012
rect 17681 54009 17693 54012
rect 17727 54009 17739 54043
rect 17681 54003 17739 54009
rect 11885 53975 11943 53981
rect 11885 53941 11897 53975
rect 11931 53972 11943 53975
rect 12710 53972 12716 53984
rect 11931 53944 12716 53972
rect 11931 53941 11943 53944
rect 11885 53935 11943 53941
rect 12710 53932 12716 53944
rect 12768 53932 12774 53984
rect 15010 53932 15016 53984
rect 15068 53932 15074 53984
rect 15657 53975 15715 53981
rect 15657 53941 15669 53975
rect 15703 53972 15715 53975
rect 15746 53972 15752 53984
rect 15703 53944 15752 53972
rect 15703 53941 15715 53944
rect 15657 53935 15715 53941
rect 15746 53932 15752 53944
rect 15804 53932 15810 53984
rect 17034 53932 17040 53984
rect 17092 53932 17098 53984
rect 18414 53932 18420 53984
rect 18472 53932 18478 53984
rect 19334 53932 19340 53984
rect 19392 53972 19398 53984
rect 19521 53975 19579 53981
rect 19521 53972 19533 53975
rect 19392 53944 19533 53972
rect 19392 53932 19398 53944
rect 19521 53941 19533 53944
rect 19567 53941 19579 53975
rect 19521 53935 19579 53941
rect 20257 53975 20315 53981
rect 20257 53941 20269 53975
rect 20303 53972 20315 53975
rect 20438 53972 20444 53984
rect 20303 53944 20444 53972
rect 20303 53941 20315 53944
rect 20257 53935 20315 53941
rect 20438 53932 20444 53944
rect 20496 53932 20502 53984
rect 20993 53975 21051 53981
rect 20993 53941 21005 53975
rect 21039 53972 21051 53975
rect 21634 53972 21640 53984
rect 21039 53944 21640 53972
rect 21039 53941 21051 53944
rect 20993 53935 21051 53941
rect 21634 53932 21640 53944
rect 21692 53932 21698 53984
rect 22097 53975 22155 53981
rect 22097 53941 22109 53975
rect 22143 53972 22155 53975
rect 22186 53972 22192 53984
rect 22143 53944 22192 53972
rect 22143 53941 22155 53944
rect 22097 53935 22155 53941
rect 22186 53932 22192 53944
rect 22244 53932 22250 53984
rect 22278 53932 22284 53984
rect 22336 53972 22342 53984
rect 22925 53975 22983 53981
rect 22925 53972 22937 53975
rect 22336 53944 22937 53972
rect 22336 53932 22342 53944
rect 22925 53941 22937 53944
rect 22971 53941 22983 53975
rect 22925 53935 22983 53941
rect 23845 53975 23903 53981
rect 23845 53941 23857 53975
rect 23891 53972 23903 53975
rect 24578 53972 24584 53984
rect 23891 53944 24584 53972
rect 23891 53941 23903 53944
rect 23845 53935 23903 53941
rect 24578 53932 24584 53944
rect 24636 53932 24642 53984
rect 25133 53975 25191 53981
rect 25133 53941 25145 53975
rect 25179 53972 25191 53975
rect 25958 53972 25964 53984
rect 25179 53944 25964 53972
rect 25179 53941 25191 53944
rect 25133 53935 25191 53941
rect 25958 53932 25964 53944
rect 26016 53932 26022 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 3970 53728 3976 53780
rect 4028 53768 4034 53780
rect 5902 53768 5908 53780
rect 4028 53740 5908 53768
rect 4028 53728 4034 53740
rect 5902 53728 5908 53740
rect 5960 53728 5966 53780
rect 16393 53771 16451 53777
rect 16393 53737 16405 53771
rect 16439 53768 16451 53771
rect 16574 53768 16580 53780
rect 16439 53740 16580 53768
rect 16439 53737 16451 53740
rect 16393 53731 16451 53737
rect 16574 53728 16580 53740
rect 16632 53728 16638 53780
rect 18506 53728 18512 53780
rect 18564 53768 18570 53780
rect 18877 53771 18935 53777
rect 18877 53768 18889 53771
rect 18564 53740 18889 53768
rect 18564 53728 18570 53740
rect 18877 53737 18889 53740
rect 18923 53737 18935 53771
rect 18877 53731 18935 53737
rect 9769 53703 9827 53709
rect 9769 53700 9781 53703
rect 4632 53672 9781 53700
rect 2961 53635 3019 53641
rect 2961 53601 2973 53635
rect 3007 53632 3019 53635
rect 3007 53604 4568 53632
rect 3007 53601 3019 53604
rect 2961 53595 3019 53601
rect 3421 53567 3479 53573
rect 3421 53533 3433 53567
rect 3467 53564 3479 53567
rect 3467 53536 4476 53564
rect 3467 53533 3479 53536
rect 3421 53527 3479 53533
rect 2406 53388 2412 53440
rect 2464 53428 2470 53440
rect 3973 53431 4031 53437
rect 3973 53428 3985 53431
rect 2464 53400 3985 53428
rect 2464 53388 2470 53400
rect 3973 53397 3985 53400
rect 4019 53397 4031 53431
rect 4448 53428 4476 53536
rect 4540 53496 4568 53604
rect 4632 53573 4660 53672
rect 9769 53669 9781 53672
rect 9815 53669 9827 53703
rect 9769 53663 9827 53669
rect 20622 53660 20628 53712
rect 20680 53700 20686 53712
rect 21821 53703 21879 53709
rect 21821 53700 21833 53703
rect 20680 53672 21833 53700
rect 20680 53660 20686 53672
rect 21821 53669 21833 53672
rect 21867 53669 21879 53703
rect 21821 53663 21879 53669
rect 22278 53660 22284 53712
rect 22336 53700 22342 53712
rect 23109 53703 23167 53709
rect 23109 53700 23121 53703
rect 22336 53672 23121 53700
rect 22336 53660 22342 53672
rect 23109 53669 23121 53672
rect 23155 53669 23167 53703
rect 23109 53663 23167 53669
rect 6273 53635 6331 53641
rect 6273 53601 6285 53635
rect 6319 53601 6331 53635
rect 6273 53595 6331 53601
rect 8113 53635 8171 53641
rect 8113 53601 8125 53635
rect 8159 53632 8171 53635
rect 8846 53632 8852 53644
rect 8159 53604 8852 53632
rect 8159 53601 8171 53604
rect 8113 53595 8171 53601
rect 4617 53567 4675 53573
rect 4617 53533 4629 53567
rect 4663 53533 4675 53567
rect 4617 53527 4675 53533
rect 5534 53524 5540 53576
rect 5592 53524 5598 53576
rect 5552 53496 5580 53524
rect 4540 53468 5580 53496
rect 6288 53496 6316 53595
rect 8846 53592 8852 53604
rect 8904 53592 8910 53644
rect 11054 53592 11060 53644
rect 11112 53592 11118 53644
rect 12158 53592 12164 53644
rect 12216 53632 12222 53644
rect 12713 53635 12771 53641
rect 12713 53632 12725 53635
rect 12216 53604 12725 53632
rect 12216 53592 12222 53604
rect 12713 53601 12725 53604
rect 12759 53601 12771 53635
rect 24397 53635 24455 53641
rect 24397 53632 24409 53635
rect 12713 53595 12771 53601
rect 23308 53604 24409 53632
rect 6730 53524 6736 53576
rect 6788 53524 6794 53576
rect 8570 53524 8576 53576
rect 8628 53524 8634 53576
rect 9122 53524 9128 53576
rect 9180 53524 9186 53576
rect 11793 53567 11851 53573
rect 11793 53533 11805 53567
rect 11839 53564 11851 53567
rect 12066 53564 12072 53576
rect 11839 53536 12072 53564
rect 11839 53533 11851 53536
rect 11793 53527 11851 53533
rect 12066 53524 12072 53536
rect 12124 53524 12130 53576
rect 12437 53567 12495 53573
rect 12437 53533 12449 53567
rect 12483 53564 12495 53567
rect 12618 53564 12624 53576
rect 12483 53536 12624 53564
rect 12483 53533 12495 53536
rect 12437 53527 12495 53533
rect 12618 53524 12624 53536
rect 12676 53524 12682 53576
rect 13998 53524 14004 53576
rect 14056 53564 14062 53576
rect 14553 53567 14611 53573
rect 14553 53564 14565 53567
rect 14056 53536 14565 53564
rect 14056 53524 14062 53536
rect 14553 53533 14565 53536
rect 14599 53564 14611 53567
rect 14829 53567 14887 53573
rect 14829 53564 14841 53567
rect 14599 53536 14841 53564
rect 14599 53533 14611 53536
rect 14553 53527 14611 53533
rect 14829 53533 14841 53536
rect 14875 53533 14887 53567
rect 14829 53527 14887 53533
rect 15470 53524 15476 53576
rect 15528 53564 15534 53576
rect 15749 53567 15807 53573
rect 15749 53564 15761 53567
rect 15528 53536 15761 53564
rect 15528 53524 15534 53536
rect 15749 53533 15761 53536
rect 15795 53564 15807 53567
rect 16117 53567 16175 53573
rect 16117 53564 16129 53567
rect 15795 53536 16129 53564
rect 15795 53533 15807 53536
rect 15749 53527 15807 53533
rect 16117 53533 16129 53536
rect 16163 53533 16175 53567
rect 16117 53527 16175 53533
rect 16574 53524 16580 53576
rect 16632 53564 16638 53576
rect 16669 53567 16727 53573
rect 16669 53564 16681 53567
rect 16632 53536 16681 53564
rect 16632 53524 16638 53536
rect 16669 53533 16681 53536
rect 16715 53533 16727 53567
rect 16669 53527 16727 53533
rect 17310 53524 17316 53576
rect 17368 53564 17374 53576
rect 17405 53567 17463 53573
rect 17405 53564 17417 53567
rect 17368 53536 17417 53564
rect 17368 53524 17374 53536
rect 17405 53533 17417 53536
rect 17451 53533 17463 53567
rect 17405 53527 17463 53533
rect 18322 53524 18328 53576
rect 18380 53564 18386 53576
rect 18693 53567 18751 53573
rect 18693 53564 18705 53567
rect 18380 53536 18705 53564
rect 18380 53524 18386 53536
rect 18693 53533 18705 53536
rect 18739 53533 18751 53567
rect 18693 53527 18751 53533
rect 19150 53524 19156 53576
rect 19208 53564 19214 53576
rect 19429 53567 19487 53573
rect 19429 53564 19441 53567
rect 19208 53536 19441 53564
rect 19208 53524 19214 53536
rect 19429 53533 19441 53536
rect 19475 53533 19487 53567
rect 19429 53527 19487 53533
rect 19886 53524 19892 53576
rect 19944 53564 19950 53576
rect 20349 53567 20407 53573
rect 20349 53564 20361 53567
rect 19944 53536 20361 53564
rect 19944 53524 19950 53536
rect 20349 53533 20361 53536
rect 20395 53564 20407 53567
rect 20717 53567 20775 53573
rect 20717 53564 20729 53567
rect 20395 53536 20729 53564
rect 20395 53533 20407 53536
rect 20349 53527 20407 53533
rect 20717 53533 20729 53536
rect 20763 53533 20775 53567
rect 20717 53527 20775 53533
rect 20990 53524 20996 53576
rect 21048 53564 21054 53576
rect 21085 53567 21143 53573
rect 21085 53564 21097 53567
rect 21048 53536 21097 53564
rect 21048 53524 21054 53536
rect 21085 53533 21097 53536
rect 21131 53533 21143 53567
rect 21085 53527 21143 53533
rect 21726 53524 21732 53576
rect 21784 53564 21790 53576
rect 22005 53567 22063 53573
rect 22005 53564 22017 53567
rect 21784 53536 22017 53564
rect 21784 53524 21790 53536
rect 22005 53533 22017 53536
rect 22051 53533 22063 53567
rect 22005 53527 22063 53533
rect 22094 53524 22100 53576
rect 22152 53564 22158 53576
rect 22649 53567 22707 53573
rect 22649 53564 22661 53567
rect 22152 53536 22661 53564
rect 22152 53524 22158 53536
rect 22649 53533 22661 53536
rect 22695 53533 22707 53567
rect 22649 53527 22707 53533
rect 22830 53524 22836 53576
rect 22888 53564 22894 53576
rect 23308 53573 23336 53604
rect 24397 53601 24409 53604
rect 24443 53601 24455 53635
rect 24397 53595 24455 53601
rect 23293 53567 23351 53573
rect 23293 53564 23305 53567
rect 22888 53536 23305 53564
rect 22888 53524 22894 53536
rect 23293 53533 23305 53536
rect 23339 53533 23351 53567
rect 23293 53527 23351 53533
rect 23937 53567 23995 53573
rect 23937 53533 23949 53567
rect 23983 53564 23995 53567
rect 24486 53564 24492 53576
rect 23983 53536 24492 53564
rect 23983 53533 23995 53536
rect 23937 53527 23995 53533
rect 24486 53524 24492 53536
rect 24544 53524 24550 53576
rect 24762 53524 24768 53576
rect 24820 53564 24826 53576
rect 25225 53567 25283 53573
rect 25225 53564 25237 53567
rect 24820 53536 25237 53564
rect 24820 53524 24826 53536
rect 25225 53533 25237 53536
rect 25271 53533 25283 53567
rect 25225 53527 25283 53533
rect 7374 53496 7380 53508
rect 6288 53468 7380 53496
rect 7374 53456 7380 53468
rect 7432 53456 7438 53508
rect 7282 53428 7288 53440
rect 4448 53400 7288 53428
rect 3973 53391 4031 53397
rect 7282 53388 7288 53400
rect 7340 53388 7346 53440
rect 14369 53431 14427 53437
rect 14369 53397 14381 53431
rect 14415 53428 14427 53431
rect 14642 53428 14648 53440
rect 14415 53400 14648 53428
rect 14415 53397 14427 53400
rect 14369 53391 14427 53397
rect 14642 53388 14648 53400
rect 14700 53388 14706 53440
rect 15657 53431 15715 53437
rect 15657 53397 15669 53431
rect 15703 53428 15715 53431
rect 15838 53428 15844 53440
rect 15703 53400 15844 53428
rect 15703 53397 15715 53400
rect 15657 53391 15715 53397
rect 15838 53388 15844 53400
rect 15896 53388 15902 53440
rect 16853 53431 16911 53437
rect 16853 53397 16865 53431
rect 16899 53428 16911 53431
rect 17034 53428 17040 53440
rect 16899 53400 17040 53428
rect 16899 53397 16911 53400
rect 16853 53391 16911 53397
rect 17034 53388 17040 53400
rect 17092 53388 17098 53440
rect 17586 53388 17592 53440
rect 17644 53388 17650 53440
rect 18233 53431 18291 53437
rect 18233 53397 18245 53431
rect 18279 53428 18291 53431
rect 18322 53428 18328 53440
rect 18279 53400 18328 53428
rect 18279 53397 18291 53400
rect 18233 53391 18291 53397
rect 18322 53388 18328 53400
rect 18380 53388 18386 53440
rect 19610 53388 19616 53440
rect 19668 53388 19674 53440
rect 20257 53431 20315 53437
rect 20257 53397 20269 53431
rect 20303 53428 20315 53431
rect 20530 53428 20536 53440
rect 20303 53400 20536 53428
rect 20303 53397 20315 53400
rect 20257 53391 20315 53397
rect 20530 53388 20536 53400
rect 20588 53388 20594 53440
rect 21266 53388 21272 53440
rect 21324 53388 21330 53440
rect 21910 53388 21916 53440
rect 21968 53428 21974 53440
rect 22465 53431 22523 53437
rect 22465 53428 22477 53431
rect 21968 53400 22477 53428
rect 21968 53388 21974 53400
rect 22465 53397 22477 53400
rect 22511 53397 22523 53431
rect 22465 53391 22523 53397
rect 23842 53388 23848 53440
rect 23900 53388 23906 53440
rect 25130 53388 25136 53440
rect 25188 53388 25194 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 17310 53184 17316 53236
rect 17368 53184 17374 53236
rect 19150 53184 19156 53236
rect 19208 53224 19214 53236
rect 19521 53227 19579 53233
rect 19521 53224 19533 53227
rect 19208 53196 19533 53224
rect 19208 53184 19214 53196
rect 19521 53193 19533 53196
rect 19567 53193 19579 53227
rect 19521 53187 19579 53193
rect 19702 53184 19708 53236
rect 19760 53184 19766 53236
rect 20990 53184 20996 53236
rect 21048 53184 21054 53236
rect 21174 53184 21180 53236
rect 21232 53184 21238 53236
rect 21726 53184 21732 53236
rect 21784 53224 21790 53236
rect 21821 53227 21879 53233
rect 21821 53224 21833 53227
rect 21784 53196 21833 53224
rect 21784 53184 21790 53196
rect 21821 53193 21833 53196
rect 21867 53193 21879 53227
rect 21821 53187 21879 53193
rect 22094 53184 22100 53236
rect 22152 53224 22158 53236
rect 22281 53227 22339 53233
rect 22281 53224 22293 53227
rect 22152 53196 22293 53224
rect 22152 53184 22158 53196
rect 22281 53193 22293 53196
rect 22327 53193 22339 53227
rect 22281 53187 22339 53193
rect 22462 53184 22468 53236
rect 22520 53224 22526 53236
rect 22557 53227 22615 53233
rect 22557 53224 22569 53227
rect 22520 53196 22569 53224
rect 22520 53184 22526 53196
rect 22557 53193 22569 53196
rect 22603 53193 22615 53227
rect 22557 53187 22615 53193
rect 23017 53227 23075 53233
rect 23017 53193 23029 53227
rect 23063 53224 23075 53227
rect 23290 53224 23296 53236
rect 23063 53196 23296 53224
rect 23063 53193 23075 53196
rect 23017 53187 23075 53193
rect 23290 53184 23296 53196
rect 23348 53184 23354 53236
rect 13630 53116 13636 53168
rect 13688 53156 13694 53168
rect 13817 53159 13875 53165
rect 13817 53156 13829 53159
rect 13688 53128 13829 53156
rect 13688 53116 13694 53128
rect 13817 53125 13829 53128
rect 13863 53125 13875 53159
rect 13817 53119 13875 53125
rect 2317 53091 2375 53097
rect 2317 53057 2329 53091
rect 2363 53088 2375 53091
rect 2406 53088 2412 53100
rect 2363 53060 2412 53088
rect 2363 53057 2375 53060
rect 2317 53051 2375 53057
rect 2406 53048 2412 53060
rect 2464 53048 2470 53100
rect 4065 53091 4123 53097
rect 4065 53057 4077 53091
rect 4111 53088 4123 53091
rect 4246 53088 4252 53100
rect 4111 53060 4252 53088
rect 4111 53057 4123 53060
rect 4065 53051 4123 53057
rect 4246 53048 4252 53060
rect 4304 53048 4310 53100
rect 5997 53091 6055 53097
rect 5997 53057 6009 53091
rect 6043 53088 6055 53091
rect 6178 53088 6184 53100
rect 6043 53060 6184 53088
rect 6043 53057 6055 53060
rect 5997 53051 6055 53057
rect 6178 53048 6184 53060
rect 6236 53048 6242 53100
rect 7190 53048 7196 53100
rect 7248 53048 7254 53100
rect 8386 53048 8392 53100
rect 8444 53088 8450 53100
rect 9125 53091 9183 53097
rect 9125 53088 9137 53091
rect 8444 53060 9137 53088
rect 8444 53048 8450 53060
rect 9125 53057 9137 53060
rect 9171 53057 9183 53091
rect 9125 53051 9183 53057
rect 9490 53048 9496 53100
rect 9548 53088 9554 53100
rect 9769 53091 9827 53097
rect 9769 53088 9781 53091
rect 9548 53060 9781 53088
rect 9548 53048 9554 53060
rect 9769 53057 9781 53060
rect 9815 53057 9827 53091
rect 9769 53051 9827 53057
rect 11882 53048 11888 53100
rect 11940 53048 11946 53100
rect 14366 53048 14372 53100
rect 14424 53088 14430 53100
rect 14461 53091 14519 53097
rect 14461 53088 14473 53091
rect 14424 53060 14473 53088
rect 14424 53048 14430 53060
rect 14461 53057 14473 53060
rect 14507 53088 14519 53091
rect 14921 53091 14979 53097
rect 14921 53088 14933 53091
rect 14507 53060 14933 53088
rect 14507 53057 14519 53060
rect 14461 53051 14519 53057
rect 14921 53057 14933 53060
rect 14967 53057 14979 53091
rect 14921 53051 14979 53057
rect 15930 53048 15936 53100
rect 15988 53088 15994 53100
rect 16393 53091 16451 53097
rect 16393 53088 16405 53091
rect 15988 53060 16405 53088
rect 15988 53048 15994 53060
rect 16393 53057 16405 53060
rect 16439 53057 16451 53091
rect 16393 53051 16451 53057
rect 18782 53048 18788 53100
rect 18840 53088 18846 53100
rect 19061 53091 19119 53097
rect 19061 53088 19073 53091
rect 18840 53060 19073 53088
rect 18840 53048 18846 53060
rect 19061 53057 19073 53060
rect 19107 53088 19119 53091
rect 19337 53091 19395 53097
rect 19337 53088 19349 53091
rect 19107 53060 19349 53088
rect 19107 53057 19119 53060
rect 19061 53051 19119 53057
rect 19337 53057 19349 53060
rect 19383 53057 19395 53091
rect 19337 53051 19395 53057
rect 20254 53048 20260 53100
rect 20312 53088 20318 53100
rect 20533 53091 20591 53097
rect 20533 53088 20545 53091
rect 20312 53060 20545 53088
rect 20312 53048 20318 53060
rect 20533 53057 20545 53060
rect 20579 53088 20591 53091
rect 20809 53091 20867 53097
rect 20809 53088 20821 53091
rect 20579 53060 20821 53088
rect 20579 53057 20591 53060
rect 20533 53051 20591 53057
rect 20809 53057 20821 53060
rect 20855 53057 20867 53091
rect 23308 53088 23336 53184
rect 23477 53091 23535 53097
rect 23477 53088 23489 53091
rect 23308 53060 23489 53088
rect 20809 53051 20867 53057
rect 23477 53057 23489 53060
rect 23523 53057 23535 53091
rect 23477 53051 23535 53057
rect 23566 53048 23572 53100
rect 23624 53088 23630 53100
rect 24121 53091 24179 53097
rect 24121 53088 24133 53091
rect 23624 53060 24133 53088
rect 23624 53048 23630 53060
rect 24121 53057 24133 53060
rect 24167 53088 24179 53091
rect 24397 53091 24455 53097
rect 24397 53088 24409 53091
rect 24167 53060 24409 53088
rect 24167 53057 24179 53060
rect 24121 53051 24179 53057
rect 24397 53057 24409 53060
rect 24443 53057 24455 53091
rect 24397 53051 24455 53057
rect 24765 53091 24823 53097
rect 24765 53057 24777 53091
rect 24811 53088 24823 53091
rect 25314 53088 25320 53100
rect 24811 53060 25320 53088
rect 24811 53057 24823 53060
rect 24765 53051 24823 53057
rect 25314 53048 25320 53060
rect 25372 53048 25378 53100
rect 3697 53023 3755 53029
rect 3697 52989 3709 53023
rect 3743 53020 3755 53023
rect 4430 53020 4436 53032
rect 3743 52992 4436 53020
rect 3743 52989 3755 52992
rect 3697 52983 3755 52989
rect 4430 52980 4436 52992
rect 4488 52980 4494 53032
rect 5537 53023 5595 53029
rect 5537 52989 5549 53023
rect 5583 53020 5595 53023
rect 6270 53020 6276 53032
rect 5583 52992 6276 53020
rect 5583 52989 5595 52992
rect 5537 52983 5595 52989
rect 6270 52980 6276 52992
rect 6328 52980 6334 53032
rect 8849 53023 8907 53029
rect 8849 52989 8861 53023
rect 8895 53020 8907 53023
rect 9214 53020 9220 53032
rect 8895 52992 9220 53020
rect 8895 52989 8907 52992
rect 8849 52983 8907 52989
rect 9214 52980 9220 52992
rect 9272 52980 9278 53032
rect 10318 52980 10324 53032
rect 10376 52980 10382 53032
rect 11790 52980 11796 53032
rect 11848 53020 11854 53032
rect 12345 53023 12403 53029
rect 12345 53020 12357 53023
rect 11848 52992 12357 53020
rect 11848 52980 11854 52992
rect 12345 52989 12357 52992
rect 12391 52989 12403 53023
rect 12345 52983 12403 52989
rect 2958 52912 2964 52964
rect 3016 52952 3022 52964
rect 7834 52952 7840 52964
rect 3016 52924 7840 52952
rect 3016 52912 3022 52924
rect 7834 52912 7840 52924
rect 7892 52912 7898 52964
rect 13998 52912 14004 52964
rect 14056 52912 14062 52964
rect 14645 52955 14703 52961
rect 14645 52921 14657 52955
rect 14691 52952 14703 52955
rect 15562 52952 15568 52964
rect 14691 52924 15568 52952
rect 14691 52921 14703 52924
rect 14645 52915 14703 52921
rect 15562 52912 15568 52924
rect 15620 52912 15626 52964
rect 1578 52844 1584 52896
rect 1636 52884 1642 52896
rect 1673 52887 1731 52893
rect 1673 52884 1685 52887
rect 1636 52856 1685 52884
rect 1636 52844 1642 52856
rect 1673 52853 1685 52856
rect 1719 52853 1731 52887
rect 1673 52847 1731 52853
rect 6546 52844 6552 52896
rect 6604 52844 6610 52896
rect 16114 52844 16120 52896
rect 16172 52844 16178 52896
rect 18874 52844 18880 52896
rect 18932 52844 18938 52896
rect 20070 52844 20076 52896
rect 20128 52884 20134 52896
rect 20349 52887 20407 52893
rect 20349 52884 20361 52887
rect 20128 52856 20361 52884
rect 20128 52844 20134 52856
rect 20349 52853 20361 52856
rect 20395 52853 20407 52887
rect 20349 52847 20407 52853
rect 23290 52844 23296 52896
rect 23348 52844 23354 52896
rect 23382 52844 23388 52896
rect 23440 52884 23446 52896
rect 23937 52887 23995 52893
rect 23937 52884 23949 52887
rect 23440 52856 23949 52884
rect 23440 52844 23446 52856
rect 23937 52853 23949 52856
rect 23983 52853 23995 52887
rect 23937 52847 23995 52853
rect 25133 52887 25191 52893
rect 25133 52853 25145 52887
rect 25179 52884 25191 52887
rect 25682 52884 25688 52896
rect 25179 52856 25688 52884
rect 25179 52853 25191 52856
rect 25133 52847 25191 52853
rect 25682 52844 25688 52856
rect 25740 52844 25746 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 3694 52680 3700 52692
rect 2976 52652 3700 52680
rect 2976 52553 3004 52652
rect 3694 52640 3700 52652
rect 3752 52640 3758 52692
rect 4246 52640 4252 52692
rect 4304 52680 4310 52692
rect 9217 52683 9275 52689
rect 9217 52680 9229 52683
rect 4304 52652 9229 52680
rect 4304 52640 4310 52652
rect 9217 52649 9229 52652
rect 9263 52649 9275 52683
rect 9217 52643 9275 52649
rect 12618 52640 12624 52692
rect 12676 52640 12682 52692
rect 13630 52640 13636 52692
rect 13688 52680 13694 52692
rect 14093 52683 14151 52689
rect 14093 52680 14105 52683
rect 13688 52652 14105 52680
rect 13688 52640 13694 52652
rect 14093 52649 14105 52652
rect 14139 52649 14151 52683
rect 14093 52643 14151 52649
rect 24581 52683 24639 52689
rect 24581 52649 24593 52683
rect 24627 52680 24639 52683
rect 24762 52680 24768 52692
rect 24627 52652 24768 52680
rect 24627 52649 24639 52652
rect 24581 52643 24639 52649
rect 24762 52640 24768 52652
rect 24820 52640 24826 52692
rect 4982 52612 4988 52624
rect 3344 52584 4988 52612
rect 2961 52547 3019 52553
rect 2961 52513 2973 52547
rect 3007 52513 3019 52547
rect 2961 52507 3019 52513
rect 3344 52485 3372 52584
rect 4982 52572 4988 52584
rect 5040 52572 5046 52624
rect 25133 52615 25191 52621
rect 25133 52581 25145 52615
rect 25179 52612 25191 52615
rect 25774 52612 25780 52624
rect 25179 52584 25780 52612
rect 25179 52581 25191 52584
rect 25133 52575 25191 52581
rect 25774 52572 25780 52584
rect 25832 52572 25838 52624
rect 6273 52547 6331 52553
rect 6273 52513 6285 52547
rect 6319 52544 6331 52547
rect 6638 52544 6644 52556
rect 6319 52516 6644 52544
rect 6319 52513 6331 52516
rect 6273 52507 6331 52513
rect 6638 52504 6644 52516
rect 6696 52504 6702 52556
rect 7742 52504 7748 52556
rect 7800 52504 7806 52556
rect 10686 52504 10692 52556
rect 10744 52544 10750 52556
rect 11241 52547 11299 52553
rect 11241 52544 11253 52547
rect 10744 52516 11253 52544
rect 10744 52504 10750 52516
rect 11241 52513 11253 52516
rect 11287 52513 11299 52547
rect 11241 52507 11299 52513
rect 3329 52479 3387 52485
rect 3329 52445 3341 52479
rect 3375 52445 3387 52479
rect 3329 52439 3387 52445
rect 3418 52436 3424 52488
rect 3476 52476 3482 52488
rect 3973 52479 4031 52485
rect 3973 52476 3985 52479
rect 3476 52448 3985 52476
rect 3476 52436 3482 52448
rect 3973 52445 3985 52448
rect 4019 52445 4031 52479
rect 3973 52439 4031 52445
rect 6733 52479 6791 52485
rect 6733 52445 6745 52479
rect 6779 52476 6791 52479
rect 6822 52476 6828 52488
rect 6779 52448 6828 52476
rect 6779 52445 6791 52448
rect 6733 52439 6791 52445
rect 6822 52436 6828 52448
rect 6880 52436 6886 52488
rect 8573 52479 8631 52485
rect 8573 52445 8585 52479
rect 8619 52476 8631 52479
rect 8846 52476 8852 52488
rect 8619 52448 8852 52476
rect 8619 52445 8631 52448
rect 8573 52439 8631 52445
rect 8846 52436 8852 52448
rect 8904 52436 8910 52488
rect 9582 52436 9588 52488
rect 9640 52476 9646 52488
rect 10781 52479 10839 52485
rect 10781 52476 10793 52479
rect 9640 52448 10793 52476
rect 9640 52436 9646 52448
rect 10781 52445 10793 52448
rect 10827 52445 10839 52479
rect 10781 52439 10839 52445
rect 12802 52436 12808 52488
rect 12860 52436 12866 52488
rect 13633 52479 13691 52485
rect 13633 52445 13645 52479
rect 13679 52476 13691 52479
rect 16298 52476 16304 52488
rect 13679 52448 16304 52476
rect 13679 52445 13691 52448
rect 13633 52439 13691 52445
rect 16298 52436 16304 52448
rect 16356 52436 16362 52488
rect 24765 52479 24823 52485
rect 24765 52445 24777 52479
rect 24811 52476 24823 52479
rect 25314 52476 25320 52488
rect 24811 52448 25320 52476
rect 24811 52445 24823 52448
rect 24765 52439 24823 52445
rect 25314 52436 25320 52448
rect 25372 52436 25378 52488
rect 9306 52368 9312 52420
rect 9364 52368 9370 52420
rect 13354 52368 13360 52420
rect 13412 52408 13418 52420
rect 13449 52411 13507 52417
rect 13449 52408 13461 52411
rect 13412 52380 13461 52408
rect 13412 52368 13418 52380
rect 13449 52377 13461 52380
rect 13495 52377 13507 52411
rect 13449 52371 13507 52377
rect 4614 52300 4620 52352
rect 4672 52300 4678 52352
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 6546 52136 6552 52148
rect 3436 52108 6552 52136
rect 3237 52071 3295 52077
rect 3237 52037 3249 52071
rect 3283 52068 3295 52071
rect 3326 52068 3332 52080
rect 3283 52040 3332 52068
rect 3283 52037 3295 52040
rect 3237 52031 3295 52037
rect 3326 52028 3332 52040
rect 3384 52028 3390 52080
rect 1581 52003 1639 52009
rect 1581 51969 1593 52003
rect 1627 52000 1639 52003
rect 3436 52000 3464 52108
rect 6546 52096 6552 52108
rect 6604 52096 6610 52148
rect 7190 52096 7196 52148
rect 7248 52096 7254 52148
rect 11882 52096 11888 52148
rect 11940 52096 11946 52148
rect 12526 52096 12532 52148
rect 12584 52096 12590 52148
rect 13265 52139 13323 52145
rect 13265 52105 13277 52139
rect 13311 52136 13323 52139
rect 13354 52136 13360 52148
rect 13311 52108 13360 52136
rect 13311 52105 13323 52108
rect 13265 52099 13323 52105
rect 13354 52096 13360 52108
rect 13412 52096 13418 52148
rect 25222 52096 25228 52148
rect 25280 52096 25286 52148
rect 3878 52028 3884 52080
rect 3936 52068 3942 52080
rect 3936 52040 4752 52068
rect 3936 52028 3942 52040
rect 1627 51972 3464 52000
rect 4065 52003 4123 52009
rect 1627 51969 1639 51972
rect 1581 51963 1639 51969
rect 4065 51969 4077 52003
rect 4111 51969 4123 52003
rect 4724 52000 4752 52040
rect 4798 52028 4804 52080
rect 4856 52028 4862 52080
rect 7469 52071 7527 52077
rect 7469 52068 7481 52071
rect 5828 52040 7481 52068
rect 5828 52000 5856 52040
rect 4724 51972 5856 52000
rect 5997 52003 6055 52009
rect 4065 51963 4123 51969
rect 5997 51969 6009 52003
rect 6043 52000 6055 52003
rect 6454 52000 6460 52012
rect 6043 51972 6460 52000
rect 6043 51969 6055 51972
rect 5997 51963 6055 51969
rect 4080 51932 4108 51963
rect 6454 51960 6460 51972
rect 6512 51960 6518 52012
rect 6564 52009 6592 52040
rect 7469 52037 7481 52040
rect 7515 52037 7527 52071
rect 7469 52031 7527 52037
rect 9674 52028 9680 52080
rect 9732 52068 9738 52080
rect 9861 52071 9919 52077
rect 9861 52068 9873 52071
rect 9732 52040 9873 52068
rect 9732 52028 9738 52040
rect 9861 52037 9873 52040
rect 9907 52037 9919 52071
rect 9861 52031 9919 52037
rect 6549 52003 6607 52009
rect 6549 51969 6561 52003
rect 6595 52000 6607 52003
rect 6595 51972 6629 52000
rect 6595 51969 6607 51972
rect 6549 51963 6607 51969
rect 8754 51960 8760 52012
rect 8812 52000 8818 52012
rect 9033 52003 9091 52009
rect 9033 52000 9045 52003
rect 8812 51972 9045 52000
rect 8812 51960 8818 51972
rect 9033 51969 9045 51972
rect 9079 51969 9091 52003
rect 9033 51963 9091 51969
rect 10870 51960 10876 52012
rect 10928 51960 10934 52012
rect 11698 51960 11704 52012
rect 11756 51960 11762 52012
rect 12342 51960 12348 52012
rect 12400 51960 12406 52012
rect 4798 51932 4804 51944
rect 4080 51904 4804 51932
rect 4798 51892 4804 51904
rect 4856 51892 4862 51944
rect 8478 51892 8484 51944
rect 8536 51892 8542 51944
rect 2225 51867 2283 51873
rect 2225 51833 2237 51867
rect 2271 51864 2283 51867
rect 9122 51864 9128 51876
rect 2271 51836 9128 51864
rect 2271 51833 2283 51836
rect 2225 51827 2283 51833
rect 9122 51824 9128 51836
rect 9180 51824 9186 51876
rect 25314 51756 25320 51808
rect 25372 51796 25378 51808
rect 25409 51799 25467 51805
rect 25409 51796 25421 51799
rect 25372 51768 25421 51796
rect 25372 51756 25378 51768
rect 25409 51765 25421 51768
rect 25455 51765 25467 51799
rect 25409 51759 25467 51765
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 9950 51552 9956 51604
rect 10008 51592 10014 51604
rect 10229 51595 10287 51601
rect 10229 51592 10241 51595
rect 10008 51564 10241 51592
rect 10008 51552 10014 51564
rect 10229 51561 10241 51564
rect 10275 51561 10287 51595
rect 10229 51555 10287 51561
rect 2866 51416 2872 51468
rect 2924 51416 2930 51468
rect 5534 51416 5540 51468
rect 5592 51416 5598 51468
rect 7006 51416 7012 51468
rect 7064 51456 7070 51468
rect 7285 51459 7343 51465
rect 7285 51456 7297 51459
rect 7064 51428 7297 51456
rect 7064 51416 7070 51428
rect 7285 51425 7297 51428
rect 7331 51425 7343 51459
rect 7285 51419 7343 51425
rect 3421 51391 3479 51397
rect 3421 51357 3433 51391
rect 3467 51357 3479 51391
rect 3421 51351 3479 51357
rect 3436 51320 3464 51351
rect 4614 51348 4620 51400
rect 4672 51348 4678 51400
rect 6638 51348 6644 51400
rect 6696 51348 6702 51400
rect 8478 51348 8484 51400
rect 8536 51348 8542 51400
rect 9030 51348 9036 51400
rect 9088 51388 9094 51400
rect 10413 51391 10471 51397
rect 10413 51388 10425 51391
rect 9088 51360 10425 51388
rect 9088 51348 9094 51360
rect 10413 51357 10425 51360
rect 10459 51357 10471 51391
rect 10413 51351 10471 51357
rect 25314 51348 25320 51400
rect 25372 51348 25378 51400
rect 5534 51320 5540 51332
rect 3436 51292 5540 51320
rect 5534 51280 5540 51292
rect 5592 51280 5598 51332
rect 3970 51212 3976 51264
rect 4028 51212 4034 51264
rect 24854 51212 24860 51264
rect 24912 51252 24918 51264
rect 25133 51255 25191 51261
rect 25133 51252 25145 51255
rect 24912 51224 25145 51252
rect 24912 51212 24918 51224
rect 25133 51221 25145 51224
rect 25179 51221 25191 51255
rect 25133 51215 25191 51221
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 1765 51051 1823 51057
rect 1765 51017 1777 51051
rect 1811 51048 1823 51051
rect 3418 51048 3424 51060
rect 1811 51020 3424 51048
rect 1811 51017 1823 51020
rect 1765 51011 1823 51017
rect 3418 51008 3424 51020
rect 3476 51008 3482 51060
rect 5534 51008 5540 51060
rect 5592 51048 5598 51060
rect 7653 51051 7711 51057
rect 7653 51048 7665 51051
rect 5592 51020 7665 51048
rect 5592 51008 5598 51020
rect 7653 51017 7665 51020
rect 7699 51017 7711 51051
rect 7653 51011 7711 51017
rect 2774 50940 2780 50992
rect 2832 50940 2838 50992
rect 4154 50940 4160 50992
rect 4212 50980 4218 50992
rect 4341 50983 4399 50989
rect 4341 50980 4353 50983
rect 4212 50952 4353 50980
rect 4212 50940 4218 50952
rect 4341 50949 4353 50952
rect 4387 50949 4399 50983
rect 4341 50943 4399 50949
rect 6730 50940 6736 50992
rect 6788 50980 6794 50992
rect 6825 50983 6883 50989
rect 6825 50980 6837 50983
rect 6788 50952 6837 50980
rect 6788 50940 6794 50952
rect 6825 50949 6837 50952
rect 6871 50949 6883 50983
rect 6825 50943 6883 50949
rect 7834 50940 7840 50992
rect 7892 50980 7898 50992
rect 9401 50983 9459 50989
rect 9401 50980 9413 50983
rect 7892 50952 9413 50980
rect 7892 50940 7898 50952
rect 9401 50949 9413 50952
rect 9447 50949 9459 50983
rect 9401 50943 9459 50949
rect 9582 50940 9588 50992
rect 9640 50940 9646 50992
rect 1578 50872 1584 50924
rect 1636 50872 1642 50924
rect 3694 50872 3700 50924
rect 3752 50872 3758 50924
rect 5442 50872 5448 50924
rect 5500 50872 5506 50924
rect 6086 50872 6092 50924
rect 6144 50912 6150 50924
rect 7009 50915 7067 50921
rect 7009 50912 7021 50915
rect 6144 50884 7021 50912
rect 6144 50872 6150 50884
rect 7009 50881 7021 50884
rect 7055 50881 7067 50915
rect 7009 50875 7067 50881
rect 7745 50915 7803 50921
rect 7745 50881 7757 50915
rect 7791 50912 7803 50915
rect 9214 50912 9220 50924
rect 7791 50884 9220 50912
rect 7791 50881 7803 50884
rect 7745 50875 7803 50881
rect 9214 50872 9220 50884
rect 9272 50872 9278 50924
rect 24765 50915 24823 50921
rect 24765 50881 24777 50915
rect 24811 50912 24823 50915
rect 25314 50912 25320 50924
rect 24811 50884 25320 50912
rect 24811 50881 24823 50884
rect 24765 50875 24823 50881
rect 25314 50872 25320 50884
rect 25372 50872 25378 50924
rect 25133 50711 25191 50717
rect 25133 50677 25145 50711
rect 25179 50708 25191 50711
rect 25498 50708 25504 50720
rect 25179 50680 25504 50708
rect 25179 50677 25191 50680
rect 25133 50671 25191 50677
rect 25498 50668 25504 50680
rect 25556 50668 25562 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 8570 50464 8576 50516
rect 8628 50504 8634 50516
rect 9217 50507 9275 50513
rect 9217 50504 9229 50507
rect 8628 50476 9229 50504
rect 8628 50464 8634 50476
rect 9217 50473 9229 50476
rect 9263 50473 9275 50507
rect 9217 50467 9275 50473
rect 2222 50328 2228 50380
rect 2280 50328 2286 50380
rect 5626 50328 5632 50380
rect 5684 50368 5690 50380
rect 7193 50371 7251 50377
rect 7193 50368 7205 50371
rect 5684 50340 7205 50368
rect 5684 50328 5690 50340
rect 7193 50337 7205 50340
rect 7239 50337 7251 50371
rect 7193 50331 7251 50337
rect 24857 50371 24915 50377
rect 24857 50337 24869 50371
rect 24903 50368 24915 50371
rect 25406 50368 25412 50380
rect 24903 50340 25412 50368
rect 24903 50337 24915 50340
rect 24857 50331 24915 50337
rect 25406 50328 25412 50340
rect 25464 50328 25470 50380
rect 3421 50303 3479 50309
rect 3421 50269 3433 50303
rect 3467 50300 3479 50303
rect 3878 50300 3884 50312
rect 3467 50272 3884 50300
rect 3467 50269 3479 50272
rect 3421 50263 3479 50269
rect 3878 50260 3884 50272
rect 3936 50260 3942 50312
rect 3970 50260 3976 50312
rect 4028 50260 4034 50312
rect 7466 50260 7472 50312
rect 7524 50260 7530 50312
rect 9398 50260 9404 50312
rect 9456 50260 9462 50312
rect 24673 50303 24731 50309
rect 24673 50269 24685 50303
rect 24719 50300 24731 50303
rect 25314 50300 25320 50312
rect 24719 50272 25320 50300
rect 24719 50269 24731 50272
rect 24673 50263 24731 50269
rect 25314 50260 25320 50272
rect 25372 50260 25378 50312
rect 22066 50204 25176 50232
rect 4246 50124 4252 50176
rect 4304 50164 4310 50176
rect 4617 50167 4675 50173
rect 4617 50164 4629 50167
rect 4304 50136 4629 50164
rect 4304 50124 4310 50136
rect 4617 50133 4629 50136
rect 4663 50133 4675 50167
rect 4617 50127 4675 50133
rect 21542 50124 21548 50176
rect 21600 50164 21606 50176
rect 22066 50164 22094 50204
rect 25148 50173 25176 50204
rect 21600 50136 22094 50164
rect 25133 50167 25191 50173
rect 21600 50124 21606 50136
rect 25133 50133 25145 50167
rect 25179 50133 25191 50167
rect 25133 50127 25191 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 10042 49960 10048 49972
rect 3988 49932 10048 49960
rect 1854 49852 1860 49904
rect 1912 49892 1918 49904
rect 2133 49895 2191 49901
rect 2133 49892 2145 49895
rect 1912 49864 2145 49892
rect 1912 49852 1918 49864
rect 2133 49861 2145 49864
rect 2179 49861 2191 49895
rect 2133 49855 2191 49861
rect 3329 49827 3387 49833
rect 3329 49793 3341 49827
rect 3375 49824 3387 49827
rect 3418 49824 3424 49836
rect 3375 49796 3424 49824
rect 3375 49793 3387 49796
rect 3329 49787 3387 49793
rect 3418 49784 3424 49796
rect 3476 49784 3482 49836
rect 3988 49833 4016 49932
rect 10042 49920 10048 49932
rect 10100 49920 10106 49972
rect 11885 49963 11943 49969
rect 11885 49929 11897 49963
rect 11931 49960 11943 49963
rect 12342 49960 12348 49972
rect 11931 49932 12348 49960
rect 11931 49929 11943 49932
rect 11885 49923 11943 49929
rect 12342 49920 12348 49932
rect 12400 49920 12406 49972
rect 4246 49852 4252 49904
rect 4304 49852 4310 49904
rect 6365 49895 6423 49901
rect 6365 49892 6377 49895
rect 5474 49864 6377 49892
rect 6365 49861 6377 49864
rect 6411 49892 6423 49895
rect 6411 49864 9444 49892
rect 6411 49861 6423 49864
rect 6365 49855 6423 49861
rect 3973 49827 4031 49833
rect 3973 49793 3985 49827
rect 4019 49793 4031 49827
rect 3973 49787 4031 49793
rect 7742 49784 7748 49836
rect 7800 49824 7806 49836
rect 9309 49827 9367 49833
rect 9309 49824 9321 49827
rect 7800 49796 9321 49824
rect 7800 49784 7806 49796
rect 9309 49793 9321 49796
rect 9355 49793 9367 49827
rect 9416 49824 9444 49864
rect 9490 49852 9496 49904
rect 9548 49852 9554 49904
rect 11054 49824 11060 49836
rect 9416 49796 11060 49824
rect 9309 49787 9367 49793
rect 11054 49784 11060 49796
rect 11112 49784 11118 49836
rect 11422 49784 11428 49836
rect 11480 49824 11486 49836
rect 11701 49827 11759 49833
rect 11701 49824 11713 49827
rect 11480 49796 11713 49824
rect 11480 49784 11486 49796
rect 11701 49793 11713 49796
rect 11747 49793 11759 49827
rect 11701 49787 11759 49793
rect 5997 49759 6055 49765
rect 5997 49725 6009 49759
rect 6043 49756 6055 49759
rect 8570 49756 8576 49768
rect 6043 49728 8576 49756
rect 6043 49725 6055 49728
rect 5997 49719 6055 49725
rect 8570 49716 8576 49728
rect 8628 49716 8634 49768
rect 19794 49716 19800 49768
rect 19852 49756 19858 49768
rect 25041 49759 25099 49765
rect 25041 49756 25053 49759
rect 19852 49728 25053 49756
rect 19852 49716 19858 49728
rect 25041 49725 25053 49728
rect 25087 49725 25099 49759
rect 25041 49719 25099 49725
rect 25317 49759 25375 49765
rect 25317 49725 25329 49759
rect 25363 49756 25375 49759
rect 25406 49756 25412 49768
rect 25363 49728 25412 49756
rect 25363 49725 25375 49728
rect 25317 49719 25375 49725
rect 25406 49716 25412 49728
rect 25464 49716 25470 49768
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 12802 49376 12808 49428
rect 12860 49376 12866 49428
rect 1486 49240 1492 49292
rect 1544 49280 1550 49292
rect 1765 49283 1823 49289
rect 1765 49280 1777 49283
rect 1544 49252 1777 49280
rect 1544 49240 1550 49252
rect 1765 49249 1777 49252
rect 1811 49249 1823 49283
rect 1765 49243 1823 49249
rect 2961 49215 3019 49221
rect 2961 49181 2973 49215
rect 3007 49181 3019 49215
rect 2961 49175 3019 49181
rect 12989 49215 13047 49221
rect 12989 49181 13001 49215
rect 13035 49212 13047 49215
rect 13538 49212 13544 49224
rect 13035 49184 13544 49212
rect 13035 49181 13047 49184
rect 12989 49175 13047 49181
rect 2976 49076 3004 49175
rect 13538 49172 13544 49184
rect 13596 49172 13602 49224
rect 24857 49215 24915 49221
rect 24857 49181 24869 49215
rect 24903 49212 24915 49215
rect 25314 49212 25320 49224
rect 24903 49184 25320 49212
rect 24903 49181 24915 49184
rect 24857 49175 24915 49181
rect 25314 49172 25320 49184
rect 25372 49172 25378 49224
rect 22066 49116 25176 49144
rect 3329 49079 3387 49085
rect 3329 49076 3341 49079
rect 2976 49048 3341 49076
rect 3329 49045 3341 49048
rect 3375 49076 3387 49079
rect 3510 49076 3516 49088
rect 3375 49048 3516 49076
rect 3375 49045 3387 49048
rect 3329 49039 3387 49045
rect 3510 49036 3516 49048
rect 3568 49036 3574 49088
rect 18966 49036 18972 49088
rect 19024 49076 19030 49088
rect 22066 49076 22094 49116
rect 25148 49085 25176 49116
rect 19024 49048 22094 49076
rect 25133 49079 25191 49085
rect 19024 49036 19030 49048
rect 25133 49045 25145 49079
rect 25179 49045 25191 49079
rect 25133 49039 25191 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 25041 48739 25099 48745
rect 25041 48705 25053 48739
rect 25087 48736 25099 48739
rect 25866 48736 25872 48748
rect 25087 48708 25872 48736
rect 25087 48705 25099 48708
rect 25041 48699 25099 48705
rect 25866 48696 25872 48708
rect 25924 48696 25930 48748
rect 25222 48628 25228 48680
rect 25280 48668 25286 48680
rect 25317 48671 25375 48677
rect 25317 48668 25329 48671
rect 25280 48640 25329 48668
rect 25280 48628 25286 48640
rect 25317 48637 25329 48640
rect 25363 48637 25375 48671
rect 25317 48631 25375 48637
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 18322 48260 18328 48272
rect 17512 48232 18328 48260
rect 17310 48152 17316 48204
rect 17368 48152 17374 48204
rect 17512 48201 17540 48232
rect 18322 48220 18328 48232
rect 18380 48260 18386 48272
rect 18690 48260 18696 48272
rect 18380 48232 18696 48260
rect 18380 48220 18386 48232
rect 18690 48220 18696 48232
rect 18748 48220 18754 48272
rect 17497 48195 17555 48201
rect 17497 48161 17509 48195
rect 17543 48161 17555 48195
rect 17497 48155 17555 48161
rect 17586 48084 17592 48136
rect 17644 48084 17650 48136
rect 18782 48084 18788 48136
rect 18840 48124 18846 48136
rect 19429 48127 19487 48133
rect 19429 48124 19441 48127
rect 18840 48096 19441 48124
rect 18840 48084 18846 48096
rect 19429 48093 19441 48096
rect 19475 48093 19487 48127
rect 19429 48087 19487 48093
rect 17678 47948 17684 48000
rect 17736 47988 17742 48000
rect 17957 47991 18015 47997
rect 17957 47988 17969 47991
rect 17736 47960 17969 47988
rect 17736 47948 17742 47960
rect 17957 47957 17969 47960
rect 18003 47957 18015 47991
rect 17957 47951 18015 47957
rect 19518 47948 19524 48000
rect 19576 47988 19582 48000
rect 20073 47991 20131 47997
rect 20073 47988 20085 47991
rect 19576 47960 20085 47988
rect 19576 47948 19582 47960
rect 20073 47957 20085 47960
rect 20119 47957 20131 47991
rect 20073 47951 20131 47957
rect 25222 47948 25228 48000
rect 25280 47948 25286 48000
rect 25314 47948 25320 48000
rect 25372 47988 25378 48000
rect 25409 47991 25467 47997
rect 25409 47988 25421 47991
rect 25372 47960 25421 47988
rect 25372 47948 25378 47960
rect 25409 47957 25421 47960
rect 25455 47957 25467 47991
rect 25409 47951 25467 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9217 47787 9275 47793
rect 9217 47753 9229 47787
rect 9263 47784 9275 47787
rect 9306 47784 9312 47796
rect 9263 47756 9312 47784
rect 9263 47753 9275 47756
rect 9217 47747 9275 47753
rect 9306 47744 9312 47756
rect 9364 47744 9370 47796
rect 11698 47744 11704 47796
rect 11756 47784 11762 47796
rect 11885 47787 11943 47793
rect 11885 47784 11897 47787
rect 11756 47756 11897 47784
rect 11756 47744 11762 47756
rect 11885 47753 11897 47756
rect 11931 47753 11943 47787
rect 11885 47747 11943 47753
rect 16114 47744 16120 47796
rect 16172 47784 16178 47796
rect 17221 47787 17279 47793
rect 17221 47784 17233 47787
rect 16172 47756 17233 47784
rect 16172 47744 16178 47756
rect 17221 47753 17233 47756
rect 17267 47753 17279 47787
rect 17221 47747 17279 47753
rect 17313 47787 17371 47793
rect 17313 47753 17325 47787
rect 17359 47784 17371 47787
rect 18230 47784 18236 47796
rect 17359 47756 18236 47784
rect 17359 47753 17371 47756
rect 17313 47747 17371 47753
rect 18230 47744 18236 47756
rect 18288 47744 18294 47796
rect 19058 47676 19064 47728
rect 19116 47676 19122 47728
rect 19518 47676 19524 47728
rect 19576 47676 19582 47728
rect 9401 47651 9459 47657
rect 9401 47617 9413 47651
rect 9447 47648 9459 47651
rect 10962 47648 10968 47660
rect 9447 47620 10968 47648
rect 9447 47617 9459 47620
rect 9401 47611 9459 47617
rect 10962 47608 10968 47620
rect 11020 47608 11026 47660
rect 11698 47608 11704 47660
rect 11756 47608 11762 47660
rect 20162 47608 20168 47660
rect 20220 47648 20226 47660
rect 20257 47651 20315 47657
rect 20257 47648 20269 47651
rect 20220 47620 20269 47648
rect 20220 47608 20226 47620
rect 20257 47617 20269 47620
rect 20303 47617 20315 47651
rect 20257 47611 20315 47617
rect 17402 47540 17408 47592
rect 17460 47540 17466 47592
rect 19797 47583 19855 47589
rect 19797 47549 19809 47583
rect 19843 47549 19855 47583
rect 19797 47543 19855 47549
rect 16853 47447 16911 47453
rect 16853 47413 16865 47447
rect 16899 47444 16911 47447
rect 16942 47444 16948 47456
rect 16899 47416 16948 47444
rect 16899 47413 16911 47416
rect 16853 47407 16911 47413
rect 16942 47404 16948 47416
rect 17000 47404 17006 47456
rect 17770 47404 17776 47456
rect 17828 47444 17834 47456
rect 18049 47447 18107 47453
rect 18049 47444 18061 47447
rect 17828 47416 18061 47444
rect 17828 47404 17834 47416
rect 18049 47413 18061 47416
rect 18095 47413 18107 47447
rect 18049 47407 18107 47413
rect 19518 47404 19524 47456
rect 19576 47444 19582 47456
rect 19812 47444 19840 47543
rect 25038 47540 25044 47592
rect 25096 47540 25102 47592
rect 25314 47540 25320 47592
rect 25372 47540 25378 47592
rect 19576 47416 19840 47444
rect 19576 47404 19582 47416
rect 20714 47404 20720 47456
rect 20772 47444 20778 47456
rect 20901 47447 20959 47453
rect 20901 47444 20913 47447
rect 20772 47416 20913 47444
rect 20772 47404 20778 47416
rect 20901 47413 20913 47416
rect 20947 47413 20959 47447
rect 20901 47407 20959 47413
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 7377 47243 7435 47249
rect 7377 47209 7389 47243
rect 7423 47240 7435 47243
rect 7466 47240 7472 47252
rect 7423 47212 7472 47240
rect 7423 47209 7435 47212
rect 7377 47203 7435 47209
rect 7466 47200 7472 47212
rect 7524 47200 7530 47252
rect 17773 47243 17831 47249
rect 17773 47209 17785 47243
rect 17819 47240 17831 47243
rect 18230 47240 18236 47252
rect 17819 47212 18236 47240
rect 17819 47209 17831 47212
rect 17773 47203 17831 47209
rect 18230 47200 18236 47212
rect 18288 47200 18294 47252
rect 18506 47200 18512 47252
rect 18564 47240 18570 47252
rect 19334 47240 19340 47252
rect 18564 47212 19340 47240
rect 18564 47200 18570 47212
rect 19334 47200 19340 47212
rect 19392 47200 19398 47252
rect 20530 47200 20536 47252
rect 20588 47240 20594 47252
rect 20901 47243 20959 47249
rect 20901 47240 20913 47243
rect 20588 47212 20913 47240
rect 20588 47200 20594 47212
rect 20901 47209 20913 47212
rect 20947 47240 20959 47243
rect 20947 47212 21680 47240
rect 20947 47209 20959 47212
rect 20901 47203 20959 47209
rect 17494 47132 17500 47184
rect 17552 47172 17558 47184
rect 18141 47175 18199 47181
rect 18141 47172 18153 47175
rect 17552 47144 18153 47172
rect 17552 47132 17558 47144
rect 18141 47141 18153 47144
rect 18187 47141 18199 47175
rect 18141 47135 18199 47141
rect 19613 47175 19671 47181
rect 19613 47141 19625 47175
rect 19659 47172 19671 47175
rect 19886 47172 19892 47184
rect 19659 47144 19892 47172
rect 19659 47141 19671 47144
rect 19613 47135 19671 47141
rect 19886 47132 19892 47144
rect 19944 47132 19950 47184
rect 10042 47064 10048 47116
rect 10100 47064 10106 47116
rect 15470 47064 15476 47116
rect 15528 47104 15534 47116
rect 15657 47107 15715 47113
rect 15657 47104 15669 47107
rect 15528 47076 15669 47104
rect 15528 47064 15534 47076
rect 15657 47073 15669 47076
rect 15703 47073 15715 47107
rect 15657 47067 15715 47073
rect 16574 47064 16580 47116
rect 16632 47104 16638 47116
rect 16632 47076 17448 47104
rect 16632 47064 16638 47076
rect 7561 47039 7619 47045
rect 7561 47005 7573 47039
rect 7607 47036 7619 47039
rect 8938 47036 8944 47048
rect 7607 47008 8944 47036
rect 7607 47005 7619 47008
rect 7561 46999 7619 47005
rect 8938 46996 8944 47008
rect 8996 46996 9002 47048
rect 17420 47045 17448 47076
rect 18782 47064 18788 47116
rect 18840 47064 18846 47116
rect 20070 47064 20076 47116
rect 20128 47064 20134 47116
rect 20162 47064 20168 47116
rect 20220 47064 20226 47116
rect 21453 47107 21511 47113
rect 21453 47073 21465 47107
rect 21499 47104 21511 47107
rect 21542 47104 21548 47116
rect 21499 47076 21548 47104
rect 21499 47073 21511 47076
rect 21453 47067 21511 47073
rect 21542 47064 21548 47076
rect 21600 47064 21606 47116
rect 12253 47039 12311 47045
rect 12253 47036 12265 47039
rect 11808 47008 12265 47036
rect 10318 46928 10324 46980
rect 10376 46928 10382 46980
rect 11054 46928 11060 46980
rect 11112 46928 11118 46980
rect 11808 46912 11836 47008
rect 12253 47005 12265 47008
rect 12299 47005 12311 47039
rect 12253 46999 12311 47005
rect 17405 47039 17463 47045
rect 17405 47005 17417 47039
rect 17451 47036 17463 47039
rect 18598 47036 18604 47048
rect 17451 47008 18604 47036
rect 17451 47005 17463 47008
rect 17405 46999 17463 47005
rect 18598 46996 18604 47008
rect 18656 46996 18662 47048
rect 19610 46996 19616 47048
rect 19668 47036 19674 47048
rect 21652 47045 21680 47212
rect 22005 47175 22063 47181
rect 22005 47141 22017 47175
rect 22051 47172 22063 47175
rect 22462 47172 22468 47184
rect 22051 47144 22468 47172
rect 22051 47141 22063 47144
rect 22005 47135 22063 47141
rect 22462 47132 22468 47144
rect 22520 47132 22526 47184
rect 23753 47107 23811 47113
rect 23753 47073 23765 47107
rect 23799 47104 23811 47107
rect 24118 47104 24124 47116
rect 23799 47076 24124 47104
rect 23799 47073 23811 47076
rect 23753 47067 23811 47073
rect 24118 47064 24124 47076
rect 24176 47064 24182 47116
rect 19981 47039 20039 47045
rect 19981 47036 19993 47039
rect 19668 47008 19993 47036
rect 19668 46996 19674 47008
rect 19981 47005 19993 47008
rect 20027 47036 20039 47039
rect 20625 47039 20683 47045
rect 20625 47036 20637 47039
rect 20027 47008 20637 47036
rect 20027 47005 20039 47008
rect 19981 46999 20039 47005
rect 20625 47005 20637 47008
rect 20671 47005 20683 47039
rect 20625 46999 20683 47005
rect 21637 47039 21695 47045
rect 21637 47005 21649 47039
rect 21683 47005 21695 47039
rect 21637 46999 21695 47005
rect 24029 47039 24087 47045
rect 24029 47005 24041 47039
rect 24075 47005 24087 47039
rect 24029 46999 24087 47005
rect 16698 46940 16804 46968
rect 11790 46860 11796 46912
rect 11848 46860 11854 46912
rect 12802 46860 12808 46912
rect 12860 46900 12866 46912
rect 12897 46903 12955 46909
rect 12897 46900 12909 46903
rect 12860 46872 12909 46900
rect 12860 46860 12866 46872
rect 12897 46869 12909 46872
rect 12943 46869 12955 46903
rect 12897 46863 12955 46869
rect 14182 46860 14188 46912
rect 14240 46860 14246 46912
rect 16776 46900 16804 46940
rect 17126 46928 17132 46980
rect 17184 46928 17190 46980
rect 18506 46928 18512 46980
rect 18564 46928 18570 46980
rect 18874 46968 18880 46980
rect 18616 46940 18880 46968
rect 16850 46900 16856 46912
rect 16776 46872 16856 46900
rect 16850 46860 16856 46872
rect 16908 46900 16914 46912
rect 17862 46900 17868 46912
rect 16908 46872 17868 46900
rect 16908 46860 16914 46872
rect 17862 46860 17868 46872
rect 17920 46860 17926 46912
rect 18616 46909 18644 46940
rect 18874 46928 18880 46940
rect 18932 46928 18938 46980
rect 21545 46971 21603 46977
rect 21545 46937 21557 46971
rect 21591 46968 21603 46971
rect 21910 46968 21916 46980
rect 21591 46940 21916 46968
rect 21591 46937 21603 46940
rect 21545 46931 21603 46937
rect 21910 46928 21916 46940
rect 21968 46928 21974 46980
rect 24044 46968 24072 46999
rect 24486 46968 24492 46980
rect 24044 46940 24492 46968
rect 24486 46928 24492 46940
rect 24544 46928 24550 46980
rect 18601 46903 18659 46909
rect 18601 46869 18613 46903
rect 18647 46869 18659 46903
rect 18601 46863 18659 46869
rect 25314 46860 25320 46912
rect 25372 46900 25378 46912
rect 25409 46903 25467 46909
rect 25409 46900 25421 46903
rect 25372 46872 25421 46900
rect 25372 46860 25378 46872
rect 25409 46869 25421 46872
rect 25455 46869 25467 46903
rect 25409 46863 25467 46869
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 9030 46656 9036 46708
rect 9088 46656 9094 46708
rect 9214 46656 9220 46708
rect 9272 46696 9278 46708
rect 10597 46699 10655 46705
rect 10597 46696 10609 46699
rect 9272 46668 10609 46696
rect 9272 46656 9278 46668
rect 10597 46665 10609 46668
rect 10643 46665 10655 46699
rect 10597 46659 10655 46665
rect 11054 46656 11060 46708
rect 11112 46696 11118 46708
rect 11885 46699 11943 46705
rect 11885 46696 11897 46699
rect 11112 46668 11897 46696
rect 11112 46656 11118 46668
rect 11885 46665 11897 46668
rect 11931 46665 11943 46699
rect 14090 46696 14096 46708
rect 11885 46659 11943 46665
rect 12544 46668 14096 46696
rect 6822 46588 6828 46640
rect 6880 46628 6886 46640
rect 8021 46631 8079 46637
rect 8021 46628 8033 46631
rect 6880 46600 8033 46628
rect 6880 46588 6886 46600
rect 8021 46597 8033 46600
rect 8067 46597 8079 46631
rect 8021 46591 8079 46597
rect 8205 46563 8263 46569
rect 8205 46560 8217 46563
rect 7668 46532 8217 46560
rect 7374 46316 7380 46368
rect 7432 46356 7438 46368
rect 7668 46365 7696 46532
rect 8205 46529 8217 46532
rect 8251 46529 8263 46563
rect 8205 46523 8263 46529
rect 8849 46563 8907 46569
rect 8849 46529 8861 46563
rect 8895 46560 8907 46563
rect 9122 46560 9128 46572
rect 8895 46532 9128 46560
rect 8895 46529 8907 46532
rect 8849 46523 8907 46529
rect 9122 46520 9128 46532
rect 9180 46520 9186 46572
rect 10781 46563 10839 46569
rect 10781 46529 10793 46563
rect 10827 46560 10839 46563
rect 12544 46560 12572 46668
rect 14090 46656 14096 46668
rect 14148 46656 14154 46708
rect 16301 46699 16359 46705
rect 15212 46668 16160 46696
rect 14182 46628 14188 46640
rect 13386 46600 14188 46628
rect 14182 46588 14188 46600
rect 14240 46588 14246 46640
rect 15212 46628 15240 46668
rect 16132 46640 16160 46668
rect 16301 46665 16313 46699
rect 16347 46696 16359 46699
rect 17402 46696 17408 46708
rect 16347 46668 17408 46696
rect 16347 46665 16359 46668
rect 16301 46659 16359 46665
rect 17402 46656 17408 46668
rect 17460 46656 17466 46708
rect 18782 46656 18788 46708
rect 18840 46696 18846 46708
rect 19061 46699 19119 46705
rect 19061 46696 19073 46699
rect 18840 46668 19073 46696
rect 18840 46656 18846 46668
rect 19061 46665 19073 46668
rect 19107 46665 19119 46699
rect 19061 46659 19119 46665
rect 19150 46656 19156 46708
rect 19208 46696 19214 46708
rect 22649 46699 22707 46705
rect 19208 46668 20208 46696
rect 19208 46656 19214 46668
rect 15286 46628 15292 46640
rect 15212 46600 15292 46628
rect 15286 46588 15292 46600
rect 15344 46588 15350 46640
rect 16114 46588 16120 46640
rect 16172 46628 16178 46640
rect 16850 46628 16856 46640
rect 16172 46600 16856 46628
rect 16172 46588 16178 46600
rect 16850 46588 16856 46600
rect 16908 46588 16914 46640
rect 17862 46588 17868 46640
rect 17920 46628 17926 46640
rect 19168 46628 19196 46656
rect 20180 46628 20208 46668
rect 22649 46665 22661 46699
rect 22695 46696 22707 46699
rect 23382 46696 23388 46708
rect 22695 46668 23388 46696
rect 22695 46665 22707 46668
rect 22649 46659 22707 46665
rect 23382 46656 23388 46668
rect 23440 46656 23446 46708
rect 22097 46631 22155 46637
rect 17920 46600 19196 46628
rect 20102 46600 20852 46628
rect 17920 46588 17926 46600
rect 10827 46532 12572 46560
rect 10827 46529 10839 46532
rect 10781 46523 10839 46529
rect 18598 46520 18604 46572
rect 18656 46520 18662 46572
rect 20824 46560 20852 46600
rect 22097 46597 22109 46631
rect 22143 46628 22155 46631
rect 22186 46628 22192 46640
rect 22143 46600 22192 46628
rect 22143 46597 22155 46600
rect 22097 46591 22155 46597
rect 22186 46588 22192 46600
rect 22244 46628 22250 46640
rect 22244 46600 22784 46628
rect 22244 46588 22250 46600
rect 22756 46572 22784 46600
rect 20824 46532 22692 46560
rect 13814 46452 13820 46504
rect 13872 46452 13878 46504
rect 14093 46495 14151 46501
rect 14093 46461 14105 46495
rect 14139 46492 14151 46495
rect 14553 46495 14611 46501
rect 14553 46492 14565 46495
rect 14139 46464 14565 46492
rect 14139 46461 14151 46464
rect 14093 46455 14151 46461
rect 14553 46461 14565 46464
rect 14599 46461 14611 46495
rect 14553 46455 14611 46461
rect 14829 46495 14887 46501
rect 14829 46461 14841 46495
rect 14875 46492 14887 46495
rect 16666 46492 16672 46504
rect 14875 46464 16672 46492
rect 14875 46461 14887 46464
rect 14829 46455 14887 46461
rect 7653 46359 7711 46365
rect 7653 46356 7665 46359
rect 7432 46328 7665 46356
rect 7432 46316 7438 46328
rect 7653 46325 7665 46328
rect 7699 46325 7711 46359
rect 7653 46319 7711 46325
rect 12345 46359 12403 46365
rect 12345 46325 12357 46359
rect 12391 46356 12403 46359
rect 12434 46356 12440 46368
rect 12391 46328 12440 46356
rect 12391 46325 12403 46328
rect 12345 46319 12403 46325
rect 12434 46316 12440 46328
rect 12492 46316 12498 46368
rect 12526 46316 12532 46368
rect 12584 46356 12590 46368
rect 14108 46356 14136 46455
rect 16666 46452 16672 46464
rect 16724 46452 16730 46504
rect 18322 46452 18328 46504
rect 18380 46452 18386 46504
rect 20533 46495 20591 46501
rect 20533 46492 20545 46495
rect 19536 46464 20545 46492
rect 19536 46368 19564 46464
rect 20533 46461 20545 46464
rect 20579 46461 20591 46495
rect 20533 46455 20591 46461
rect 20809 46495 20867 46501
rect 20809 46461 20821 46495
rect 20855 46492 20867 46495
rect 21174 46492 21180 46504
rect 20855 46464 21180 46492
rect 20855 46461 20867 46464
rect 20809 46455 20867 46461
rect 21174 46452 21180 46464
rect 21232 46452 21238 46504
rect 22554 46452 22560 46504
rect 22612 46452 22618 46504
rect 22664 46492 22692 46532
rect 22738 46520 22744 46572
rect 22796 46520 22802 46572
rect 25041 46563 25099 46569
rect 25041 46529 25053 46563
rect 25087 46560 25099 46563
rect 25958 46560 25964 46572
rect 25087 46532 25964 46560
rect 25087 46529 25099 46532
rect 25041 46523 25099 46529
rect 25958 46520 25964 46532
rect 26016 46520 26022 46572
rect 23658 46492 23664 46504
rect 22664 46464 23664 46492
rect 23658 46452 23664 46464
rect 23716 46452 23722 46504
rect 25314 46452 25320 46504
rect 25372 46452 25378 46504
rect 12584 46328 14136 46356
rect 16853 46359 16911 46365
rect 12584 46316 12590 46328
rect 16853 46325 16865 46359
rect 16899 46356 16911 46359
rect 17310 46356 17316 46368
rect 16899 46328 17316 46356
rect 16899 46325 16911 46328
rect 16853 46319 16911 46325
rect 17310 46316 17316 46328
rect 17368 46356 17374 46368
rect 17586 46356 17592 46368
rect 17368 46328 17592 46356
rect 17368 46316 17374 46328
rect 17586 46316 17592 46328
rect 17644 46316 17650 46368
rect 19518 46316 19524 46368
rect 19576 46316 19582 46368
rect 23109 46359 23167 46365
rect 23109 46325 23121 46359
rect 23155 46356 23167 46359
rect 25038 46356 25044 46368
rect 23155 46328 25044 46356
rect 23155 46325 23167 46328
rect 23109 46319 23167 46325
rect 25038 46316 25044 46328
rect 25096 46316 25102 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 11422 46112 11428 46164
rect 11480 46112 11486 46164
rect 14182 46112 14188 46164
rect 14240 46112 14246 46164
rect 16206 46112 16212 46164
rect 16264 46152 16270 46164
rect 16482 46152 16488 46164
rect 16264 46124 16488 46152
rect 16264 46112 16270 46124
rect 16482 46112 16488 46124
rect 16540 46112 16546 46164
rect 16666 46112 16672 46164
rect 16724 46112 16730 46164
rect 17126 46112 17132 46164
rect 17184 46152 17190 46164
rect 17773 46155 17831 46161
rect 17773 46152 17785 46155
rect 17184 46124 17785 46152
rect 17184 46112 17190 46124
rect 17773 46121 17785 46124
rect 17819 46121 17831 46155
rect 17773 46115 17831 46121
rect 6178 46044 6184 46096
rect 6236 46084 6242 46096
rect 7745 46087 7803 46093
rect 7745 46084 7757 46087
rect 6236 46056 7757 46084
rect 6236 46044 6242 46056
rect 7745 46053 7757 46056
rect 7791 46053 7803 46087
rect 7745 46047 7803 46053
rect 8478 46044 8484 46096
rect 8536 46084 8542 46096
rect 9125 46087 9183 46093
rect 9125 46084 9137 46087
rect 8536 46056 9137 46084
rect 8536 46044 8542 46056
rect 9125 46053 9137 46056
rect 9171 46053 9183 46087
rect 9125 46047 9183 46053
rect 10873 46019 10931 46025
rect 10873 45985 10885 46019
rect 10919 46016 10931 46019
rect 11790 46016 11796 46028
rect 10919 45988 11796 46016
rect 10919 45985 10931 45988
rect 10873 45979 10931 45985
rect 11790 45976 11796 45988
rect 11848 45976 11854 46028
rect 11885 46019 11943 46025
rect 11885 45985 11897 46019
rect 11931 46016 11943 46019
rect 12526 46016 12532 46028
rect 11931 45988 12532 46016
rect 11931 45985 11943 45988
rect 11885 45979 11943 45985
rect 12526 45976 12532 45988
rect 12584 46016 12590 46028
rect 12710 46016 12716 46028
rect 12584 45988 12716 46016
rect 12584 45976 12590 45988
rect 12710 45976 12716 45988
rect 12768 45976 12774 46028
rect 16206 45976 16212 46028
rect 16264 45976 16270 46028
rect 20622 45976 20628 46028
rect 20680 46016 20686 46028
rect 20717 46019 20775 46025
rect 20717 46016 20729 46019
rect 20680 45988 20729 46016
rect 20680 45976 20686 45988
rect 20717 45985 20729 45988
rect 20763 45985 20775 46019
rect 20717 45979 20775 45985
rect 20901 46019 20959 46025
rect 20901 45985 20913 46019
rect 20947 46016 20959 46019
rect 21910 46016 21916 46028
rect 20947 45988 21916 46016
rect 20947 45985 20959 45988
rect 20901 45979 20959 45985
rect 21910 45976 21916 45988
rect 21968 45976 21974 46028
rect 22370 45976 22376 46028
rect 22428 46016 22434 46028
rect 22428 45988 24624 46016
rect 22428 45976 22434 45988
rect 17034 45908 17040 45960
rect 17092 45948 17098 45960
rect 17313 45951 17371 45957
rect 17313 45948 17325 45951
rect 17092 45920 17325 45948
rect 17092 45908 17098 45920
rect 17313 45917 17325 45920
rect 17359 45917 17371 45951
rect 17313 45911 17371 45917
rect 17586 45908 17592 45960
rect 17644 45948 17650 45960
rect 18417 45951 18475 45957
rect 18417 45948 18429 45951
rect 17644 45920 18429 45948
rect 17644 45908 17650 45920
rect 18417 45917 18429 45920
rect 18463 45917 18475 45951
rect 18417 45911 18475 45917
rect 24026 45908 24032 45960
rect 24084 45908 24090 45960
rect 24596 45957 24624 45988
rect 24581 45951 24639 45957
rect 24581 45917 24593 45951
rect 24627 45917 24639 45951
rect 24581 45911 24639 45917
rect 7929 45883 7987 45889
rect 7929 45849 7941 45883
rect 7975 45849 7987 45883
rect 7929 45843 7987 45849
rect 9309 45883 9367 45889
rect 9309 45849 9321 45883
rect 9355 45849 9367 45883
rect 9309 45843 9367 45849
rect 10965 45883 11023 45889
rect 10965 45849 10977 45883
rect 11011 45880 11023 45883
rect 11882 45880 11888 45892
rect 11011 45852 11888 45880
rect 11011 45849 11023 45852
rect 10965 45843 11023 45849
rect 7944 45812 7972 45843
rect 8389 45815 8447 45821
rect 8389 45812 8401 45815
rect 7944 45784 8401 45812
rect 8389 45781 8401 45784
rect 8435 45812 8447 45815
rect 8754 45812 8760 45824
rect 8435 45784 8760 45812
rect 8435 45781 8447 45784
rect 8389 45775 8447 45781
rect 8754 45772 8760 45784
rect 8812 45772 8818 45824
rect 9324 45812 9352 45843
rect 11882 45840 11888 45852
rect 11940 45840 11946 45892
rect 12161 45883 12219 45889
rect 12161 45849 12173 45883
rect 12207 45880 12219 45883
rect 14182 45880 14188 45892
rect 12207 45852 12434 45880
rect 13386 45852 14188 45880
rect 12207 45849 12219 45852
rect 12161 45843 12219 45849
rect 9674 45812 9680 45824
rect 9324 45784 9680 45812
rect 9674 45772 9680 45784
rect 9732 45772 9738 45824
rect 11057 45815 11115 45821
rect 11057 45781 11069 45815
rect 11103 45812 11115 45815
rect 11422 45812 11428 45824
rect 11103 45784 11428 45812
rect 11103 45781 11115 45784
rect 11057 45775 11115 45781
rect 11422 45772 11428 45784
rect 11480 45772 11486 45824
rect 12406 45812 12434 45852
rect 14182 45840 14188 45852
rect 14240 45880 14246 45892
rect 14550 45880 14556 45892
rect 14240 45852 14556 45880
rect 14240 45840 14246 45852
rect 14550 45840 14556 45852
rect 14608 45840 14614 45892
rect 15378 45840 15384 45892
rect 15436 45840 15442 45892
rect 15933 45883 15991 45889
rect 15933 45849 15945 45883
rect 15979 45880 15991 45883
rect 16850 45880 16856 45892
rect 15979 45852 16856 45880
rect 15979 45849 15991 45852
rect 15933 45843 15991 45849
rect 16850 45840 16856 45852
rect 16908 45840 16914 45892
rect 19242 45840 19248 45892
rect 19300 45880 19306 45892
rect 20438 45880 20444 45892
rect 19300 45852 20444 45880
rect 19300 45840 19306 45852
rect 20438 45840 20444 45852
rect 20496 45880 20502 45892
rect 20625 45883 20683 45889
rect 20625 45880 20637 45883
rect 20496 45852 20637 45880
rect 20496 45840 20502 45852
rect 20625 45849 20637 45852
rect 20671 45880 20683 45883
rect 21269 45883 21327 45889
rect 21269 45880 21281 45883
rect 20671 45852 21281 45880
rect 20671 45849 20683 45852
rect 20625 45843 20683 45849
rect 21269 45849 21281 45852
rect 21315 45849 21327 45883
rect 23658 45880 23664 45892
rect 23322 45852 23664 45880
rect 21269 45843 21327 45849
rect 23658 45840 23664 45852
rect 23716 45840 23722 45892
rect 23753 45883 23811 45889
rect 23753 45849 23765 45883
rect 23799 45880 23811 45883
rect 24946 45880 24952 45892
rect 23799 45852 24952 45880
rect 23799 45849 23811 45852
rect 23753 45843 23811 45849
rect 24946 45840 24952 45852
rect 25004 45840 25010 45892
rect 12802 45812 12808 45824
rect 12406 45784 12808 45812
rect 12802 45772 12808 45784
rect 12860 45772 12866 45824
rect 13446 45772 13452 45824
rect 13504 45812 13510 45824
rect 13633 45815 13691 45821
rect 13633 45812 13645 45815
rect 13504 45784 13645 45812
rect 13504 45772 13510 45784
rect 13633 45781 13645 45784
rect 13679 45781 13691 45815
rect 13633 45775 13691 45781
rect 14461 45815 14519 45821
rect 14461 45781 14473 45815
rect 14507 45812 14519 45815
rect 14918 45812 14924 45824
rect 14507 45784 14924 45812
rect 14507 45781 14519 45784
rect 14461 45775 14519 45781
rect 14918 45772 14924 45784
rect 14976 45772 14982 45824
rect 16114 45772 16120 45824
rect 16172 45812 16178 45824
rect 16574 45812 16580 45824
rect 16172 45784 16580 45812
rect 16172 45772 16178 45784
rect 16574 45772 16580 45784
rect 16632 45772 16638 45824
rect 20254 45772 20260 45824
rect 20312 45772 20318 45824
rect 22281 45815 22339 45821
rect 22281 45781 22293 45815
rect 22327 45812 22339 45815
rect 22370 45812 22376 45824
rect 22327 45784 22376 45812
rect 22327 45781 22339 45784
rect 22281 45775 22339 45781
rect 22370 45772 22376 45784
rect 22428 45772 22434 45824
rect 23474 45772 23480 45824
rect 23532 45812 23538 45824
rect 25225 45815 25283 45821
rect 25225 45812 25237 45815
rect 23532 45784 25237 45812
rect 23532 45772 23538 45784
rect 25225 45781 25237 45784
rect 25271 45781 25283 45815
rect 25225 45775 25283 45781
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 3970 45568 3976 45620
rect 4028 45608 4034 45620
rect 9490 45608 9496 45620
rect 4028 45580 9496 45608
rect 4028 45568 4034 45580
rect 9490 45568 9496 45580
rect 9548 45568 9554 45620
rect 11054 45568 11060 45620
rect 11112 45608 11118 45620
rect 11241 45611 11299 45617
rect 11241 45608 11253 45611
rect 11112 45580 11253 45608
rect 11112 45568 11118 45580
rect 11241 45577 11253 45580
rect 11287 45577 11299 45611
rect 11241 45571 11299 45577
rect 13814 45568 13820 45620
rect 13872 45608 13878 45620
rect 14553 45611 14611 45617
rect 14553 45608 14565 45611
rect 13872 45580 14565 45608
rect 13872 45568 13878 45580
rect 14553 45577 14565 45580
rect 14599 45577 14611 45611
rect 14553 45571 14611 45577
rect 18141 45611 18199 45617
rect 18141 45577 18153 45611
rect 18187 45608 18199 45611
rect 18322 45608 18328 45620
rect 18187 45580 18328 45608
rect 18187 45577 18199 45580
rect 18141 45571 18199 45577
rect 18322 45568 18328 45580
rect 18380 45568 18386 45620
rect 8570 45500 8576 45552
rect 8628 45540 8634 45552
rect 8665 45543 8723 45549
rect 8665 45540 8677 45543
rect 8628 45512 8677 45540
rect 8628 45500 8634 45512
rect 8665 45509 8677 45512
rect 8711 45540 8723 45543
rect 9306 45540 9312 45552
rect 8711 45512 9312 45540
rect 8711 45509 8723 45512
rect 8665 45503 8723 45509
rect 9306 45500 9312 45512
rect 9364 45500 9370 45552
rect 11072 45540 11100 45568
rect 10534 45512 11100 45540
rect 11514 45500 11520 45552
rect 11572 45540 11578 45552
rect 11701 45543 11759 45549
rect 11701 45540 11713 45543
rect 11572 45512 11713 45540
rect 11572 45500 11578 45512
rect 11701 45509 11713 45512
rect 11747 45509 11759 45543
rect 11701 45503 11759 45509
rect 16850 45500 16856 45552
rect 16908 45500 16914 45552
rect 20622 45540 20628 45552
rect 20286 45512 20628 45540
rect 20622 45500 20628 45512
rect 20680 45500 20686 45552
rect 20714 45500 20720 45552
rect 20772 45500 20778 45552
rect 23382 45540 23388 45552
rect 23046 45512 23388 45540
rect 23382 45500 23388 45512
rect 23440 45500 23446 45552
rect 23474 45500 23480 45552
rect 23532 45500 23538 45552
rect 11885 45475 11943 45481
rect 11885 45441 11897 45475
rect 11931 45472 11943 45475
rect 12250 45472 12256 45484
rect 11931 45444 12256 45472
rect 11931 45441 11943 45444
rect 11885 45435 11943 45441
rect 12250 45432 12256 45444
rect 12308 45432 12314 45484
rect 13722 45432 13728 45484
rect 13780 45432 13786 45484
rect 14734 45432 14740 45484
rect 14792 45472 14798 45484
rect 15197 45475 15255 45481
rect 15197 45472 15209 45475
rect 14792 45444 15209 45472
rect 14792 45432 14798 45444
rect 15197 45441 15209 45444
rect 15243 45441 15255 45475
rect 15197 45435 15255 45441
rect 17402 45432 17408 45484
rect 17460 45472 17466 45484
rect 17497 45475 17555 45481
rect 17497 45472 17509 45475
rect 17460 45444 17509 45472
rect 17460 45432 17466 45444
rect 17497 45441 17509 45444
rect 17543 45441 17555 45475
rect 17497 45435 17555 45441
rect 18322 45432 18328 45484
rect 18380 45472 18386 45484
rect 18785 45475 18843 45481
rect 18785 45472 18797 45475
rect 18380 45444 18797 45472
rect 18380 45432 18386 45444
rect 18785 45441 18797 45444
rect 18831 45441 18843 45475
rect 18785 45435 18843 45441
rect 23753 45475 23811 45481
rect 23753 45441 23765 45475
rect 23799 45472 23811 45475
rect 24026 45472 24032 45484
rect 23799 45444 24032 45472
rect 23799 45441 23811 45444
rect 23753 45435 23811 45441
rect 24026 45432 24032 45444
rect 24084 45432 24090 45484
rect 9033 45407 9091 45413
rect 9033 45373 9045 45407
rect 9079 45373 9091 45407
rect 9033 45367 9091 45373
rect 11149 45407 11207 45413
rect 11149 45373 11161 45407
rect 11195 45404 11207 45407
rect 11238 45404 11244 45416
rect 11195 45376 11244 45404
rect 11195 45373 11207 45376
rect 11149 45367 11207 45373
rect 6457 45271 6515 45277
rect 6457 45237 6469 45271
rect 6503 45268 6515 45271
rect 6546 45268 6552 45280
rect 6503 45240 6552 45268
rect 6503 45237 6515 45240
rect 6457 45231 6515 45237
rect 6546 45228 6552 45240
rect 6604 45228 6610 45280
rect 9048 45268 9076 45367
rect 11238 45364 11244 45376
rect 11296 45364 11302 45416
rect 13814 45364 13820 45416
rect 13872 45364 13878 45416
rect 13909 45407 13967 45413
rect 13909 45373 13921 45407
rect 13955 45373 13967 45407
rect 13909 45367 13967 45373
rect 20993 45407 21051 45413
rect 20993 45373 21005 45407
rect 21039 45404 21051 45407
rect 21174 45404 21180 45416
rect 21039 45376 21180 45404
rect 21039 45373 21051 45376
rect 20993 45367 21051 45373
rect 10318 45296 10324 45348
rect 10376 45336 10382 45348
rect 10781 45339 10839 45345
rect 10781 45336 10793 45339
rect 10376 45308 10793 45336
rect 10376 45296 10382 45308
rect 10781 45305 10793 45308
rect 10827 45336 10839 45339
rect 12158 45336 12164 45348
rect 10827 45308 12164 45336
rect 10827 45305 10839 45308
rect 10781 45299 10839 45305
rect 12158 45296 12164 45308
rect 12216 45296 12222 45348
rect 13357 45339 13415 45345
rect 13357 45305 13369 45339
rect 13403 45336 13415 45339
rect 13538 45336 13544 45348
rect 13403 45308 13544 45336
rect 13403 45305 13415 45308
rect 13357 45299 13415 45305
rect 13538 45296 13544 45308
rect 13596 45296 13602 45348
rect 13630 45296 13636 45348
rect 13688 45336 13694 45348
rect 13924 45336 13952 45367
rect 21174 45364 21180 45376
rect 21232 45364 21238 45416
rect 24213 45407 24271 45413
rect 24213 45373 24225 45407
rect 24259 45404 24271 45407
rect 24486 45404 24492 45416
rect 24259 45376 24492 45404
rect 24259 45373 24271 45376
rect 24213 45367 24271 45373
rect 24486 45364 24492 45376
rect 24544 45364 24550 45416
rect 24762 45364 24768 45416
rect 24820 45364 24826 45416
rect 13688 45308 13952 45336
rect 13688 45296 13694 45308
rect 10042 45268 10048 45280
rect 9048 45240 10048 45268
rect 10042 45228 10048 45240
rect 10100 45228 10106 45280
rect 12250 45228 12256 45280
rect 12308 45228 12314 45280
rect 15378 45228 15384 45280
rect 15436 45268 15442 45280
rect 15562 45268 15568 45280
rect 15436 45240 15568 45268
rect 15436 45228 15442 45240
rect 15562 45228 15568 45240
rect 15620 45228 15626 45280
rect 19150 45228 19156 45280
rect 19208 45268 19214 45280
rect 19245 45271 19303 45277
rect 19245 45268 19257 45271
rect 19208 45240 19257 45268
rect 19208 45228 19214 45240
rect 19245 45237 19257 45240
rect 19291 45237 19303 45271
rect 19245 45231 19303 45237
rect 21910 45228 21916 45280
rect 21968 45268 21974 45280
rect 22005 45271 22063 45277
rect 22005 45268 22017 45271
rect 21968 45240 22017 45268
rect 21968 45228 21974 45240
rect 22005 45237 22017 45240
rect 22051 45237 22063 45271
rect 22005 45231 22063 45237
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 6086 45024 6092 45076
rect 6144 45024 6150 45076
rect 6638 45024 6644 45076
rect 6696 45024 6702 45076
rect 7834 45024 7840 45076
rect 7892 45064 7898 45076
rect 8205 45067 8263 45073
rect 8205 45064 8217 45067
rect 7892 45036 8217 45064
rect 7892 45024 7898 45036
rect 8205 45033 8217 45036
rect 8251 45033 8263 45067
rect 8205 45027 8263 45033
rect 8662 45024 8668 45076
rect 8720 45064 8726 45076
rect 10413 45067 10471 45073
rect 10413 45064 10425 45067
rect 8720 45036 10425 45064
rect 8720 45024 8726 45036
rect 10413 45033 10425 45036
rect 10459 45033 10471 45067
rect 10413 45027 10471 45033
rect 12066 45024 12072 45076
rect 12124 45024 12130 45076
rect 16574 45024 16580 45076
rect 16632 45064 16638 45076
rect 19429 45067 19487 45073
rect 16632 45036 16804 45064
rect 16632 45024 16638 45036
rect 7282 44956 7288 45008
rect 7340 44956 7346 45008
rect 8846 44956 8852 45008
rect 8904 44996 8910 45008
rect 9125 44999 9183 45005
rect 9125 44996 9137 44999
rect 8904 44968 9137 44996
rect 8904 44956 8910 44968
rect 9125 44965 9137 44968
rect 9171 44965 9183 44999
rect 9125 44959 9183 44965
rect 10870 44956 10876 45008
rect 10928 44996 10934 45008
rect 11057 44999 11115 45005
rect 11057 44996 11069 44999
rect 10928 44968 11069 44996
rect 10928 44956 10934 44968
rect 11057 44965 11069 44968
rect 11103 44965 11115 44999
rect 11057 44959 11115 44965
rect 5902 44820 5908 44872
rect 5960 44820 5966 44872
rect 7650 44820 7656 44872
rect 7708 44860 7714 44872
rect 8021 44863 8079 44869
rect 8021 44860 8033 44863
rect 7708 44832 8033 44860
rect 7708 44820 7714 44832
rect 8021 44829 8033 44832
rect 8067 44829 8079 44863
rect 8021 44823 8079 44829
rect 12526 44820 12532 44872
rect 12584 44860 12590 44872
rect 13357 44863 13415 44869
rect 13357 44860 13369 44863
rect 12584 44832 13369 44860
rect 12584 44820 12590 44832
rect 13357 44829 13369 44832
rect 13403 44860 13415 44863
rect 13630 44860 13636 44872
rect 13403 44832 13636 44860
rect 13403 44829 13415 44832
rect 13357 44823 13415 44829
rect 13630 44820 13636 44832
rect 13688 44820 13694 44872
rect 15289 44863 15347 44869
rect 15289 44829 15301 44863
rect 15335 44829 15347 44863
rect 15289 44823 15347 44829
rect 6638 44752 6644 44804
rect 6696 44792 6702 44804
rect 6733 44795 6791 44801
rect 6733 44792 6745 44795
rect 6696 44764 6745 44792
rect 6696 44752 6702 44764
rect 6733 44761 6745 44764
rect 6779 44761 6791 44795
rect 6733 44755 6791 44761
rect 7282 44752 7288 44804
rect 7340 44792 7346 44804
rect 7469 44795 7527 44801
rect 7469 44792 7481 44795
rect 7340 44764 7481 44792
rect 7340 44752 7346 44764
rect 7469 44761 7481 44764
rect 7515 44761 7527 44795
rect 7469 44755 7527 44761
rect 8478 44752 8484 44804
rect 8536 44792 8542 44804
rect 9309 44795 9367 44801
rect 9309 44792 9321 44795
rect 8536 44764 9321 44792
rect 8536 44752 8542 44764
rect 9309 44761 9321 44764
rect 9355 44792 9367 44795
rect 9677 44795 9735 44801
rect 9677 44792 9689 44795
rect 9355 44764 9689 44792
rect 9355 44761 9367 44764
rect 9309 44755 9367 44761
rect 9677 44761 9689 44764
rect 9723 44761 9735 44795
rect 9677 44755 9735 44761
rect 10045 44795 10103 44801
rect 10045 44761 10057 44795
rect 10091 44792 10103 44795
rect 10502 44792 10508 44804
rect 10091 44764 10508 44792
rect 10091 44761 10103 44764
rect 10045 44755 10103 44761
rect 10502 44752 10508 44764
rect 10560 44752 10566 44804
rect 11238 44752 11244 44804
rect 11296 44752 11302 44804
rect 11701 44795 11759 44801
rect 11701 44761 11713 44795
rect 11747 44792 11759 44795
rect 12161 44795 12219 44801
rect 12161 44792 12173 44795
rect 11747 44764 12173 44792
rect 11747 44761 11759 44764
rect 11701 44755 11759 44761
rect 12161 44761 12173 44764
rect 12207 44792 12219 44795
rect 14274 44792 14280 44804
rect 12207 44764 14280 44792
rect 12207 44761 12219 44764
rect 12161 44755 12219 44761
rect 14274 44752 14280 44764
rect 14332 44752 14338 44804
rect 12713 44727 12771 44733
rect 12713 44693 12725 44727
rect 12759 44724 12771 44727
rect 12802 44724 12808 44736
rect 12759 44696 12808 44724
rect 12759 44693 12771 44696
rect 12713 44687 12771 44693
rect 12802 44684 12808 44696
rect 12860 44684 12866 44736
rect 15304 44724 15332 44823
rect 15562 44752 15568 44804
rect 15620 44752 15626 44804
rect 16776 44792 16804 45036
rect 19429 45033 19441 45067
rect 19475 45064 19487 45067
rect 20162 45064 20168 45076
rect 19475 45036 20168 45064
rect 19475 45033 19487 45036
rect 19429 45027 19487 45033
rect 20162 45024 20168 45036
rect 20220 45024 20226 45076
rect 24946 45024 24952 45076
rect 25004 45064 25010 45076
rect 25225 45067 25283 45073
rect 25225 45064 25237 45067
rect 25004 45036 25237 45064
rect 25004 45024 25010 45036
rect 25225 45033 25237 45036
rect 25271 45033 25283 45067
rect 25225 45027 25283 45033
rect 18233 44999 18291 45005
rect 18233 44965 18245 44999
rect 18279 44996 18291 44999
rect 19518 44996 19524 45008
rect 18279 44968 19524 44996
rect 18279 44965 18291 44968
rect 18233 44959 18291 44965
rect 19518 44956 19524 44968
rect 19576 44956 19582 45008
rect 22189 44931 22247 44937
rect 22189 44897 22201 44931
rect 22235 44928 22247 44931
rect 24026 44928 24032 44940
rect 22235 44900 24032 44928
rect 22235 44897 22247 44900
rect 22189 44891 22247 44897
rect 18874 44820 18880 44872
rect 18932 44820 18938 44872
rect 21174 44820 21180 44872
rect 21232 44860 21238 44872
rect 22002 44860 22008 44872
rect 21232 44832 22008 44860
rect 21232 44820 21238 44832
rect 22002 44820 22008 44832
rect 22060 44860 22066 44872
rect 22204 44860 22232 44891
rect 24026 44888 24032 44900
rect 24084 44888 24090 44940
rect 24581 44863 24639 44869
rect 24581 44860 24593 44863
rect 22060 44832 22232 44860
rect 23952 44832 24593 44860
rect 22060 44820 22066 44832
rect 17586 44792 17592 44804
rect 16776 44778 17592 44792
rect 16790 44764 17592 44778
rect 17586 44752 17592 44764
rect 17644 44752 17650 44804
rect 20622 44792 20628 44804
rect 20470 44764 20628 44792
rect 20622 44752 20628 44764
rect 20680 44752 20686 44804
rect 20901 44795 20959 44801
rect 20901 44761 20913 44795
rect 20947 44792 20959 44795
rect 21358 44792 21364 44804
rect 20947 44764 21364 44792
rect 20947 44761 20959 44764
rect 20901 44755 20959 44761
rect 21358 44752 21364 44764
rect 21416 44752 21422 44804
rect 21542 44752 21548 44804
rect 21600 44792 21606 44804
rect 22465 44795 22523 44801
rect 22465 44792 22477 44795
rect 21600 44764 22477 44792
rect 21600 44752 21606 44764
rect 22465 44761 22477 44764
rect 22511 44761 22523 44795
rect 22465 44755 22523 44761
rect 23474 44752 23480 44804
rect 23532 44752 23538 44804
rect 16206 44724 16212 44736
rect 15304 44696 16212 44724
rect 16206 44684 16212 44696
rect 16264 44724 16270 44736
rect 16482 44724 16488 44736
rect 16264 44696 16488 44724
rect 16264 44684 16270 44696
rect 16482 44684 16488 44696
rect 16540 44684 16546 44736
rect 17034 44684 17040 44736
rect 17092 44684 17098 44736
rect 21266 44684 21272 44736
rect 21324 44724 21330 44736
rect 21818 44724 21824 44736
rect 21324 44696 21824 44724
rect 21324 44684 21330 44696
rect 21818 44684 21824 44696
rect 21876 44684 21882 44736
rect 22738 44684 22744 44736
rect 22796 44724 22802 44736
rect 23952 44733 23980 44832
rect 24581 44829 24593 44832
rect 24627 44829 24639 44863
rect 24581 44823 24639 44829
rect 23937 44727 23995 44733
rect 23937 44724 23949 44727
rect 22796 44696 23949 44724
rect 22796 44684 22802 44696
rect 23937 44693 23949 44696
rect 23983 44693 23995 44727
rect 23937 44687 23995 44693
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 5994 44480 6000 44532
rect 6052 44520 6058 44532
rect 9125 44523 9183 44529
rect 9125 44520 9137 44523
rect 6052 44492 9137 44520
rect 6052 44480 6058 44492
rect 9125 44489 9137 44492
rect 9171 44489 9183 44523
rect 9125 44483 9183 44489
rect 9490 44480 9496 44532
rect 9548 44520 9554 44532
rect 9677 44523 9735 44529
rect 9677 44520 9689 44523
rect 9548 44492 9689 44520
rect 9548 44480 9554 44492
rect 9677 44489 9689 44492
rect 9723 44489 9735 44523
rect 9677 44483 9735 44489
rect 11882 44480 11888 44532
rect 11940 44480 11946 44532
rect 12253 44523 12311 44529
rect 12253 44489 12265 44523
rect 12299 44520 12311 44523
rect 14366 44520 14372 44532
rect 12299 44492 14372 44520
rect 12299 44489 12311 44492
rect 12253 44483 12311 44489
rect 14366 44480 14372 44492
rect 14424 44480 14430 44532
rect 21358 44480 21364 44532
rect 21416 44480 21422 44532
rect 21818 44480 21824 44532
rect 21876 44520 21882 44532
rect 22465 44523 22523 44529
rect 22465 44520 22477 44523
rect 21876 44492 22477 44520
rect 21876 44480 21882 44492
rect 22465 44489 22477 44492
rect 22511 44489 22523 44523
rect 22465 44483 22523 44489
rect 22557 44523 22615 44529
rect 22557 44489 22569 44523
rect 22603 44520 22615 44523
rect 23290 44520 23296 44532
rect 22603 44492 23296 44520
rect 22603 44489 22615 44492
rect 22557 44483 22615 44489
rect 23290 44480 23296 44492
rect 23348 44480 23354 44532
rect 6454 44412 6460 44464
rect 6512 44452 6518 44464
rect 6549 44455 6607 44461
rect 6549 44452 6561 44455
rect 6512 44424 6561 44452
rect 6512 44412 6518 44424
rect 6549 44421 6561 44424
rect 6595 44421 6607 44455
rect 6549 44415 6607 44421
rect 8386 44412 8392 44464
rect 8444 44452 8450 44464
rect 10873 44455 10931 44461
rect 10873 44452 10885 44455
rect 8444 44424 10885 44452
rect 8444 44412 8450 44424
rect 10873 44421 10885 44424
rect 10919 44421 10931 44455
rect 10873 44415 10931 44421
rect 17586 44412 17592 44464
rect 17644 44412 17650 44464
rect 21910 44412 21916 44464
rect 21968 44452 21974 44464
rect 21968 44424 22094 44452
rect 21968 44412 21974 44424
rect 6181 44387 6239 44393
rect 6181 44353 6193 44387
rect 6227 44384 6239 44387
rect 6733 44387 6791 44393
rect 6733 44384 6745 44387
rect 6227 44356 6745 44384
rect 6227 44353 6239 44356
rect 6181 44347 6239 44353
rect 6733 44353 6745 44356
rect 6779 44384 6791 44387
rect 6822 44384 6828 44396
rect 6779 44356 6828 44384
rect 6779 44353 6791 44356
rect 6733 44347 6791 44353
rect 6822 44344 6828 44356
rect 6880 44344 6886 44396
rect 8757 44387 8815 44393
rect 8757 44353 8769 44387
rect 8803 44384 8815 44387
rect 9214 44384 9220 44396
rect 8803 44356 9220 44384
rect 8803 44353 8815 44356
rect 8757 44347 8815 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 11057 44387 11115 44393
rect 11057 44353 11069 44387
rect 11103 44384 11115 44387
rect 11103 44356 11652 44384
rect 11103 44353 11115 44356
rect 11057 44347 11115 44353
rect 11624 44260 11652 44356
rect 14550 44344 14556 44396
rect 14608 44344 14614 44396
rect 14918 44344 14924 44396
rect 14976 44384 14982 44396
rect 16025 44387 16083 44393
rect 16025 44384 16037 44387
rect 14976 44356 16037 44384
rect 14976 44344 14982 44356
rect 16025 44353 16037 44356
rect 16071 44384 16083 44387
rect 16666 44384 16672 44396
rect 16071 44356 16672 44384
rect 16071 44353 16083 44356
rect 16025 44347 16083 44353
rect 16666 44344 16672 44356
rect 16724 44344 16730 44396
rect 19061 44387 19119 44393
rect 19061 44353 19073 44387
rect 19107 44384 19119 44387
rect 19150 44384 19156 44396
rect 19107 44356 19156 44384
rect 19107 44353 19119 44356
rect 19061 44347 19119 44353
rect 19150 44344 19156 44356
rect 19208 44344 19214 44396
rect 20162 44344 20168 44396
rect 20220 44384 20226 44396
rect 20717 44387 20775 44393
rect 20717 44384 20729 44387
rect 20220 44356 20729 44384
rect 20220 44344 20226 44356
rect 20717 44353 20729 44356
rect 20763 44353 20775 44387
rect 22066 44384 22094 44424
rect 23293 44387 23351 44393
rect 23293 44384 23305 44387
rect 22066 44356 23305 44384
rect 20717 44347 20775 44353
rect 23293 44353 23305 44356
rect 23339 44353 23351 44387
rect 23293 44347 23351 44353
rect 12342 44276 12348 44328
rect 12400 44276 12406 44328
rect 12437 44319 12495 44325
rect 12437 44285 12449 44319
rect 12483 44285 12495 44319
rect 12437 44279 12495 44285
rect 11606 44208 11612 44260
rect 11664 44208 11670 44260
rect 12250 44208 12256 44260
rect 12308 44248 12314 44260
rect 12452 44248 12480 44279
rect 12710 44276 12716 44328
rect 12768 44316 12774 44328
rect 13173 44319 13231 44325
rect 13173 44316 13185 44319
rect 12768 44288 13185 44316
rect 12768 44276 12774 44288
rect 13173 44285 13185 44288
rect 13219 44285 13231 44319
rect 13173 44279 13231 44285
rect 13446 44276 13452 44328
rect 13504 44276 13510 44328
rect 14568 44316 14596 44344
rect 16301 44319 16359 44325
rect 16301 44316 16313 44319
rect 14568 44288 16313 44316
rect 16301 44285 16313 44288
rect 16347 44285 16359 44319
rect 16301 44279 16359 44285
rect 16482 44276 16488 44328
rect 16540 44316 16546 44328
rect 16853 44319 16911 44325
rect 16853 44316 16865 44319
rect 16540 44288 16865 44316
rect 16540 44276 16546 44288
rect 16853 44285 16865 44288
rect 16899 44285 16911 44319
rect 16853 44279 16911 44285
rect 17126 44276 17132 44328
rect 17184 44316 17190 44328
rect 17770 44316 17776 44328
rect 17184 44288 17776 44316
rect 17184 44276 17190 44288
rect 17770 44276 17776 44288
rect 17828 44276 17834 44328
rect 22741 44319 22799 44325
rect 22741 44285 22753 44319
rect 22787 44316 22799 44319
rect 23566 44316 23572 44328
rect 22787 44288 23572 44316
rect 22787 44285 22799 44288
rect 22741 44279 22799 44285
rect 23566 44276 23572 44288
rect 23624 44276 23630 44328
rect 24489 44319 24547 44325
rect 24489 44285 24501 44319
rect 24535 44316 24547 44319
rect 24670 44316 24676 44328
rect 24535 44288 24676 44316
rect 24535 44285 24547 44288
rect 24489 44279 24547 44285
rect 24670 44276 24676 44288
rect 24728 44276 24734 44328
rect 24762 44276 24768 44328
rect 24820 44276 24826 44328
rect 12308 44220 12480 44248
rect 12308 44208 12314 44220
rect 7193 44183 7251 44189
rect 7193 44149 7205 44183
rect 7239 44180 7251 44183
rect 7282 44180 7288 44192
rect 7239 44152 7288 44180
rect 7239 44149 7251 44152
rect 7193 44143 7251 44149
rect 7282 44140 7288 44152
rect 7340 44140 7346 44192
rect 14734 44140 14740 44192
rect 14792 44180 14798 44192
rect 14921 44183 14979 44189
rect 14921 44180 14933 44183
rect 14792 44152 14933 44180
rect 14792 44140 14798 44152
rect 14921 44149 14933 44152
rect 14967 44149 14979 44183
rect 14921 44143 14979 44149
rect 15194 44140 15200 44192
rect 15252 44180 15258 44192
rect 15381 44183 15439 44189
rect 15381 44180 15393 44183
rect 15252 44152 15393 44180
rect 15252 44140 15258 44152
rect 15381 44149 15393 44152
rect 15427 44149 15439 44183
rect 15381 44143 15439 44149
rect 18322 44140 18328 44192
rect 18380 44180 18386 44192
rect 18601 44183 18659 44189
rect 18601 44180 18613 44183
rect 18380 44152 18613 44180
rect 18380 44140 18386 44152
rect 18601 44149 18613 44152
rect 18647 44149 18659 44183
rect 18601 44143 18659 44149
rect 19610 44140 19616 44192
rect 19668 44180 19674 44192
rect 19705 44183 19763 44189
rect 19705 44180 19717 44183
rect 19668 44152 19717 44180
rect 19668 44140 19674 44152
rect 19705 44149 19717 44152
rect 19751 44149 19763 44183
rect 19705 44143 19763 44149
rect 22094 44140 22100 44192
rect 22152 44140 22158 44192
rect 22830 44140 22836 44192
rect 22888 44180 22894 44192
rect 23937 44183 23995 44189
rect 23937 44180 23949 44183
rect 22888 44152 23949 44180
rect 22888 44140 22894 44152
rect 23937 44149 23949 44152
rect 23983 44149 23995 44183
rect 23937 44143 23995 44149
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 7558 43936 7564 43988
rect 7616 43976 7622 43988
rect 8021 43979 8079 43985
rect 8021 43976 8033 43979
rect 7616 43948 8033 43976
rect 7616 43936 7622 43948
rect 8021 43945 8033 43948
rect 8067 43945 8079 43979
rect 8021 43939 8079 43945
rect 8573 43979 8631 43985
rect 8573 43945 8585 43979
rect 8619 43976 8631 43979
rect 9398 43976 9404 43988
rect 8619 43948 9404 43976
rect 8619 43945 8631 43948
rect 8573 43939 8631 43945
rect 8036 43704 8064 43939
rect 9398 43936 9404 43948
rect 9456 43936 9462 43988
rect 9953 43979 10011 43985
rect 9953 43945 9965 43979
rect 9999 43976 10011 43979
rect 12342 43976 12348 43988
rect 9999 43948 12348 43976
rect 9999 43945 10011 43948
rect 9953 43939 10011 43945
rect 12342 43936 12348 43948
rect 12400 43936 12406 43988
rect 13814 43936 13820 43988
rect 13872 43976 13878 43988
rect 15381 43979 15439 43985
rect 15381 43976 15393 43979
rect 13872 43948 15393 43976
rect 13872 43936 13878 43948
rect 15381 43945 15393 43948
rect 15427 43945 15439 43979
rect 15381 43939 15439 43945
rect 15562 43936 15568 43988
rect 15620 43976 15626 43988
rect 15620 43948 17816 43976
rect 15620 43936 15626 43948
rect 10229 43911 10287 43917
rect 10229 43908 10241 43911
rect 9324 43880 10241 43908
rect 9324 43852 9352 43880
rect 10229 43877 10241 43880
rect 10275 43877 10287 43911
rect 10229 43871 10287 43877
rect 9306 43800 9312 43852
rect 9364 43800 9370 43852
rect 9490 43800 9496 43852
rect 9548 43800 9554 43852
rect 10244 43840 10272 43871
rect 10962 43868 10968 43920
rect 11020 43908 11026 43920
rect 11977 43911 12035 43917
rect 11977 43908 11989 43911
rect 11020 43880 11989 43908
rect 11020 43868 11026 43880
rect 11977 43877 11989 43880
rect 12023 43877 12035 43911
rect 16114 43908 16120 43920
rect 11977 43871 12035 43877
rect 12406 43880 16120 43908
rect 12406 43840 12434 43880
rect 16114 43868 16120 43880
rect 16172 43868 16178 43920
rect 10244 43812 12434 43840
rect 12618 43800 12624 43852
rect 12676 43840 12682 43852
rect 12676 43812 14320 43840
rect 12676 43800 12682 43812
rect 8389 43775 8447 43781
rect 8389 43741 8401 43775
rect 8435 43772 8447 43775
rect 10226 43772 10232 43784
rect 8435 43744 10232 43772
rect 8435 43741 8447 43744
rect 8389 43735 8447 43741
rect 10226 43732 10232 43744
rect 10284 43732 10290 43784
rect 14292 43781 14320 43812
rect 14734 43800 14740 43852
rect 14792 43840 14798 43852
rect 15933 43843 15991 43849
rect 15933 43840 15945 43843
rect 14792 43812 15945 43840
rect 14792 43800 14798 43812
rect 15933 43809 15945 43812
rect 15979 43809 15991 43843
rect 15933 43803 15991 43809
rect 17678 43800 17684 43852
rect 17736 43800 17742 43852
rect 17788 43849 17816 43948
rect 22646 43936 22652 43988
rect 22704 43976 22710 43988
rect 22704 43948 22968 43976
rect 22704 43936 22710 43948
rect 19334 43908 19340 43920
rect 18432 43880 19340 43908
rect 17773 43843 17831 43849
rect 17773 43809 17785 43843
rect 17819 43809 17831 43843
rect 17773 43803 17831 43809
rect 14277 43775 14335 43781
rect 14277 43741 14289 43775
rect 14323 43741 14335 43775
rect 14277 43735 14335 43741
rect 15749 43775 15807 43781
rect 15749 43741 15761 43775
rect 15795 43772 15807 43775
rect 18432 43772 18460 43880
rect 19334 43868 19340 43880
rect 19392 43868 19398 43920
rect 22830 43908 22836 43920
rect 21928 43880 22836 43908
rect 18509 43843 18567 43849
rect 18509 43809 18521 43843
rect 18555 43840 18567 43843
rect 21082 43840 21088 43852
rect 18555 43812 21088 43840
rect 18555 43809 18567 43812
rect 18509 43803 18567 43809
rect 15795 43744 18460 43772
rect 15795 43741 15807 43744
rect 15749 43735 15807 43741
rect 9585 43707 9643 43713
rect 9585 43704 9597 43707
rect 8036 43676 9597 43704
rect 9585 43673 9597 43676
rect 9631 43704 9643 43707
rect 10778 43704 10784 43716
rect 9631 43676 10784 43704
rect 9631 43673 9643 43676
rect 9585 43667 9643 43673
rect 10778 43664 10784 43676
rect 10836 43664 10842 43716
rect 12437 43707 12495 43713
rect 12437 43673 12449 43707
rect 12483 43704 12495 43707
rect 16850 43704 16856 43716
rect 12483 43676 16856 43704
rect 12483 43673 12495 43676
rect 12437 43667 12495 43673
rect 16850 43664 16856 43676
rect 16908 43664 16914 43716
rect 17589 43707 17647 43713
rect 17589 43673 17601 43707
rect 17635 43704 17647 43707
rect 18524 43704 18552 43803
rect 21082 43800 21088 43812
rect 21140 43800 21146 43852
rect 21177 43843 21235 43849
rect 21177 43809 21189 43843
rect 21223 43840 21235 43843
rect 21928 43840 21956 43880
rect 22830 43868 22836 43880
rect 22888 43868 22894 43920
rect 22940 43908 22968 43948
rect 23474 43936 23480 43988
rect 23532 43936 23538 43988
rect 25682 43908 25688 43920
rect 22940 43880 25688 43908
rect 25682 43868 25688 43880
rect 25740 43868 25746 43920
rect 21223 43812 21956 43840
rect 22097 43843 22155 43849
rect 21223 43809 21235 43812
rect 21177 43803 21235 43809
rect 22097 43809 22109 43843
rect 22143 43840 22155 43843
rect 22738 43840 22744 43852
rect 22143 43812 22744 43840
rect 22143 43809 22155 43812
rect 22097 43803 22155 43809
rect 22738 43800 22744 43812
rect 22796 43800 22802 43852
rect 23109 43843 23167 43849
rect 23109 43809 23121 43843
rect 23155 43840 23167 43843
rect 24670 43840 24676 43852
rect 23155 43812 24676 43840
rect 23155 43809 23167 43812
rect 23109 43803 23167 43809
rect 24670 43800 24676 43812
rect 24728 43800 24734 43852
rect 21453 43775 21511 43781
rect 21453 43741 21465 43775
rect 21499 43772 21511 43775
rect 21499 43744 22048 43772
rect 21499 43741 21511 43744
rect 21453 43735 21511 43741
rect 22020 43716 22048 43744
rect 22186 43732 22192 43784
rect 22244 43772 22250 43784
rect 22281 43775 22339 43781
rect 22281 43772 22293 43775
rect 22244 43744 22293 43772
rect 22244 43732 22250 43744
rect 22281 43741 22293 43744
rect 22327 43741 22339 43775
rect 22281 43735 22339 43741
rect 24026 43732 24032 43784
rect 24084 43772 24090 43784
rect 24581 43775 24639 43781
rect 24581 43772 24593 43775
rect 24084 43744 24593 43772
rect 24084 43732 24090 43744
rect 24581 43741 24593 43744
rect 24627 43741 24639 43775
rect 24581 43735 24639 43741
rect 17635 43676 18552 43704
rect 19628 43676 19932 43704
rect 17635 43673 17647 43676
rect 17589 43667 17647 43673
rect 12342 43596 12348 43648
rect 12400 43596 12406 43648
rect 14918 43596 14924 43648
rect 14976 43596 14982 43648
rect 15838 43596 15844 43648
rect 15896 43596 15902 43648
rect 17218 43596 17224 43648
rect 17276 43596 17282 43648
rect 17770 43596 17776 43648
rect 17828 43636 17834 43648
rect 18233 43639 18291 43645
rect 18233 43636 18245 43639
rect 17828 43608 18245 43636
rect 17828 43596 17834 43608
rect 18233 43605 18245 43608
rect 18279 43636 18291 43639
rect 19628 43636 19656 43676
rect 18279 43608 19656 43636
rect 18279 43605 18291 43608
rect 18233 43599 18291 43605
rect 19702 43596 19708 43648
rect 19760 43596 19766 43648
rect 19904 43636 19932 43676
rect 20622 43664 20628 43716
rect 20680 43664 20686 43716
rect 22002 43664 22008 43716
rect 22060 43664 22066 43716
rect 23658 43664 23664 43716
rect 23716 43704 23722 43716
rect 23753 43707 23811 43713
rect 23753 43704 23765 43707
rect 23716 43676 23765 43704
rect 23716 43664 23722 43676
rect 23753 43673 23765 43676
rect 23799 43704 23811 43707
rect 24121 43707 24179 43713
rect 24121 43704 24133 43707
rect 23799 43676 24133 43704
rect 23799 43673 23811 43676
rect 23753 43667 23811 43673
rect 24121 43673 24133 43676
rect 24167 43673 24179 43707
rect 24121 43667 24179 43673
rect 21266 43636 21272 43648
rect 19904 43608 21272 43636
rect 21266 43596 21272 43608
rect 21324 43596 21330 43648
rect 22189 43639 22247 43645
rect 22189 43605 22201 43639
rect 22235 43636 22247 43639
rect 22462 43636 22468 43648
rect 22235 43608 22468 43636
rect 22235 43605 22247 43608
rect 22189 43599 22247 43605
rect 22462 43596 22468 43608
rect 22520 43596 22526 43648
rect 22646 43596 22652 43648
rect 22704 43596 22710 43648
rect 23474 43596 23480 43648
rect 23532 43636 23538 43648
rect 24578 43636 24584 43648
rect 23532 43608 24584 43636
rect 23532 43596 23538 43608
rect 24578 43596 24584 43608
rect 24636 43596 24642 43648
rect 24946 43596 24952 43648
rect 25004 43636 25010 43648
rect 25225 43639 25283 43645
rect 25225 43636 25237 43639
rect 25004 43608 25237 43636
rect 25004 43596 25010 43608
rect 25225 43605 25237 43608
rect 25271 43605 25283 43639
rect 25225 43599 25283 43605
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 7742 43392 7748 43444
rect 7800 43432 7806 43444
rect 8113 43435 8171 43441
rect 8113 43432 8125 43435
rect 7800 43404 8125 43432
rect 7800 43392 7806 43404
rect 8113 43401 8125 43404
rect 8159 43401 8171 43435
rect 8113 43395 8171 43401
rect 12802 43392 12808 43444
rect 12860 43392 12866 43444
rect 15381 43435 15439 43441
rect 15381 43401 15393 43435
rect 15427 43432 15439 43435
rect 15470 43432 15476 43444
rect 15427 43404 15476 43432
rect 15427 43401 15439 43404
rect 15381 43395 15439 43401
rect 15470 43392 15476 43404
rect 15528 43392 15534 43444
rect 16574 43432 16580 43444
rect 16224 43404 16580 43432
rect 9398 43324 9404 43376
rect 9456 43324 9462 43376
rect 10042 43324 10048 43376
rect 10100 43364 10106 43376
rect 12820 43364 12848 43392
rect 12989 43367 13047 43373
rect 12989 43364 13001 43367
rect 10100 43336 10456 43364
rect 12820 43336 13001 43364
rect 10100 43324 10106 43336
rect 10428 43308 10456 43336
rect 12989 43333 13001 43336
rect 13035 43333 13047 43367
rect 12989 43327 13047 43333
rect 1302 43256 1308 43308
rect 1360 43296 1366 43308
rect 1673 43299 1731 43305
rect 1673 43296 1685 43299
rect 1360 43268 1685 43296
rect 1360 43256 1366 43268
rect 1673 43265 1685 43268
rect 1719 43296 1731 43299
rect 2133 43299 2191 43305
rect 2133 43296 2145 43299
rect 1719 43268 2145 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 2133 43265 2145 43268
rect 2179 43265 2191 43299
rect 2133 43259 2191 43265
rect 7834 43256 7840 43308
rect 7892 43296 7898 43308
rect 7929 43299 7987 43305
rect 7929 43296 7941 43299
rect 7892 43268 7941 43296
rect 7892 43256 7898 43268
rect 7929 43265 7941 43268
rect 7975 43265 7987 43299
rect 7929 43259 7987 43265
rect 10410 43256 10416 43308
rect 10468 43256 10474 43308
rect 14826 43296 14832 43308
rect 14122 43268 14832 43296
rect 14826 43256 14832 43268
rect 14884 43296 14890 43308
rect 16025 43299 16083 43305
rect 16025 43296 16037 43299
rect 14884 43268 16037 43296
rect 14884 43256 14890 43268
rect 16025 43265 16037 43268
rect 16071 43265 16083 43299
rect 16025 43259 16083 43265
rect 10137 43231 10195 43237
rect 10137 43197 10149 43231
rect 10183 43228 10195 43231
rect 11054 43228 11060 43240
rect 10183 43200 11060 43228
rect 10183 43197 10195 43200
rect 10137 43191 10195 43197
rect 11054 43188 11060 43200
rect 11112 43188 11118 43240
rect 11146 43188 11152 43240
rect 11204 43188 11210 43240
rect 12710 43188 12716 43240
rect 12768 43188 12774 43240
rect 15470 43188 15476 43240
rect 15528 43188 15534 43240
rect 15562 43188 15568 43240
rect 15620 43188 15626 43240
rect 1857 43163 1915 43169
rect 1857 43129 1869 43163
rect 1903 43160 1915 43163
rect 3786 43160 3792 43172
rect 1903 43132 3792 43160
rect 1903 43129 1915 43132
rect 1857 43123 1915 43129
rect 3786 43120 3792 43132
rect 3844 43120 3850 43172
rect 14461 43163 14519 43169
rect 14461 43129 14473 43163
rect 14507 43160 14519 43163
rect 15286 43160 15292 43172
rect 14507 43132 15292 43160
rect 14507 43129 14519 43132
rect 14461 43123 14519 43129
rect 15286 43120 15292 43132
rect 15344 43120 15350 43172
rect 15488 43160 15516 43188
rect 16224 43169 16252 43404
rect 16574 43392 16580 43404
rect 16632 43392 16638 43444
rect 17221 43435 17279 43441
rect 17221 43401 17233 43435
rect 17267 43432 17279 43435
rect 17494 43432 17500 43444
rect 17267 43404 17500 43432
rect 17267 43401 17279 43404
rect 17221 43395 17279 43401
rect 17494 43392 17500 43404
rect 17552 43392 17558 43444
rect 19426 43392 19432 43444
rect 19484 43392 19490 43444
rect 19702 43392 19708 43444
rect 19760 43432 19766 43444
rect 19760 43404 20392 43432
rect 19760 43392 19766 43404
rect 19444 43364 19472 43392
rect 19444 43336 19932 43364
rect 17313 43299 17371 43305
rect 17313 43265 17325 43299
rect 17359 43296 17371 43299
rect 17770 43296 17776 43308
rect 17359 43268 17776 43296
rect 17359 43265 17371 43268
rect 17313 43259 17371 43265
rect 17770 43256 17776 43268
rect 17828 43256 17834 43308
rect 19904 43305 19932 43336
rect 20364 43305 20392 43404
rect 22278 43392 22284 43444
rect 22336 43392 22342 43444
rect 22370 43392 22376 43444
rect 22428 43432 22434 43444
rect 22428 43404 22508 43432
rect 22428 43392 22434 43404
rect 19889 43299 19947 43305
rect 17126 43188 17132 43240
rect 17184 43188 17190 43240
rect 17862 43188 17868 43240
rect 17920 43228 17926 43240
rect 18524 43228 18552 43282
rect 19889 43265 19901 43299
rect 19935 43265 19947 43299
rect 19889 43259 19947 43265
rect 20349 43299 20407 43305
rect 20349 43265 20361 43299
rect 20395 43265 20407 43299
rect 20349 43259 20407 43265
rect 21358 43256 21364 43308
rect 21416 43296 21422 43308
rect 21726 43296 21732 43308
rect 21416 43268 21732 43296
rect 21416 43256 21422 43268
rect 21726 43256 21732 43268
rect 21784 43296 21790 43308
rect 22373 43299 22431 43305
rect 22373 43296 22385 43299
rect 21784 43268 22385 43296
rect 21784 43256 21790 43268
rect 22373 43265 22385 43268
rect 22419 43265 22431 43299
rect 22373 43259 22431 43265
rect 22480 43240 22508 43404
rect 23382 43392 23388 43444
rect 23440 43432 23446 43444
rect 23440 43404 23888 43432
rect 23440 43392 23446 43404
rect 23860 43308 23888 43404
rect 24946 43324 24952 43376
rect 25004 43324 25010 43376
rect 23842 43256 23848 43308
rect 23900 43256 23906 43308
rect 19518 43228 19524 43240
rect 17920 43200 19524 43228
rect 17920 43188 17926 43200
rect 19518 43188 19524 43200
rect 19576 43188 19582 43240
rect 19610 43188 19616 43240
rect 19668 43188 19674 43240
rect 22189 43231 22247 43237
rect 22189 43197 22201 43231
rect 22235 43197 22247 43231
rect 22189 43191 22247 43197
rect 16209 43163 16267 43169
rect 16209 43160 16221 43163
rect 15488 43132 16221 43160
rect 16209 43129 16221 43132
rect 16255 43129 16267 43163
rect 16209 43123 16267 43129
rect 17681 43163 17739 43169
rect 17681 43129 17693 43163
rect 17727 43160 17739 43163
rect 18414 43160 18420 43172
rect 17727 43132 18420 43160
rect 17727 43129 17739 43132
rect 17681 43123 17739 43129
rect 18414 43120 18420 43132
rect 18472 43120 18478 43172
rect 22204 43160 22232 43191
rect 22462 43188 22468 43240
rect 22520 43188 22526 43240
rect 25225 43231 25283 43237
rect 22664 43200 25176 43228
rect 22370 43160 22376 43172
rect 22204 43132 22376 43160
rect 22370 43120 22376 43132
rect 22428 43120 22434 43172
rect 3510 43052 3516 43104
rect 3568 43092 3574 43104
rect 8662 43092 8668 43104
rect 3568 43064 8668 43092
rect 3568 43052 3574 43064
rect 8662 43052 8668 43064
rect 8720 43052 8726 43104
rect 12802 43052 12808 43104
rect 12860 43092 12866 43104
rect 13446 43092 13452 43104
rect 12860 43064 13452 43092
rect 12860 43052 12866 43064
rect 13446 43052 13452 43064
rect 13504 43052 13510 43104
rect 15013 43095 15071 43101
rect 15013 43061 15025 43095
rect 15059 43092 15071 43095
rect 15102 43092 15108 43104
rect 15059 43064 15108 43092
rect 15059 43061 15071 43064
rect 15013 43055 15071 43061
rect 15102 43052 15108 43064
rect 15160 43052 15166 43104
rect 18141 43095 18199 43101
rect 18141 43061 18153 43095
rect 18187 43092 18199 43095
rect 18874 43092 18880 43104
rect 18187 43064 18880 43092
rect 18187 43061 18199 43064
rect 18141 43055 18199 43061
rect 18874 43052 18880 43064
rect 18932 43052 18938 43104
rect 19518 43052 19524 43104
rect 19576 43092 19582 43104
rect 20622 43092 20628 43104
rect 19576 43064 20628 43092
rect 19576 43052 19582 43064
rect 20622 43052 20628 43064
rect 20680 43052 20686 43104
rect 20990 43052 20996 43104
rect 21048 43052 21054 43104
rect 21358 43052 21364 43104
rect 21416 43052 21422 43104
rect 21450 43052 21456 43104
rect 21508 43092 21514 43104
rect 21637 43095 21695 43101
rect 21637 43092 21649 43095
rect 21508 43064 21649 43092
rect 21508 43052 21514 43064
rect 21637 43061 21649 43064
rect 21683 43092 21695 43095
rect 22664 43092 22692 43200
rect 22741 43163 22799 43169
rect 22741 43129 22753 43163
rect 22787 43160 22799 43163
rect 23382 43160 23388 43172
rect 22787 43132 23388 43160
rect 22787 43129 22799 43132
rect 22741 43123 22799 43129
rect 23382 43120 23388 43132
rect 23440 43120 23446 43172
rect 25148 43160 25176 43200
rect 25225 43197 25237 43231
rect 25271 43228 25283 43231
rect 25314 43228 25320 43240
rect 25271 43200 25320 43228
rect 25271 43197 25283 43200
rect 25225 43191 25283 43197
rect 25314 43188 25320 43200
rect 25372 43188 25378 43240
rect 26050 43160 26056 43172
rect 25148 43132 26056 43160
rect 26050 43120 26056 43132
rect 26108 43120 26114 43172
rect 21683 43064 22692 43092
rect 23109 43095 23167 43101
rect 21683 43061 21695 43064
rect 21637 43055 21695 43061
rect 23109 43061 23121 43095
rect 23155 43092 23167 43095
rect 23290 43092 23296 43104
rect 23155 43064 23296 43092
rect 23155 43061 23167 43064
rect 23109 43055 23167 43061
rect 23290 43052 23296 43064
rect 23348 43052 23354 43104
rect 23477 43095 23535 43101
rect 23477 43061 23489 43095
rect 23523 43092 23535 43095
rect 23566 43092 23572 43104
rect 23523 43064 23572 43092
rect 23523 43061 23535 43064
rect 23477 43055 23535 43061
rect 23566 43052 23572 43064
rect 23624 43092 23630 43104
rect 24302 43092 24308 43104
rect 23624 43064 24308 43092
rect 23624 43052 23630 43064
rect 24302 43052 24308 43064
rect 24360 43052 24366 43104
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 14918 42848 14924 42900
rect 14976 42888 14982 42900
rect 15178 42891 15236 42897
rect 15178 42888 15190 42891
rect 14976 42860 15190 42888
rect 14976 42848 14982 42860
rect 15178 42857 15190 42860
rect 15224 42857 15236 42891
rect 15178 42851 15236 42857
rect 17494 42848 17500 42900
rect 17552 42888 17558 42900
rect 19702 42888 19708 42900
rect 17552 42860 19708 42888
rect 17552 42848 17558 42860
rect 19702 42848 19708 42860
rect 19760 42848 19766 42900
rect 22544 42891 22602 42897
rect 22544 42857 22556 42891
rect 22590 42888 22602 42891
rect 24581 42891 24639 42897
rect 24581 42888 24593 42891
rect 22590 42860 24593 42888
rect 22590 42857 22602 42860
rect 22544 42851 22602 42857
rect 24581 42857 24593 42860
rect 24627 42857 24639 42891
rect 24581 42851 24639 42857
rect 13446 42780 13452 42832
rect 13504 42820 13510 42832
rect 19610 42820 19616 42832
rect 13504 42792 15056 42820
rect 13504 42780 13510 42792
rect 4709 42755 4767 42761
rect 4709 42721 4721 42755
rect 4755 42752 4767 42755
rect 4798 42752 4804 42764
rect 4755 42724 4804 42752
rect 4755 42721 4767 42724
rect 4709 42715 4767 42721
rect 4798 42712 4804 42724
rect 4856 42712 4862 42764
rect 5442 42712 5448 42764
rect 5500 42752 5506 42764
rect 5721 42755 5779 42761
rect 5721 42752 5733 42755
rect 5500 42724 5733 42752
rect 5500 42712 5506 42724
rect 5721 42721 5733 42724
rect 5767 42721 5779 42755
rect 9677 42755 9735 42761
rect 9677 42752 9689 42755
rect 5721 42715 5779 42721
rect 8588 42724 9689 42752
rect 8588 42696 8616 42724
rect 9677 42721 9689 42724
rect 9723 42721 9735 42755
rect 9677 42715 9735 42721
rect 10410 42712 10416 42764
rect 10468 42752 10474 42764
rect 11057 42755 11115 42761
rect 11057 42752 11069 42755
rect 10468 42724 11069 42752
rect 10468 42712 10474 42724
rect 11057 42721 11069 42724
rect 11103 42721 11115 42755
rect 11057 42715 11115 42721
rect 12618 42712 12624 42764
rect 12676 42752 12682 42764
rect 12805 42755 12863 42761
rect 12805 42752 12817 42755
rect 12676 42724 12817 42752
rect 12676 42712 12682 42724
rect 12805 42721 12817 42724
rect 12851 42721 12863 42755
rect 15028 42752 15056 42792
rect 16224 42792 19616 42820
rect 16224 42752 16252 42792
rect 15028 42724 16252 42752
rect 16669 42755 16727 42761
rect 12805 42715 12863 42721
rect 16669 42721 16681 42755
rect 16715 42752 16727 42755
rect 17310 42752 17316 42764
rect 16715 42724 17316 42752
rect 16715 42721 16727 42724
rect 16669 42715 16727 42721
rect 17310 42712 17316 42724
rect 17368 42712 17374 42764
rect 17788 42761 17816 42792
rect 19610 42780 19616 42792
rect 19668 42780 19674 42832
rect 19720 42761 19748 42848
rect 21542 42820 21548 42832
rect 21192 42792 21548 42820
rect 17773 42755 17831 42761
rect 17773 42721 17785 42755
rect 17819 42721 17831 42755
rect 17773 42715 17831 42721
rect 19705 42755 19763 42761
rect 19705 42721 19717 42755
rect 19751 42721 19763 42755
rect 19705 42715 19763 42721
rect 19889 42755 19947 42761
rect 19889 42721 19901 42755
rect 19935 42752 19947 42755
rect 20254 42752 20260 42764
rect 19935 42724 20260 42752
rect 19935 42721 19947 42724
rect 19889 42715 19947 42721
rect 20254 42712 20260 42724
rect 20312 42712 20318 42764
rect 21192 42761 21220 42792
rect 21542 42780 21548 42792
rect 21600 42820 21606 42832
rect 21726 42820 21732 42832
rect 21600 42792 21732 42820
rect 21600 42780 21606 42792
rect 21726 42780 21732 42792
rect 21784 42780 21790 42832
rect 23566 42780 23572 42832
rect 23624 42820 23630 42832
rect 25774 42820 25780 42832
rect 23624 42792 25780 42820
rect 23624 42780 23630 42792
rect 25774 42780 25780 42792
rect 25832 42780 25838 42832
rect 21177 42755 21235 42761
rect 21177 42721 21189 42755
rect 21223 42721 21235 42755
rect 21177 42715 21235 42721
rect 21266 42712 21272 42764
rect 21324 42712 21330 42764
rect 22002 42712 22008 42764
rect 22060 42752 22066 42764
rect 22281 42755 22339 42761
rect 22281 42752 22293 42755
rect 22060 42724 22293 42752
rect 22060 42712 22066 42724
rect 22281 42721 22293 42724
rect 22327 42752 22339 42755
rect 25314 42752 25320 42764
rect 22327 42724 25320 42752
rect 22327 42721 22339 42724
rect 22281 42715 22339 42721
rect 25314 42712 25320 42724
rect 25372 42712 25378 42764
rect 8570 42644 8576 42696
rect 8628 42644 8634 42696
rect 14182 42644 14188 42696
rect 14240 42684 14246 42696
rect 14921 42687 14979 42693
rect 14921 42684 14933 42687
rect 14240 42656 14933 42684
rect 14240 42644 14246 42656
rect 14921 42653 14933 42656
rect 14967 42653 14979 42687
rect 14921 42647 14979 42653
rect 16758 42644 16764 42696
rect 16816 42684 16822 42696
rect 17589 42687 17647 42693
rect 17589 42684 17601 42687
rect 16816 42656 17601 42684
rect 16816 42644 16822 42656
rect 17589 42653 17601 42656
rect 17635 42684 17647 42687
rect 18325 42687 18383 42693
rect 18325 42684 18337 42687
rect 17635 42656 18337 42684
rect 17635 42653 17647 42656
rect 17589 42647 17647 42653
rect 18325 42653 18337 42656
rect 18371 42653 18383 42687
rect 18325 42647 18383 42653
rect 21361 42687 21419 42693
rect 21361 42653 21373 42687
rect 21407 42684 21419 42687
rect 21450 42684 21456 42696
rect 21407 42656 21456 42684
rect 21407 42653 21419 42656
rect 21361 42647 21419 42653
rect 21450 42644 21456 42656
rect 21508 42644 21514 42696
rect 24026 42644 24032 42696
rect 24084 42644 24090 42696
rect 25222 42644 25228 42696
rect 25280 42644 25286 42696
rect 4893 42619 4951 42625
rect 4893 42585 4905 42619
rect 4939 42585 4951 42619
rect 4893 42579 4951 42585
rect 5905 42619 5963 42625
rect 5905 42585 5917 42619
rect 5951 42585 5963 42619
rect 5905 42579 5963 42585
rect 10229 42619 10287 42625
rect 10229 42585 10241 42619
rect 10275 42616 10287 42619
rect 10505 42619 10563 42625
rect 10505 42616 10517 42619
rect 10275 42588 10517 42616
rect 10275 42585 10287 42588
rect 10229 42579 10287 42585
rect 10505 42585 10517 42588
rect 10551 42616 10563 42619
rect 11238 42616 11244 42628
rect 10551 42588 11244 42616
rect 10551 42585 10563 42588
rect 10505 42579 10563 42585
rect 4908 42548 4936 42579
rect 5258 42548 5264 42560
rect 4908 42520 5264 42548
rect 5258 42508 5264 42520
rect 5316 42508 5322 42560
rect 5920 42548 5948 42579
rect 11238 42576 11244 42588
rect 11296 42576 11302 42628
rect 11330 42576 11336 42628
rect 11388 42576 11394 42628
rect 12618 42616 12624 42628
rect 12558 42588 12624 42616
rect 12618 42576 12624 42588
rect 12676 42616 12682 42628
rect 12676 42588 13952 42616
rect 12676 42576 12682 42588
rect 6362 42548 6368 42560
rect 5920 42520 6368 42548
rect 6362 42508 6368 42520
rect 6420 42508 6426 42560
rect 7742 42508 7748 42560
rect 7800 42548 7806 42560
rect 7929 42551 7987 42557
rect 7929 42548 7941 42551
rect 7800 42520 7941 42548
rect 7800 42508 7806 42520
rect 7929 42517 7941 42520
rect 7975 42517 7987 42551
rect 7929 42511 7987 42517
rect 8938 42508 8944 42560
rect 8996 42548 9002 42560
rect 9125 42551 9183 42557
rect 9125 42548 9137 42551
rect 8996 42520 9137 42548
rect 8996 42508 9002 42520
rect 9125 42517 9137 42520
rect 9171 42517 9183 42551
rect 9125 42511 9183 42517
rect 9398 42508 9404 42560
rect 9456 42548 9462 42560
rect 9493 42551 9551 42557
rect 9493 42548 9505 42551
rect 9456 42520 9505 42548
rect 9456 42508 9462 42520
rect 9493 42517 9505 42520
rect 9539 42517 9551 42551
rect 9493 42511 9551 42517
rect 9582 42508 9588 42560
rect 9640 42508 9646 42560
rect 11256 42548 11284 42576
rect 12636 42548 12664 42576
rect 11256 42520 12664 42548
rect 13354 42508 13360 42560
rect 13412 42508 13418 42560
rect 13924 42557 13952 42588
rect 15654 42576 15660 42628
rect 15712 42576 15718 42628
rect 17497 42619 17555 42625
rect 16546 42588 17172 42616
rect 13909 42551 13967 42557
rect 13909 42517 13921 42551
rect 13955 42548 13967 42551
rect 14826 42548 14832 42560
rect 13955 42520 14832 42548
rect 13955 42517 13967 42520
rect 13909 42511 13967 42517
rect 14826 42508 14832 42520
rect 14884 42508 14890 42560
rect 15838 42508 15844 42560
rect 15896 42548 15902 42560
rect 16546 42548 16574 42588
rect 17144 42557 17172 42588
rect 17497 42585 17509 42619
rect 17543 42616 17555 42619
rect 18233 42619 18291 42625
rect 18233 42616 18245 42619
rect 17543 42588 18245 42616
rect 17543 42585 17555 42588
rect 17497 42579 17555 42585
rect 18233 42585 18245 42588
rect 18279 42616 18291 42619
rect 19794 42616 19800 42628
rect 18279 42588 19800 42616
rect 18279 42585 18291 42588
rect 18233 42579 18291 42585
rect 19794 42576 19800 42588
rect 19852 42616 19858 42628
rect 20530 42616 20536 42628
rect 19852 42588 20536 42616
rect 19852 42576 19858 42588
rect 20530 42576 20536 42588
rect 20588 42576 20594 42628
rect 20622 42576 20628 42628
rect 20680 42616 20686 42628
rect 23842 42616 23848 42628
rect 20680 42588 22968 42616
rect 23782 42588 23848 42616
rect 20680 42576 20686 42588
rect 15896 42520 16574 42548
rect 17129 42551 17187 42557
rect 15896 42508 15902 42520
rect 17129 42517 17141 42551
rect 17175 42517 17187 42551
rect 17129 42511 17187 42517
rect 19978 42508 19984 42560
rect 20036 42508 20042 42560
rect 20346 42508 20352 42560
rect 20404 42508 20410 42560
rect 21729 42551 21787 42557
rect 21729 42517 21741 42551
rect 21775 42548 21787 42551
rect 22186 42548 22192 42560
rect 21775 42520 22192 42548
rect 21775 42517 21787 42520
rect 21729 42511 21787 42517
rect 22186 42508 22192 42520
rect 22244 42508 22250 42560
rect 22940 42548 22968 42588
rect 23842 42576 23848 42588
rect 23900 42576 23906 42628
rect 23860 42548 23888 42576
rect 24044 42557 24072 42644
rect 22940 42520 23888 42548
rect 24029 42551 24087 42557
rect 24029 42517 24041 42551
rect 24075 42517 24087 42551
rect 24029 42511 24087 42517
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 4982 42304 4988 42356
rect 5040 42304 5046 42356
rect 9585 42347 9643 42353
rect 9585 42313 9597 42347
rect 9631 42344 9643 42347
rect 11330 42344 11336 42356
rect 9631 42316 11336 42344
rect 9631 42313 9643 42316
rect 9585 42307 9643 42313
rect 11330 42304 11336 42316
rect 11388 42304 11394 42356
rect 11698 42304 11704 42356
rect 11756 42304 11762 42356
rect 13354 42304 13360 42356
rect 13412 42304 13418 42356
rect 13722 42304 13728 42356
rect 13780 42304 13786 42356
rect 14366 42304 14372 42356
rect 14424 42344 14430 42356
rect 17129 42347 17187 42353
rect 17129 42344 17141 42347
rect 14424 42316 17141 42344
rect 14424 42304 14430 42316
rect 17129 42313 17141 42316
rect 17175 42313 17187 42347
rect 17129 42307 17187 42313
rect 17589 42347 17647 42353
rect 17589 42313 17601 42347
rect 17635 42344 17647 42347
rect 18417 42347 18475 42353
rect 18417 42344 18429 42347
rect 17635 42316 18429 42344
rect 17635 42313 17647 42316
rect 17589 42307 17647 42313
rect 18417 42313 18429 42316
rect 18463 42344 18475 42347
rect 18782 42344 18788 42356
rect 18463 42316 18788 42344
rect 18463 42313 18475 42316
rect 18417 42307 18475 42313
rect 18782 42304 18788 42316
rect 18840 42304 18846 42356
rect 19794 42344 19800 42356
rect 19352 42316 19800 42344
rect 3418 42236 3424 42288
rect 3476 42236 3482 42288
rect 3878 42236 3884 42288
rect 3936 42276 3942 42288
rect 4157 42279 4215 42285
rect 4157 42276 4169 42279
rect 3936 42248 4169 42276
rect 3936 42236 3942 42248
rect 4157 42245 4169 42248
rect 4203 42245 4215 42279
rect 8386 42276 8392 42288
rect 4157 42239 4215 42245
rect 7852 42248 8392 42276
rect 3605 42211 3663 42217
rect 3605 42177 3617 42211
rect 3651 42177 3663 42211
rect 3605 42171 3663 42177
rect 3145 42143 3203 42149
rect 3145 42109 3157 42143
rect 3191 42140 3203 42143
rect 3620 42140 3648 42171
rect 4338 42168 4344 42220
rect 4396 42168 4402 42220
rect 7852 42217 7880 42248
rect 8386 42236 8392 42248
rect 8444 42236 8450 42288
rect 14734 42276 14740 42288
rect 10060 42248 12296 42276
rect 5077 42211 5135 42217
rect 5077 42177 5089 42211
rect 5123 42208 5135 42211
rect 7837 42211 7895 42217
rect 5123 42180 5580 42208
rect 5123 42177 5135 42180
rect 5077 42171 5135 42177
rect 4890 42140 4896 42152
rect 3191 42112 4896 42140
rect 3191 42109 3203 42112
rect 3145 42103 3203 42109
rect 4890 42100 4896 42112
rect 4948 42100 4954 42152
rect 5552 42013 5580 42180
rect 7837 42177 7849 42211
rect 7883 42177 7895 42211
rect 7837 42171 7895 42177
rect 9214 42168 9220 42220
rect 9272 42168 9278 42220
rect 9490 42168 9496 42220
rect 9548 42208 9554 42220
rect 10060 42217 10088 42248
rect 10045 42211 10103 42217
rect 10045 42208 10057 42211
rect 9548 42180 10057 42208
rect 9548 42168 9554 42180
rect 10045 42177 10057 42180
rect 10091 42177 10103 42211
rect 10045 42171 10103 42177
rect 11790 42168 11796 42220
rect 11848 42208 11854 42220
rect 12069 42211 12127 42217
rect 12069 42208 12081 42211
rect 11848 42180 12081 42208
rect 11848 42168 11854 42180
rect 12069 42177 12081 42180
rect 12115 42177 12127 42211
rect 12069 42171 12127 42177
rect 7742 42100 7748 42152
rect 7800 42140 7806 42152
rect 12268 42149 12296 42248
rect 13188 42248 14740 42276
rect 13188 42149 13216 42248
rect 14734 42236 14740 42248
rect 14792 42236 14798 42288
rect 14918 42236 14924 42288
rect 14976 42276 14982 42288
rect 15105 42279 15163 42285
rect 15105 42276 15117 42279
rect 14976 42248 15117 42276
rect 14976 42236 14982 42248
rect 15105 42245 15117 42248
rect 15151 42245 15163 42279
rect 15105 42239 15163 42245
rect 16206 42236 16212 42288
rect 16264 42276 16270 42288
rect 19352 42276 19380 42316
rect 19794 42304 19800 42316
rect 19852 42344 19858 42356
rect 19852 42316 20852 42344
rect 19852 42304 19858 42316
rect 20622 42276 20628 42288
rect 16264 42248 16896 42276
rect 16264 42236 16270 42248
rect 13722 42168 13728 42220
rect 13780 42208 13786 42220
rect 14829 42211 14887 42217
rect 14829 42208 14841 42211
rect 13780 42180 14841 42208
rect 13780 42168 13786 42180
rect 14829 42177 14841 42180
rect 14875 42208 14887 42211
rect 15562 42208 15568 42220
rect 14875 42180 15568 42208
rect 14875 42177 14887 42180
rect 14829 42171 14887 42177
rect 15562 42168 15568 42180
rect 15620 42168 15626 42220
rect 16117 42211 16175 42217
rect 16117 42177 16129 42211
rect 16163 42208 16175 42211
rect 16574 42208 16580 42220
rect 16163 42180 16580 42208
rect 16163 42177 16175 42180
rect 16117 42171 16175 42177
rect 16574 42168 16580 42180
rect 16632 42168 16638 42220
rect 8113 42143 8171 42149
rect 8113 42140 8125 42143
rect 7800 42112 8125 42140
rect 7800 42100 7806 42112
rect 8113 42109 8125 42112
rect 8159 42109 8171 42143
rect 8113 42103 8171 42109
rect 12161 42143 12219 42149
rect 12161 42109 12173 42143
rect 12207 42109 12219 42143
rect 12161 42103 12219 42109
rect 12253 42143 12311 42149
rect 12253 42109 12265 42143
rect 12299 42109 12311 42143
rect 12253 42103 12311 42109
rect 13173 42143 13231 42149
rect 13173 42109 13185 42143
rect 13219 42109 13231 42143
rect 13173 42103 13231 42109
rect 13265 42143 13323 42149
rect 13265 42109 13277 42143
rect 13311 42140 13323 42143
rect 13354 42140 13360 42152
rect 13311 42112 13360 42140
rect 13311 42109 13323 42112
rect 13265 42103 13323 42109
rect 12176 42072 12204 42103
rect 13354 42100 13360 42112
rect 13412 42100 13418 42152
rect 16868 42149 16896 42248
rect 18708 42248 19380 42276
rect 20194 42248 20628 42276
rect 17497 42211 17555 42217
rect 17497 42177 17509 42211
rect 17543 42208 17555 42211
rect 18708 42208 18736 42248
rect 20622 42236 20628 42248
rect 20680 42236 20686 42288
rect 20824 42276 20852 42316
rect 21266 42304 21272 42356
rect 21324 42344 21330 42356
rect 22554 42344 22560 42356
rect 21324 42316 22560 42344
rect 21324 42304 21330 42316
rect 22554 42304 22560 42316
rect 22612 42304 22618 42356
rect 25133 42347 25191 42353
rect 25133 42344 25145 42347
rect 23124 42316 25145 42344
rect 23124 42276 23152 42316
rect 25133 42313 25145 42316
rect 25179 42313 25191 42347
rect 25133 42307 25191 42313
rect 20824 42248 23152 42276
rect 23842 42236 23848 42288
rect 23900 42236 23906 42288
rect 24394 42236 24400 42288
rect 24452 42236 24458 42288
rect 17543 42180 18736 42208
rect 20809 42211 20867 42217
rect 17543 42177 17555 42180
rect 17497 42171 17555 42177
rect 20809 42177 20821 42211
rect 20855 42208 20867 42211
rect 21453 42211 21511 42217
rect 21453 42208 21465 42211
rect 20855 42180 21465 42208
rect 20855 42177 20867 42180
rect 20809 42171 20867 42177
rect 21453 42177 21465 42180
rect 21499 42208 21511 42211
rect 21818 42208 21824 42220
rect 21499 42180 21824 42208
rect 21499 42177 21511 42180
rect 21453 42171 21511 42177
rect 21818 42168 21824 42180
rect 21876 42168 21882 42220
rect 22554 42168 22560 42220
rect 22612 42208 22618 42220
rect 25317 42211 25375 42217
rect 22612 42180 23152 42208
rect 22612 42168 22618 42180
rect 16853 42143 16911 42149
rect 16853 42109 16865 42143
rect 16899 42140 16911 42143
rect 17681 42143 17739 42149
rect 17681 42140 17693 42143
rect 16899 42112 17693 42140
rect 16899 42109 16911 42112
rect 16853 42103 16911 42109
rect 17681 42109 17693 42112
rect 17727 42109 17739 42143
rect 17681 42103 17739 42109
rect 18693 42143 18751 42149
rect 18693 42109 18705 42143
rect 18739 42109 18751 42143
rect 18693 42103 18751 42109
rect 18969 42143 19027 42149
rect 18969 42109 18981 42143
rect 19015 42140 19027 42143
rect 20990 42140 20996 42152
rect 19015 42112 20996 42140
rect 19015 42109 19027 42112
rect 18969 42103 19027 42109
rect 14734 42072 14740 42084
rect 12176 42044 14740 42072
rect 14734 42032 14740 42044
rect 14792 42032 14798 42084
rect 5537 42007 5595 42013
rect 5537 41973 5549 42007
rect 5583 42004 5595 42007
rect 6178 42004 6184 42016
rect 5583 41976 6184 42004
rect 5583 41973 5595 41976
rect 5537 41967 5595 41973
rect 6178 41964 6184 41976
rect 6236 41964 6242 42016
rect 10502 41964 10508 42016
rect 10560 42004 10566 42016
rect 10689 42007 10747 42013
rect 10689 42004 10701 42007
rect 10560 41976 10701 42004
rect 10560 41964 10566 41976
rect 10689 41973 10701 41976
rect 10735 41973 10747 42007
rect 10689 41967 10747 41973
rect 13906 41964 13912 42016
rect 13964 42004 13970 42016
rect 14185 42007 14243 42013
rect 14185 42004 14197 42007
rect 13964 41976 14197 42004
rect 13964 41964 13970 41976
rect 14185 41973 14197 41976
rect 14231 41973 14243 42007
rect 14185 41967 14243 41973
rect 15470 41964 15476 42016
rect 15528 41964 15534 42016
rect 15838 41964 15844 42016
rect 15896 42004 15902 42016
rect 18141 42007 18199 42013
rect 18141 42004 18153 42007
rect 15896 41976 18153 42004
rect 15896 41964 15902 41976
rect 18141 41973 18153 41976
rect 18187 41973 18199 42007
rect 18708 42004 18736 42103
rect 20990 42100 20996 42112
rect 21048 42100 21054 42152
rect 22189 42143 22247 42149
rect 22189 42109 22201 42143
rect 22235 42140 22247 42143
rect 22830 42140 22836 42152
rect 22235 42112 22836 42140
rect 22235 42109 22247 42112
rect 22189 42103 22247 42109
rect 22830 42100 22836 42112
rect 22888 42100 22894 42152
rect 23124 42140 23152 42180
rect 25317 42177 25329 42211
rect 25363 42208 25375 42211
rect 25363 42180 25452 42208
rect 25363 42177 25375 42180
rect 25317 42171 25375 42177
rect 24673 42143 24731 42149
rect 23124 42112 24624 42140
rect 20070 42032 20076 42084
rect 20128 42072 20134 42084
rect 21269 42075 21327 42081
rect 21269 42072 21281 42075
rect 20128 42044 21281 42072
rect 20128 42032 20134 42044
rect 21269 42041 21281 42044
rect 21315 42041 21327 42075
rect 24596 42072 24624 42112
rect 24673 42109 24685 42143
rect 24719 42140 24731 42143
rect 24719 42112 25360 42140
rect 24719 42109 24731 42112
rect 24673 42103 24731 42109
rect 25332 42084 25360 42112
rect 24854 42072 24860 42084
rect 24596 42044 24860 42072
rect 21269 42035 21327 42041
rect 24854 42032 24860 42044
rect 24912 42032 24918 42084
rect 25314 42032 25320 42084
rect 25372 42032 25378 42084
rect 25424 42016 25452 42180
rect 18966 42004 18972 42016
rect 18708 41976 18972 42004
rect 18141 41967 18199 41973
rect 18966 41964 18972 41976
rect 19024 42004 19030 42016
rect 19426 42004 19432 42016
rect 19024 41976 19432 42004
rect 19024 41964 19030 41976
rect 19426 41964 19432 41976
rect 19484 41964 19490 42016
rect 20162 41964 20168 42016
rect 20220 42004 20226 42016
rect 20441 42007 20499 42013
rect 20441 42004 20453 42007
rect 20220 41976 20453 42004
rect 20220 41964 20226 41976
rect 20441 41973 20453 41976
rect 20487 41973 20499 42007
rect 20441 41967 20499 41973
rect 20898 41964 20904 42016
rect 20956 41964 20962 42016
rect 22554 41964 22560 42016
rect 22612 42004 22618 42016
rect 22925 42007 22983 42013
rect 22925 42004 22937 42007
rect 22612 41976 22937 42004
rect 22612 41964 22618 41976
rect 22925 41973 22937 41976
rect 22971 41973 22983 42007
rect 22925 41967 22983 41973
rect 23198 41964 23204 42016
rect 23256 42004 23262 42016
rect 25406 42004 25412 42016
rect 23256 41976 25412 42004
rect 23256 41964 23262 41976
rect 25406 41964 25412 41976
rect 25464 41964 25470 42016
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 4065 41803 4123 41809
rect 4065 41769 4077 41803
rect 4111 41800 4123 41803
rect 4338 41800 4344 41812
rect 4111 41772 4344 41800
rect 4111 41769 4123 41772
rect 4065 41763 4123 41769
rect 4338 41760 4344 41772
rect 4396 41760 4402 41812
rect 8021 41803 8079 41809
rect 8021 41769 8033 41803
rect 8067 41800 8079 41803
rect 8570 41800 8576 41812
rect 8067 41772 8576 41800
rect 8067 41769 8079 41772
rect 8021 41763 8079 41769
rect 8570 41760 8576 41772
rect 8628 41760 8634 41812
rect 9401 41803 9459 41809
rect 9401 41769 9413 41803
rect 9447 41800 9459 41803
rect 9490 41800 9496 41812
rect 9447 41772 9496 41800
rect 9447 41769 9459 41772
rect 9401 41763 9459 41769
rect 9490 41760 9496 41772
rect 9548 41760 9554 41812
rect 11517 41803 11575 41809
rect 11517 41769 11529 41803
rect 11563 41800 11575 41803
rect 12618 41800 12624 41812
rect 11563 41772 12624 41800
rect 11563 41769 11575 41772
rect 11517 41763 11575 41769
rect 3694 41692 3700 41744
rect 3752 41732 3758 41744
rect 4525 41735 4583 41741
rect 4525 41732 4537 41735
rect 3752 41704 4537 41732
rect 3752 41692 3758 41704
rect 4525 41701 4537 41704
rect 4571 41701 4583 41735
rect 4525 41695 4583 41701
rect 8297 41735 8355 41741
rect 8297 41701 8309 41735
rect 8343 41732 8355 41735
rect 8343 41704 9260 41732
rect 8343 41701 8355 41704
rect 8297 41695 8355 41701
rect 6273 41667 6331 41673
rect 6273 41633 6285 41667
rect 6319 41664 6331 41667
rect 8386 41664 8392 41676
rect 6319 41636 8392 41664
rect 6319 41633 6331 41636
rect 6273 41627 6331 41633
rect 8386 41624 8392 41636
rect 8444 41624 8450 41676
rect 7558 41556 7564 41608
rect 7616 41596 7622 41608
rect 8496 41596 8524 41704
rect 9232 41676 9260 41704
rect 9214 41624 9220 41676
rect 9272 41664 9278 41676
rect 11532 41664 11560 41763
rect 12618 41760 12624 41772
rect 12676 41760 12682 41812
rect 14366 41760 14372 41812
rect 14424 41800 14430 41812
rect 16666 41800 16672 41812
rect 14424 41772 16672 41800
rect 14424 41760 14430 41772
rect 16666 41760 16672 41772
rect 16724 41760 16730 41812
rect 17586 41760 17592 41812
rect 17644 41800 17650 41812
rect 18693 41803 18751 41809
rect 18693 41800 18705 41803
rect 17644 41772 18705 41800
rect 17644 41760 17650 41772
rect 18693 41769 18705 41772
rect 18739 41800 18751 41803
rect 18739 41772 22094 41800
rect 18739 41769 18751 41772
rect 18693 41763 18751 41769
rect 16684 41732 16712 41760
rect 22066 41732 22094 41772
rect 22554 41760 22560 41812
rect 22612 41800 22618 41812
rect 25222 41800 25228 41812
rect 22612 41772 25228 41800
rect 22612 41760 22618 41772
rect 24029 41735 24087 41741
rect 16684 41704 17080 41732
rect 22066 41704 23520 41732
rect 9272 41636 11560 41664
rect 14553 41667 14611 41673
rect 9272 41624 9278 41636
rect 7616 41568 8524 41596
rect 9784 41582 9812 41636
rect 14553 41633 14565 41667
rect 14599 41664 14611 41667
rect 15194 41664 15200 41676
rect 14599 41636 15200 41664
rect 14599 41633 14611 41636
rect 14553 41627 14611 41633
rect 15194 41624 15200 41636
rect 15252 41624 15258 41676
rect 16025 41667 16083 41673
rect 16025 41633 16037 41667
rect 16071 41664 16083 41667
rect 16574 41664 16580 41676
rect 16071 41636 16580 41664
rect 16071 41633 16083 41636
rect 16025 41627 16083 41633
rect 16574 41624 16580 41636
rect 16632 41624 16638 41676
rect 16942 41624 16948 41676
rect 17000 41624 17006 41676
rect 17052 41673 17080 41704
rect 17037 41667 17095 41673
rect 17037 41633 17049 41667
rect 17083 41633 17095 41667
rect 17862 41664 17868 41676
rect 17037 41627 17095 41633
rect 17236 41636 17868 41664
rect 11149 41599 11207 41605
rect 7616 41556 7622 41568
rect 11149 41565 11161 41599
rect 11195 41596 11207 41599
rect 11698 41596 11704 41608
rect 11195 41568 11704 41596
rect 11195 41565 11207 41568
rect 11149 41559 11207 41565
rect 11698 41556 11704 41568
rect 11756 41596 11762 41608
rect 12710 41596 12716 41608
rect 11756 41568 12716 41596
rect 11756 41556 11762 41568
rect 12710 41556 12716 41568
rect 12768 41596 12774 41608
rect 12897 41599 12955 41605
rect 12897 41596 12909 41599
rect 12768 41568 12909 41596
rect 12768 41556 12774 41568
rect 12897 41565 12909 41568
rect 12943 41596 12955 41599
rect 14182 41596 14188 41608
rect 12943 41568 14188 41596
rect 12943 41565 12955 41568
rect 12897 41559 12955 41565
rect 14182 41556 14188 41568
rect 14240 41596 14246 41608
rect 14277 41599 14335 41605
rect 14277 41596 14289 41599
rect 14240 41568 14289 41596
rect 14240 41556 14246 41568
rect 14277 41565 14289 41568
rect 14323 41565 14335 41599
rect 14277 41559 14335 41565
rect 15654 41556 15660 41608
rect 15712 41596 15718 41608
rect 17236 41596 17264 41636
rect 17862 41624 17868 41636
rect 17920 41624 17926 41676
rect 19426 41624 19432 41676
rect 19484 41664 19490 41676
rect 19521 41667 19579 41673
rect 19521 41664 19533 41667
rect 19484 41636 19533 41664
rect 19484 41624 19490 41636
rect 19521 41633 19533 41636
rect 19567 41633 19579 41667
rect 19521 41627 19579 41633
rect 22002 41624 22008 41676
rect 22060 41664 22066 41676
rect 22189 41667 22247 41673
rect 22189 41664 22201 41667
rect 22060 41636 22201 41664
rect 22060 41624 22066 41636
rect 22189 41633 22201 41636
rect 22235 41633 22247 41667
rect 22189 41627 22247 41633
rect 22738 41624 22744 41676
rect 22796 41664 22802 41676
rect 23385 41667 23443 41673
rect 23385 41664 23397 41667
rect 22796 41636 23397 41664
rect 22796 41624 22802 41636
rect 23385 41633 23397 41636
rect 23431 41633 23443 41667
rect 23385 41627 23443 41633
rect 15712 41568 17264 41596
rect 15712 41556 15718 41568
rect 17310 41556 17316 41608
rect 17368 41596 17374 41608
rect 17681 41599 17739 41605
rect 17681 41596 17693 41599
rect 17368 41568 17693 41596
rect 17368 41556 17374 41568
rect 17681 41565 17693 41568
rect 17727 41596 17739 41599
rect 20714 41596 20720 41608
rect 17727 41568 20720 41596
rect 17727 41565 17739 41568
rect 17681 41559 17739 41565
rect 20714 41556 20720 41568
rect 20772 41556 20778 41608
rect 20806 41556 20812 41608
rect 20864 41556 20870 41608
rect 22830 41556 22836 41608
rect 22888 41596 22894 41608
rect 23201 41599 23259 41605
rect 23201 41596 23213 41599
rect 22888 41568 23213 41596
rect 22888 41556 22894 41568
rect 23201 41565 23213 41568
rect 23247 41565 23259 41599
rect 23492 41596 23520 41704
rect 24029 41701 24041 41735
rect 24075 41732 24087 41735
rect 24486 41732 24492 41744
rect 24075 41704 24492 41732
rect 24075 41701 24087 41704
rect 24029 41695 24087 41701
rect 24486 41692 24492 41704
rect 24544 41692 24550 41744
rect 25056 41732 25084 41772
rect 25222 41760 25228 41772
rect 25280 41760 25286 41812
rect 25056 41704 25176 41732
rect 23842 41624 23848 41676
rect 23900 41664 23906 41676
rect 24762 41664 24768 41676
rect 23900 41636 24768 41664
rect 23900 41624 23906 41636
rect 24762 41624 24768 41636
rect 24820 41624 24826 41676
rect 25038 41624 25044 41676
rect 25096 41624 25102 41676
rect 25148 41673 25176 41704
rect 25133 41667 25191 41673
rect 25133 41633 25145 41667
rect 25179 41633 25191 41667
rect 25133 41627 25191 41633
rect 23492 41568 25084 41596
rect 23201 41559 23259 41565
rect 25056 41540 25084 41568
rect 4709 41531 4767 41537
rect 4709 41497 4721 41531
rect 4755 41528 4767 41531
rect 5074 41528 5080 41540
rect 4755 41500 5080 41528
rect 4755 41497 4767 41500
rect 4709 41491 4767 41497
rect 5074 41488 5080 41500
rect 5132 41488 5138 41540
rect 6546 41488 6552 41540
rect 6604 41488 6610 41540
rect 10873 41531 10931 41537
rect 10873 41497 10885 41531
rect 10919 41528 10931 41531
rect 11238 41528 11244 41540
rect 10919 41500 11244 41528
rect 10919 41497 10931 41500
rect 10873 41491 10931 41497
rect 11238 41488 11244 41500
rect 11296 41488 11302 41540
rect 12066 41488 12072 41540
rect 12124 41528 12130 41540
rect 18969 41531 19027 41537
rect 18969 41528 18981 41531
rect 12124 41500 12434 41528
rect 12124 41488 12130 41500
rect 12406 41460 12434 41500
rect 16316 41500 18981 41528
rect 13357 41463 13415 41469
rect 13357 41460 13369 41463
rect 12406 41432 13369 41460
rect 13357 41429 13369 41432
rect 13403 41460 13415 41463
rect 16316 41460 16344 41500
rect 18969 41497 18981 41500
rect 19015 41528 19027 41531
rect 20349 41531 20407 41537
rect 20349 41528 20361 41531
rect 19015 41500 20361 41528
rect 19015 41497 19027 41500
rect 18969 41491 19027 41497
rect 20349 41497 20361 41500
rect 20395 41528 20407 41531
rect 20898 41528 20904 41540
rect 20395 41500 20904 41528
rect 20395 41497 20407 41500
rect 20349 41491 20407 41497
rect 20898 41488 20904 41500
rect 20956 41528 20962 41540
rect 21266 41528 21272 41540
rect 20956 41500 21272 41528
rect 20956 41488 20962 41500
rect 21266 41488 21272 41500
rect 21324 41528 21330 41540
rect 21453 41531 21511 41537
rect 21453 41528 21465 41531
rect 21324 41500 21465 41528
rect 21324 41488 21330 41500
rect 21453 41497 21465 41500
rect 21499 41497 21511 41531
rect 21453 41491 21511 41497
rect 21542 41488 21548 41540
rect 21600 41528 21606 41540
rect 23293 41531 23351 41537
rect 23293 41528 23305 41531
rect 21600 41500 23305 41528
rect 21600 41488 21606 41500
rect 23293 41497 23305 41500
rect 23339 41497 23351 41531
rect 23293 41491 23351 41497
rect 25038 41488 25044 41540
rect 25096 41528 25102 41540
rect 25590 41528 25596 41540
rect 25096 41500 25596 41528
rect 25096 41488 25102 41500
rect 25590 41488 25596 41500
rect 25648 41488 25654 41540
rect 13403 41432 16344 41460
rect 13403 41429 13415 41432
rect 13357 41423 13415 41429
rect 16390 41420 16396 41472
rect 16448 41460 16454 41472
rect 16485 41463 16543 41469
rect 16485 41460 16497 41463
rect 16448 41432 16497 41460
rect 16448 41420 16454 41432
rect 16485 41429 16497 41432
rect 16531 41429 16543 41463
rect 16485 41423 16543 41429
rect 16853 41463 16911 41469
rect 16853 41429 16865 41463
rect 16899 41460 16911 41463
rect 17586 41460 17592 41472
rect 16899 41432 17592 41460
rect 16899 41429 16911 41432
rect 16853 41423 16911 41429
rect 17586 41420 17592 41432
rect 17644 41420 17650 41472
rect 18325 41463 18383 41469
rect 18325 41429 18337 41463
rect 18371 41460 18383 41463
rect 18506 41460 18512 41472
rect 18371 41432 18512 41460
rect 18371 41429 18383 41432
rect 18325 41423 18383 41429
rect 18506 41420 18512 41432
rect 18564 41420 18570 41472
rect 20990 41420 20996 41472
rect 21048 41420 21054 41472
rect 22462 41420 22468 41472
rect 22520 41460 22526 41472
rect 22738 41460 22744 41472
rect 22520 41432 22744 41460
rect 22520 41420 22526 41432
rect 22738 41420 22744 41432
rect 22796 41420 22802 41472
rect 22830 41420 22836 41472
rect 22888 41420 22894 41472
rect 24210 41420 24216 41472
rect 24268 41420 24274 41472
rect 24578 41420 24584 41472
rect 24636 41420 24642 41472
rect 24946 41420 24952 41472
rect 25004 41420 25010 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 4062 41216 4068 41268
rect 4120 41256 4126 41268
rect 10873 41259 10931 41265
rect 10873 41256 10885 41259
rect 4120 41228 10885 41256
rect 4120 41216 4126 41228
rect 10873 41225 10885 41228
rect 10919 41256 10931 41259
rect 10962 41256 10968 41268
rect 10919 41228 10968 41256
rect 10919 41225 10931 41228
rect 10873 41219 10931 41225
rect 10962 41216 10968 41228
rect 11020 41216 11026 41268
rect 11333 41259 11391 41265
rect 11333 41225 11345 41259
rect 11379 41256 11391 41259
rect 12066 41256 12072 41268
rect 11379 41228 12072 41256
rect 11379 41225 11391 41228
rect 11333 41219 11391 41225
rect 7558 41148 7564 41200
rect 7616 41148 7622 41200
rect 10410 41188 10416 41200
rect 8496 41160 10416 41188
rect 1302 41080 1308 41132
rect 1360 41120 1366 41132
rect 1581 41123 1639 41129
rect 1581 41120 1593 41123
rect 1360 41092 1593 41120
rect 1360 41080 1366 41092
rect 1581 41089 1593 41092
rect 1627 41120 1639 41123
rect 2041 41123 2099 41129
rect 2041 41120 2053 41123
rect 1627 41092 2053 41120
rect 1627 41089 1639 41092
rect 1581 41083 1639 41089
rect 2041 41089 2053 41092
rect 2087 41089 2099 41123
rect 2041 41083 2099 41089
rect 8110 41012 8116 41064
rect 8168 41012 8174 41064
rect 8386 41012 8392 41064
rect 8444 41052 8450 41064
rect 8496 41052 8524 41160
rect 10410 41148 10416 41160
rect 10468 41148 10474 41200
rect 9677 41123 9735 41129
rect 9677 41089 9689 41123
rect 9723 41120 9735 41123
rect 10594 41120 10600 41132
rect 9723 41092 10600 41120
rect 9723 41089 9735 41092
rect 9677 41083 9735 41089
rect 10594 41080 10600 41092
rect 10652 41120 10658 41132
rect 11348 41120 11376 41219
rect 12066 41216 12072 41228
rect 12124 41216 12130 41268
rect 13265 41259 13323 41265
rect 13265 41225 13277 41259
rect 13311 41256 13323 41259
rect 13722 41256 13728 41268
rect 13311 41228 13728 41256
rect 13311 41225 13323 41228
rect 13265 41219 13323 41225
rect 13722 41216 13728 41228
rect 13780 41216 13786 41268
rect 13814 41216 13820 41268
rect 13872 41256 13878 41268
rect 14826 41256 14832 41268
rect 13872 41228 14832 41256
rect 13872 41216 13878 41228
rect 14826 41216 14832 41228
rect 14884 41216 14890 41268
rect 15749 41259 15807 41265
rect 15749 41225 15761 41259
rect 15795 41256 15807 41259
rect 15838 41256 15844 41268
rect 15795 41228 15844 41256
rect 15795 41225 15807 41228
rect 15749 41219 15807 41225
rect 15838 41216 15844 41228
rect 15896 41216 15902 41268
rect 17129 41259 17187 41265
rect 17129 41225 17141 41259
rect 17175 41256 17187 41259
rect 17218 41256 17224 41268
rect 17175 41228 17224 41256
rect 17175 41225 17187 41228
rect 17129 41219 17187 41225
rect 17218 41216 17224 41228
rect 17276 41216 17282 41268
rect 18414 41216 18420 41268
rect 18472 41256 18478 41268
rect 18509 41259 18567 41265
rect 18509 41256 18521 41259
rect 18472 41228 18521 41256
rect 18472 41216 18478 41228
rect 18509 41225 18521 41228
rect 18555 41225 18567 41259
rect 18509 41219 18567 41225
rect 18690 41216 18696 41268
rect 18748 41256 18754 41268
rect 19058 41256 19064 41268
rect 18748 41228 19064 41256
rect 18748 41216 18754 41228
rect 19058 41216 19064 41228
rect 19116 41216 19122 41268
rect 19886 41216 19892 41268
rect 19944 41216 19950 41268
rect 19978 41216 19984 41268
rect 20036 41256 20042 41268
rect 20625 41259 20683 41265
rect 20625 41256 20637 41259
rect 20036 41228 20637 41256
rect 20036 41216 20042 41228
rect 20625 41225 20637 41228
rect 20671 41225 20683 41259
rect 20625 41219 20683 41225
rect 20806 41216 20812 41268
rect 20864 41256 20870 41268
rect 22002 41256 22008 41268
rect 20864 41228 22008 41256
rect 20864 41216 20870 41228
rect 22002 41216 22008 41228
rect 22060 41216 22066 41268
rect 22646 41216 22652 41268
rect 22704 41216 22710 41268
rect 22741 41259 22799 41265
rect 22741 41225 22753 41259
rect 22787 41256 22799 41259
rect 22830 41256 22836 41268
rect 22787 41228 22836 41256
rect 22787 41225 22799 41228
rect 22741 41219 22799 41225
rect 22830 41216 22836 41228
rect 22888 41216 22894 41268
rect 23109 41259 23167 41265
rect 23109 41225 23121 41259
rect 23155 41256 23167 41259
rect 23934 41256 23940 41268
rect 23155 41228 23940 41256
rect 23155 41225 23167 41228
rect 23109 41219 23167 41225
rect 23934 41216 23940 41228
rect 23992 41216 23998 41268
rect 11422 41148 11428 41200
rect 11480 41188 11486 41200
rect 16482 41188 16488 41200
rect 11480 41160 12434 41188
rect 11480 41148 11486 41160
rect 10652 41092 11376 41120
rect 12069 41123 12127 41129
rect 10652 41080 10658 41092
rect 12069 41089 12081 41123
rect 12115 41089 12127 41123
rect 12069 41083 12127 41089
rect 8444 41024 8524 41052
rect 8757 41055 8815 41061
rect 8444 41012 8450 41024
rect 8757 41021 8769 41055
rect 8803 41052 8815 41055
rect 9306 41052 9312 41064
rect 8803 41024 9312 41052
rect 8803 41021 8815 41024
rect 8757 41015 8815 41021
rect 9306 41012 9312 41024
rect 9364 41012 9370 41064
rect 10686 41012 10692 41064
rect 10744 41052 10750 41064
rect 12084 41052 12112 41083
rect 10744 41024 12112 41052
rect 12161 41055 12219 41061
rect 10744 41012 10750 41024
rect 12161 41021 12173 41055
rect 12207 41021 12219 41055
rect 12161 41015 12219 41021
rect 3418 40944 3424 40996
rect 3476 40984 3482 40996
rect 8846 40984 8852 40996
rect 3476 40956 7144 40984
rect 3476 40944 3482 40956
rect 1765 40919 1823 40925
rect 1765 40885 1777 40919
rect 1811 40916 1823 40919
rect 3694 40916 3700 40928
rect 1811 40888 3700 40916
rect 1811 40885 1823 40888
rect 1765 40879 1823 40885
rect 3694 40876 3700 40888
rect 3752 40876 3758 40928
rect 6638 40876 6644 40928
rect 6696 40876 6702 40928
rect 7116 40916 7144 40956
rect 8588 40956 8852 40984
rect 8588 40916 8616 40956
rect 8846 40944 8852 40956
rect 8904 40984 8910 40996
rect 10134 40984 10140 40996
rect 8904 40956 10140 40984
rect 8904 40944 8910 40956
rect 10134 40944 10140 40956
rect 10192 40944 10198 40996
rect 11606 40944 11612 40996
rect 11664 40984 11670 40996
rect 11701 40987 11759 40993
rect 11701 40984 11713 40987
rect 11664 40956 11713 40984
rect 11664 40944 11670 40956
rect 11701 40953 11713 40956
rect 11747 40953 11759 40987
rect 12176 40984 12204 41015
rect 12250 41012 12256 41064
rect 12308 41012 12314 41064
rect 12406 41052 12434 41160
rect 15028 41160 16488 41188
rect 12805 41123 12863 41129
rect 12805 41089 12817 41123
rect 12851 41120 12863 41123
rect 13446 41120 13452 41132
rect 12851 41092 13452 41120
rect 12851 41089 12863 41092
rect 12805 41083 12863 41089
rect 13446 41080 13452 41092
rect 13504 41080 13510 41132
rect 13630 41080 13636 41132
rect 13688 41080 13694 41132
rect 15028 41129 15056 41160
rect 16482 41148 16488 41160
rect 16540 41188 16546 41200
rect 18966 41188 18972 41200
rect 16540 41160 18972 41188
rect 16540 41148 16546 41160
rect 18966 41148 18972 41160
rect 19024 41148 19030 41200
rect 19076 41160 21128 41188
rect 15013 41123 15071 41129
rect 15013 41089 15025 41123
rect 15059 41089 15071 41123
rect 15013 41083 15071 41089
rect 15286 41080 15292 41132
rect 15344 41120 15350 41132
rect 15841 41123 15899 41129
rect 15344 41092 15608 41120
rect 15344 41080 15350 41092
rect 15580 41064 15608 41092
rect 15841 41089 15853 41123
rect 15887 41089 15899 41123
rect 15841 41083 15899 41089
rect 14737 41055 14795 41061
rect 12406 41024 13768 41052
rect 13538 40984 13544 40996
rect 12176 40956 13544 40984
rect 11701 40947 11759 40953
rect 13538 40944 13544 40956
rect 13596 40944 13602 40996
rect 7116 40888 8616 40916
rect 9125 40919 9183 40925
rect 9125 40885 9137 40919
rect 9171 40916 9183 40919
rect 9214 40916 9220 40928
rect 9171 40888 9220 40916
rect 9171 40885 9183 40888
rect 9125 40879 9183 40885
rect 9214 40876 9220 40888
rect 9272 40876 9278 40928
rect 10410 40876 10416 40928
rect 10468 40916 10474 40928
rect 11057 40919 11115 40925
rect 11057 40916 11069 40919
rect 10468 40888 11069 40916
rect 10468 40876 10474 40888
rect 11057 40885 11069 40888
rect 11103 40916 11115 40919
rect 11422 40916 11428 40928
rect 11103 40888 11428 40916
rect 11103 40885 11115 40888
rect 11057 40879 11115 40885
rect 11422 40876 11428 40888
rect 11480 40876 11486 40928
rect 11974 40876 11980 40928
rect 12032 40916 12038 40928
rect 13446 40916 13452 40928
rect 12032 40888 13452 40916
rect 12032 40876 12038 40888
rect 13446 40876 13452 40888
rect 13504 40876 13510 40928
rect 13740 40916 13768 41024
rect 14737 41021 14749 41055
rect 14783 41052 14795 41055
rect 15470 41052 15476 41064
rect 14783 41024 15476 41052
rect 14783 41021 14795 41024
rect 14737 41015 14795 41021
rect 15470 41012 15476 41024
rect 15528 41012 15534 41064
rect 15562 41012 15568 41064
rect 15620 41012 15626 41064
rect 15856 41052 15884 41083
rect 15930 41080 15936 41132
rect 15988 41120 15994 41132
rect 17221 41123 17279 41129
rect 17221 41120 17233 41123
rect 15988 41092 17233 41120
rect 15988 41080 15994 41092
rect 17221 41089 17233 41092
rect 17267 41089 17279 41123
rect 17221 41083 17279 41089
rect 18598 41080 18604 41132
rect 18656 41080 18662 41132
rect 15856 41024 15976 41052
rect 15948 40984 15976 41024
rect 17034 41012 17040 41064
rect 17092 41012 17098 41064
rect 18322 41012 18328 41064
rect 18380 41012 18386 41064
rect 17957 40987 18015 40993
rect 17957 40984 17969 40987
rect 15948 40956 17969 40984
rect 17957 40953 17969 40956
rect 18003 40984 18015 40987
rect 19076 40984 19104 41160
rect 19797 41123 19855 41129
rect 19797 41089 19809 41123
rect 19843 41120 19855 41123
rect 19886 41120 19892 41132
rect 19843 41092 19892 41120
rect 19843 41089 19855 41092
rect 19797 41083 19855 41089
rect 19886 41080 19892 41092
rect 19944 41080 19950 41132
rect 20993 41123 21051 41129
rect 20993 41089 21005 41123
rect 21039 41089 21051 41123
rect 21100 41120 21128 41160
rect 21174 41148 21180 41200
rect 21232 41188 21238 41200
rect 21232 41160 24808 41188
rect 21232 41148 21238 41160
rect 22462 41120 22468 41132
rect 21100 41092 22468 41120
rect 20993 41083 21051 41089
rect 19150 41012 19156 41064
rect 19208 41052 19214 41064
rect 19981 41055 20039 41061
rect 19981 41052 19993 41055
rect 19208 41024 19993 41052
rect 19208 41012 19214 41024
rect 19981 41021 19993 41024
rect 20027 41021 20039 41055
rect 19981 41015 20039 41021
rect 18003 40956 19104 40984
rect 21008 40984 21036 41083
rect 22462 41080 22468 41092
rect 22520 41080 22526 41132
rect 24486 41080 24492 41132
rect 24544 41080 24550 41132
rect 24780 41129 24808 41160
rect 24765 41123 24823 41129
rect 24765 41089 24777 41123
rect 24811 41089 24823 41123
rect 24765 41083 24823 41089
rect 21082 41012 21088 41064
rect 21140 41012 21146 41064
rect 21269 41055 21327 41061
rect 21269 41021 21281 41055
rect 21315 41052 21327 41055
rect 21910 41052 21916 41064
rect 21315 41024 21916 41052
rect 21315 41021 21327 41024
rect 21269 41015 21327 41021
rect 21910 41012 21916 41024
rect 21968 41012 21974 41064
rect 22557 41055 22615 41061
rect 22557 41021 22569 41055
rect 22603 41052 22615 41055
rect 22738 41052 22744 41064
rect 22603 41024 22744 41052
rect 22603 41021 22615 41024
rect 22557 41015 22615 41021
rect 22738 41012 22744 41024
rect 22796 41012 22802 41064
rect 23750 41012 23756 41064
rect 23808 41012 23814 41064
rect 21008 40956 21956 40984
rect 18003 40953 18015 40956
rect 17957 40947 18015 40953
rect 15286 40916 15292 40928
rect 13740 40888 15292 40916
rect 15286 40876 15292 40888
rect 15344 40876 15350 40928
rect 16209 40919 16267 40925
rect 16209 40885 16221 40919
rect 16255 40916 16267 40919
rect 16298 40916 16304 40928
rect 16255 40888 16304 40916
rect 16255 40885 16267 40888
rect 16209 40879 16267 40885
rect 16298 40876 16304 40888
rect 16356 40876 16362 40928
rect 17586 40876 17592 40928
rect 17644 40876 17650 40928
rect 18690 40876 18696 40928
rect 18748 40916 18754 40928
rect 18969 40919 19027 40925
rect 18969 40916 18981 40919
rect 18748 40888 18981 40916
rect 18748 40876 18754 40888
rect 18969 40885 18981 40888
rect 19015 40885 19027 40919
rect 18969 40879 19027 40885
rect 19426 40876 19432 40928
rect 19484 40876 19490 40928
rect 21082 40876 21088 40928
rect 21140 40916 21146 40928
rect 21450 40916 21456 40928
rect 21140 40888 21456 40916
rect 21140 40876 21146 40888
rect 21450 40876 21456 40888
rect 21508 40916 21514 40928
rect 21821 40919 21879 40925
rect 21821 40916 21833 40919
rect 21508 40888 21833 40916
rect 21508 40876 21514 40888
rect 21821 40885 21833 40888
rect 21867 40885 21879 40919
rect 21928 40916 21956 40956
rect 22002 40944 22008 40996
rect 22060 40984 22066 40996
rect 22060 40956 23520 40984
rect 22060 40944 22066 40956
rect 22097 40919 22155 40925
rect 22097 40916 22109 40919
rect 21928 40888 22109 40916
rect 21821 40879 21879 40885
rect 22097 40885 22109 40888
rect 22143 40916 22155 40919
rect 22462 40916 22468 40928
rect 22143 40888 22468 40916
rect 22143 40885 22155 40888
rect 22097 40879 22155 40885
rect 22462 40876 22468 40888
rect 22520 40876 22526 40928
rect 23492 40925 23520 40956
rect 23477 40919 23535 40925
rect 23477 40885 23489 40919
rect 23523 40916 23535 40919
rect 24854 40916 24860 40928
rect 23523 40888 24860 40916
rect 23523 40885 23535 40888
rect 23477 40879 23535 40885
rect 24854 40876 24860 40888
rect 24912 40876 24918 40928
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 8110 40672 8116 40724
rect 8168 40712 8174 40724
rect 8389 40715 8447 40721
rect 8389 40712 8401 40715
rect 8168 40684 8401 40712
rect 8168 40672 8174 40684
rect 8389 40681 8401 40684
rect 8435 40681 8447 40715
rect 8389 40675 8447 40681
rect 10962 40672 10968 40724
rect 11020 40712 11026 40724
rect 11020 40684 12434 40712
rect 11020 40672 11026 40684
rect 7098 40604 7104 40656
rect 7156 40644 7162 40656
rect 10410 40644 10416 40656
rect 7156 40616 10416 40644
rect 7156 40604 7162 40616
rect 10410 40604 10416 40616
rect 10468 40644 10474 40656
rect 12406 40644 12434 40684
rect 13538 40672 13544 40724
rect 13596 40712 13602 40724
rect 13722 40712 13728 40724
rect 13596 40684 13728 40712
rect 13596 40672 13602 40684
rect 13722 40672 13728 40684
rect 13780 40672 13786 40724
rect 13909 40715 13967 40721
rect 13909 40681 13921 40715
rect 13955 40712 13967 40715
rect 13998 40712 14004 40724
rect 13955 40684 14004 40712
rect 13955 40681 13967 40684
rect 13909 40675 13967 40681
rect 13998 40672 14004 40684
rect 14056 40672 14062 40724
rect 14734 40672 14740 40724
rect 14792 40712 14798 40724
rect 15841 40715 15899 40721
rect 15841 40712 15853 40715
rect 14792 40684 15853 40712
rect 14792 40672 14798 40684
rect 15841 40681 15853 40684
rect 15887 40681 15899 40715
rect 15841 40675 15899 40681
rect 17310 40672 17316 40724
rect 17368 40712 17374 40724
rect 21913 40715 21971 40721
rect 21913 40712 21925 40715
rect 17368 40684 21925 40712
rect 17368 40672 17374 40684
rect 21913 40681 21925 40684
rect 21959 40681 21971 40715
rect 21913 40675 21971 40681
rect 22462 40672 22468 40724
rect 22520 40712 22526 40724
rect 25130 40712 25136 40724
rect 22520 40684 25136 40712
rect 22520 40672 22526 40684
rect 25130 40672 25136 40684
rect 25188 40672 25194 40724
rect 14458 40644 14464 40656
rect 10468 40616 10824 40644
rect 12406 40616 14464 40644
rect 10468 40604 10474 40616
rect 9030 40536 9036 40588
rect 9088 40576 9094 40588
rect 9309 40579 9367 40585
rect 9309 40576 9321 40579
rect 9088 40548 9321 40576
rect 9088 40536 9094 40548
rect 9309 40545 9321 40548
rect 9355 40545 9367 40579
rect 10796 40576 10824 40616
rect 14458 40604 14464 40616
rect 14516 40644 14522 40656
rect 16758 40644 16764 40656
rect 14516 40616 16764 40644
rect 14516 40604 14522 40616
rect 16758 40604 16764 40616
rect 16816 40604 16822 40656
rect 21726 40604 21732 40656
rect 21784 40604 21790 40656
rect 22002 40604 22008 40656
rect 22060 40644 22066 40656
rect 23845 40647 23903 40653
rect 23845 40644 23857 40647
rect 22060 40616 23857 40644
rect 22060 40604 22066 40616
rect 23845 40613 23857 40616
rect 23891 40613 23903 40647
rect 23845 40607 23903 40613
rect 10965 40579 11023 40585
rect 10965 40576 10977 40579
rect 10796 40548 10977 40576
rect 9309 40539 9367 40545
rect 10965 40545 10977 40548
rect 11011 40545 11023 40579
rect 10965 40539 11023 40545
rect 11701 40579 11759 40585
rect 11701 40545 11713 40579
rect 11747 40545 11759 40579
rect 11701 40539 11759 40545
rect 7190 40468 7196 40520
rect 7248 40508 7254 40520
rect 7745 40511 7803 40517
rect 7745 40508 7757 40511
rect 7248 40480 7757 40508
rect 7248 40468 7254 40480
rect 7745 40477 7757 40480
rect 7791 40508 7803 40511
rect 11716 40508 11744 40539
rect 12066 40536 12072 40588
rect 12124 40576 12130 40588
rect 12897 40579 12955 40585
rect 12897 40576 12909 40579
rect 12124 40548 12909 40576
rect 12124 40536 12130 40548
rect 12897 40545 12909 40548
rect 12943 40545 12955 40579
rect 12897 40539 12955 40545
rect 13081 40579 13139 40585
rect 13081 40545 13093 40579
rect 13127 40576 13139 40579
rect 13998 40576 14004 40588
rect 13127 40548 14004 40576
rect 13127 40545 13139 40548
rect 13081 40539 13139 40545
rect 13998 40536 14004 40548
rect 14056 40536 14062 40588
rect 14826 40536 14832 40588
rect 14884 40576 14890 40588
rect 15197 40579 15255 40585
rect 15197 40576 15209 40579
rect 14884 40548 15209 40576
rect 14884 40536 14890 40548
rect 15197 40545 15209 40548
rect 15243 40545 15255 40579
rect 15197 40539 15255 40545
rect 16298 40536 16304 40588
rect 16356 40536 16362 40588
rect 16393 40579 16451 40585
rect 16393 40545 16405 40579
rect 16439 40545 16451 40579
rect 16393 40539 16451 40545
rect 17129 40579 17187 40585
rect 17129 40545 17141 40579
rect 17175 40576 17187 40579
rect 17402 40576 17408 40588
rect 17175 40548 17408 40576
rect 17175 40545 17187 40548
rect 17129 40539 17187 40545
rect 7791 40480 11744 40508
rect 7791 40477 7803 40480
rect 7745 40471 7803 40477
rect 11974 40468 11980 40520
rect 12032 40468 12038 40520
rect 12526 40468 12532 40520
rect 12584 40508 12590 40520
rect 13173 40511 13231 40517
rect 13173 40508 13185 40511
rect 12584 40480 13185 40508
rect 12584 40468 12590 40480
rect 13173 40477 13185 40480
rect 13219 40477 13231 40511
rect 13173 40471 13231 40477
rect 13446 40468 13452 40520
rect 13504 40508 13510 40520
rect 16408 40508 16436 40539
rect 17402 40536 17408 40548
rect 17460 40536 17466 40588
rect 18506 40536 18512 40588
rect 18564 40576 18570 40588
rect 18601 40579 18659 40585
rect 18601 40576 18613 40579
rect 18564 40548 18613 40576
rect 18564 40536 18570 40548
rect 18601 40545 18613 40548
rect 18647 40545 18659 40579
rect 18601 40539 18659 40545
rect 18877 40579 18935 40585
rect 18877 40545 18889 40579
rect 18923 40576 18935 40579
rect 18966 40576 18972 40588
rect 18923 40548 18972 40576
rect 18923 40545 18935 40548
rect 18877 40539 18935 40545
rect 18966 40536 18972 40548
rect 19024 40536 19030 40588
rect 20714 40536 20720 40588
rect 20772 40576 20778 40588
rect 21269 40579 21327 40585
rect 21269 40576 21281 40579
rect 20772 40548 21281 40576
rect 20772 40536 20778 40548
rect 21269 40545 21281 40548
rect 21315 40545 21327 40579
rect 21744 40576 21772 40604
rect 21910 40576 21916 40588
rect 21744 40548 21916 40576
rect 21269 40539 21327 40545
rect 21910 40536 21916 40548
rect 21968 40536 21974 40588
rect 22554 40536 22560 40588
rect 22612 40576 22618 40588
rect 22649 40579 22707 40585
rect 22649 40576 22661 40579
rect 22612 40548 22661 40576
rect 22612 40536 22618 40548
rect 22649 40545 22661 40548
rect 22695 40545 22707 40579
rect 25498 40576 25504 40588
rect 22649 40539 22707 40545
rect 23860 40548 25504 40576
rect 20438 40508 20444 40520
rect 13504 40480 16436 40508
rect 18892 40480 20444 40508
rect 13504 40468 13510 40480
rect 8846 40400 8852 40452
rect 8904 40440 8910 40452
rect 9585 40443 9643 40449
rect 9585 40440 9597 40443
rect 8904 40412 9597 40440
rect 8904 40400 8910 40412
rect 9585 40409 9597 40412
rect 9631 40409 9643 40443
rect 9585 40403 9643 40409
rect 10778 40400 10784 40452
rect 10836 40440 10842 40452
rect 11238 40440 11244 40452
rect 10836 40412 11244 40440
rect 10836 40400 10842 40412
rect 11238 40400 11244 40412
rect 11296 40440 11302 40452
rect 11885 40443 11943 40449
rect 11885 40440 11897 40443
rect 11296 40412 11897 40440
rect 11296 40400 11302 40412
rect 11885 40409 11897 40412
rect 11931 40409 11943 40443
rect 11885 40403 11943 40409
rect 14461 40443 14519 40449
rect 14461 40409 14473 40443
rect 14507 40440 14519 40443
rect 14550 40440 14556 40452
rect 14507 40412 14556 40440
rect 14507 40409 14519 40412
rect 14461 40403 14519 40409
rect 14550 40400 14556 40412
rect 14608 40440 14614 40452
rect 14918 40440 14924 40452
rect 14608 40412 14924 40440
rect 14608 40400 14614 40412
rect 14918 40400 14924 40412
rect 14976 40400 14982 40452
rect 16209 40443 16267 40449
rect 16209 40409 16221 40443
rect 16255 40440 16267 40443
rect 16255 40412 17356 40440
rect 16255 40409 16267 40412
rect 16209 40403 16267 40409
rect 8757 40375 8815 40381
rect 8757 40341 8769 40375
rect 8803 40372 8815 40375
rect 9030 40372 9036 40384
rect 8803 40344 9036 40372
rect 8803 40341 8815 40344
rect 8757 40335 8815 40341
rect 9030 40332 9036 40344
rect 9088 40332 9094 40384
rect 9306 40332 9312 40384
rect 9364 40372 9370 40384
rect 9493 40375 9551 40381
rect 9493 40372 9505 40375
rect 9364 40344 9505 40372
rect 9364 40332 9370 40344
rect 9493 40341 9505 40344
rect 9539 40341 9551 40375
rect 9493 40335 9551 40341
rect 9953 40375 10011 40381
rect 9953 40341 9965 40375
rect 9999 40372 10011 40375
rect 10318 40372 10324 40384
rect 9999 40344 10324 40372
rect 9999 40341 10011 40344
rect 9953 40335 10011 40341
rect 10318 40332 10324 40344
rect 10376 40332 10382 40384
rect 10410 40332 10416 40384
rect 10468 40332 10474 40384
rect 10873 40375 10931 40381
rect 10873 40341 10885 40375
rect 10919 40372 10931 40375
rect 10962 40372 10968 40384
rect 10919 40344 10968 40372
rect 10919 40341 10931 40344
rect 10873 40335 10931 40341
rect 10962 40332 10968 40344
rect 11020 40332 11026 40384
rect 11054 40332 11060 40384
rect 11112 40372 11118 40384
rect 11422 40372 11428 40384
rect 11112 40344 11428 40372
rect 11112 40332 11118 40344
rect 11422 40332 11428 40344
rect 11480 40332 11486 40384
rect 12345 40375 12403 40381
rect 12345 40341 12357 40375
rect 12391 40372 12403 40375
rect 12710 40372 12716 40384
rect 12391 40344 12716 40372
rect 12391 40341 12403 40344
rect 12345 40335 12403 40341
rect 12710 40332 12716 40344
rect 12768 40332 12774 40384
rect 13538 40332 13544 40384
rect 13596 40332 13602 40384
rect 17328 40372 17356 40412
rect 17862 40400 17868 40452
rect 17920 40400 17926 40452
rect 18506 40400 18512 40452
rect 18564 40440 18570 40452
rect 18892 40440 18920 40480
rect 20438 40468 20444 40480
rect 20496 40468 20502 40520
rect 21174 40468 21180 40520
rect 21232 40508 21238 40520
rect 21634 40508 21640 40520
rect 21232 40480 21640 40508
rect 21232 40468 21238 40480
rect 21634 40468 21640 40480
rect 21692 40468 21698 40520
rect 22097 40511 22155 40517
rect 22097 40477 22109 40511
rect 22143 40508 22155 40511
rect 22186 40508 22192 40520
rect 22143 40480 22192 40508
rect 22143 40477 22155 40480
rect 22097 40471 22155 40477
rect 22186 40468 22192 40480
rect 22244 40468 22250 40520
rect 22925 40511 22983 40517
rect 22925 40477 22937 40511
rect 22971 40508 22983 40511
rect 23750 40508 23756 40520
rect 22971 40480 23756 40508
rect 22971 40477 22983 40480
rect 22925 40471 22983 40477
rect 23750 40468 23756 40480
rect 23808 40468 23814 40520
rect 18564 40412 18920 40440
rect 18564 40400 18570 40412
rect 19886 40400 19892 40452
rect 19944 40440 19950 40452
rect 20349 40443 20407 40449
rect 20349 40440 20361 40443
rect 19944 40412 20361 40440
rect 19944 40400 19950 40412
rect 20349 40409 20361 40412
rect 20395 40440 20407 40443
rect 20395 40412 21220 40440
rect 20395 40409 20407 40412
rect 20349 40403 20407 40409
rect 18966 40372 18972 40384
rect 17328 40344 18972 40372
rect 18966 40332 18972 40344
rect 19024 40332 19030 40384
rect 19518 40332 19524 40384
rect 19576 40372 19582 40384
rect 20717 40375 20775 40381
rect 20717 40372 20729 40375
rect 19576 40344 20729 40372
rect 19576 40332 19582 40344
rect 20717 40341 20729 40344
rect 20763 40341 20775 40375
rect 20717 40335 20775 40341
rect 21082 40332 21088 40384
rect 21140 40332 21146 40384
rect 21192 40372 21220 40412
rect 21726 40400 21732 40452
rect 21784 40440 21790 40452
rect 22833 40443 22891 40449
rect 22833 40440 22845 40443
rect 21784 40412 22845 40440
rect 21784 40400 21790 40412
rect 22833 40409 22845 40412
rect 22879 40409 22891 40443
rect 23860 40440 23888 40548
rect 25498 40536 25504 40548
rect 25556 40536 25562 40588
rect 24029 40511 24087 40517
rect 24029 40477 24041 40511
rect 24075 40508 24087 40511
rect 24210 40508 24216 40520
rect 24075 40480 24216 40508
rect 24075 40477 24087 40480
rect 24029 40471 24087 40477
rect 24210 40468 24216 40480
rect 24268 40508 24274 40520
rect 24486 40508 24492 40520
rect 24268 40480 24492 40508
rect 24268 40468 24274 40480
rect 24486 40468 24492 40480
rect 24544 40468 24550 40520
rect 24581 40511 24639 40517
rect 24581 40477 24593 40511
rect 24627 40477 24639 40511
rect 24581 40471 24639 40477
rect 22833 40403 22891 40409
rect 22940 40412 23888 40440
rect 22462 40372 22468 40384
rect 21192 40344 22468 40372
rect 22462 40332 22468 40344
rect 22520 40372 22526 40384
rect 22940 40372 22968 40412
rect 24302 40400 24308 40452
rect 24360 40440 24366 40452
rect 24596 40440 24624 40471
rect 24360 40412 24624 40440
rect 24360 40400 24366 40412
rect 22520 40344 22968 40372
rect 22520 40332 22526 40344
rect 23290 40332 23296 40384
rect 23348 40332 23354 40384
rect 25222 40332 25228 40384
rect 25280 40332 25286 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 11054 40128 11060 40180
rect 11112 40168 11118 40180
rect 11330 40168 11336 40180
rect 11112 40140 11336 40168
rect 11112 40128 11118 40140
rect 11330 40128 11336 40140
rect 11388 40168 11394 40180
rect 13446 40168 13452 40180
rect 11388 40140 13452 40168
rect 11388 40128 11394 40140
rect 13446 40128 13452 40140
rect 13504 40128 13510 40180
rect 15289 40171 15347 40177
rect 15289 40137 15301 40171
rect 15335 40168 15347 40171
rect 15930 40168 15936 40180
rect 15335 40140 15936 40168
rect 15335 40137 15347 40140
rect 15289 40131 15347 40137
rect 15930 40128 15936 40140
rect 15988 40128 15994 40180
rect 16850 40128 16856 40180
rect 16908 40128 16914 40180
rect 19426 40128 19432 40180
rect 19484 40168 19490 40180
rect 19521 40171 19579 40177
rect 19521 40168 19533 40171
rect 19484 40140 19533 40168
rect 19484 40128 19490 40140
rect 19521 40137 19533 40140
rect 19567 40137 19579 40171
rect 19521 40131 19579 40137
rect 19978 40128 19984 40180
rect 20036 40128 20042 40180
rect 21358 40168 21364 40180
rect 20916 40140 21364 40168
rect 8849 40103 8907 40109
rect 8849 40069 8861 40103
rect 8895 40100 8907 40103
rect 9030 40100 9036 40112
rect 8895 40072 9036 40100
rect 8895 40069 8907 40072
rect 8849 40063 8907 40069
rect 9030 40060 9036 40072
rect 9088 40060 9094 40112
rect 9214 40060 9220 40112
rect 9272 40100 9278 40112
rect 9272 40072 9430 40100
rect 9272 40060 9278 40072
rect 11974 40060 11980 40112
rect 12032 40060 12038 40112
rect 13630 40100 13636 40112
rect 13202 40072 13636 40100
rect 13630 40060 13636 40072
rect 13688 40100 13694 40112
rect 13817 40103 13875 40109
rect 13817 40100 13829 40103
rect 13688 40072 13829 40100
rect 13688 40060 13694 40072
rect 13817 40069 13829 40072
rect 13863 40069 13875 40103
rect 13817 40063 13875 40069
rect 14921 40103 14979 40109
rect 14921 40069 14933 40103
rect 14967 40100 14979 40103
rect 15749 40103 15807 40109
rect 15749 40100 15761 40103
rect 14967 40072 15761 40100
rect 14967 40069 14979 40072
rect 14921 40063 14979 40069
rect 15749 40069 15761 40072
rect 15795 40069 15807 40103
rect 15749 40063 15807 40069
rect 16758 40060 16764 40112
rect 16816 40100 16822 40112
rect 17221 40103 17279 40109
rect 17221 40100 17233 40103
rect 16816 40072 17233 40100
rect 16816 40060 16822 40072
rect 17221 40069 17233 40072
rect 17267 40069 17279 40103
rect 17221 40063 17279 40069
rect 17770 40060 17776 40112
rect 17828 40100 17834 40112
rect 18049 40103 18107 40109
rect 18049 40100 18061 40103
rect 17828 40072 18061 40100
rect 17828 40060 17834 40072
rect 18049 40069 18061 40072
rect 18095 40069 18107 40103
rect 18049 40063 18107 40069
rect 18322 40060 18328 40112
rect 18380 40100 18386 40112
rect 19613 40103 19671 40109
rect 19613 40100 19625 40103
rect 18380 40072 19625 40100
rect 18380 40060 18386 40072
rect 19613 40069 19625 40072
rect 19659 40069 19671 40103
rect 19613 40063 19671 40069
rect 10873 40035 10931 40041
rect 10873 40001 10885 40035
rect 10919 40032 10931 40035
rect 11698 40032 11704 40044
rect 10919 40004 11704 40032
rect 10919 40001 10931 40004
rect 10873 39995 10931 40001
rect 11698 39992 11704 40004
rect 11756 39992 11762 40044
rect 15378 40032 15384 40044
rect 14752 40004 15384 40032
rect 10502 39924 10508 39976
rect 10560 39964 10566 39976
rect 14752 39973 14780 40004
rect 15378 39992 15384 40004
rect 15436 39992 15442 40044
rect 17310 39992 17316 40044
rect 17368 39992 17374 40044
rect 20916 40032 20944 40140
rect 21358 40128 21364 40140
rect 21416 40168 21422 40180
rect 22373 40171 22431 40177
rect 22373 40168 22385 40171
rect 21416 40140 22385 40168
rect 21416 40128 21422 40140
rect 22373 40137 22385 40140
rect 22419 40137 22431 40171
rect 22373 40131 22431 40137
rect 22741 40171 22799 40177
rect 22741 40137 22753 40171
rect 22787 40168 22799 40171
rect 24946 40168 24952 40180
rect 22787 40140 24952 40168
rect 22787 40137 22799 40140
rect 22741 40131 22799 40137
rect 24946 40128 24952 40140
rect 25004 40128 25010 40180
rect 20990 40060 20996 40112
rect 21048 40100 21054 40112
rect 21910 40100 21916 40112
rect 21048 40072 21916 40100
rect 21048 40060 21054 40072
rect 21910 40060 21916 40072
rect 21968 40100 21974 40112
rect 24762 40100 24768 40112
rect 21968 40072 23612 40100
rect 24610 40072 24768 40100
rect 21968 40060 21974 40072
rect 21177 40035 21235 40041
rect 21177 40032 21189 40035
rect 17420 40004 21189 40032
rect 10597 39967 10655 39973
rect 10597 39964 10609 39967
rect 10560 39936 10609 39964
rect 10560 39924 10566 39936
rect 10597 39933 10609 39936
rect 10643 39933 10655 39967
rect 10597 39927 10655 39933
rect 14737 39967 14795 39973
rect 14737 39933 14749 39967
rect 14783 39933 14795 39967
rect 14737 39927 14795 39933
rect 14826 39924 14832 39976
rect 14884 39924 14890 39976
rect 15930 39924 15936 39976
rect 15988 39964 15994 39976
rect 17420 39964 17448 40004
rect 21177 40001 21189 40004
rect 21223 40001 21235 40035
rect 21177 39995 21235 40001
rect 21453 40035 21511 40041
rect 21453 40001 21465 40035
rect 21499 40032 21511 40035
rect 22186 40032 22192 40044
rect 21499 40004 22192 40032
rect 21499 40001 21511 40004
rect 21453 39995 21511 40001
rect 22186 39992 22192 40004
rect 22244 39992 22250 40044
rect 15988 39936 17448 39964
rect 17497 39967 17555 39973
rect 15988 39924 15994 39936
rect 17497 39933 17509 39967
rect 17543 39933 17555 39967
rect 17497 39927 17555 39933
rect 17512 39896 17540 39927
rect 18874 39924 18880 39976
rect 18932 39964 18938 39976
rect 19337 39967 19395 39973
rect 19337 39964 19349 39967
rect 18932 39936 19349 39964
rect 18932 39924 18938 39936
rect 19337 39933 19349 39936
rect 19383 39933 19395 39967
rect 19337 39927 19395 39933
rect 21634 39924 21640 39976
rect 21692 39964 21698 39976
rect 22002 39964 22008 39976
rect 21692 39936 22008 39964
rect 21692 39924 21698 39936
rect 22002 39924 22008 39936
rect 22060 39924 22066 39976
rect 23584 39973 23612 40072
rect 24762 40060 24768 40072
rect 24820 40060 24826 40112
rect 25314 39992 25320 40044
rect 25372 39992 25378 40044
rect 22097 39967 22155 39973
rect 22097 39933 22109 39967
rect 22143 39964 22155 39967
rect 22281 39967 22339 39973
rect 22143 39936 22232 39964
rect 22143 39933 22155 39936
rect 22097 39927 22155 39933
rect 22204 39908 22232 39936
rect 22281 39933 22293 39967
rect 22327 39933 22339 39967
rect 22281 39927 22339 39933
rect 23569 39967 23627 39973
rect 23569 39933 23581 39967
rect 23615 39933 23627 39967
rect 23569 39927 23627 39933
rect 13372 39868 17540 39896
rect 6638 39788 6644 39840
rect 6696 39828 6702 39840
rect 8570 39828 8576 39840
rect 6696 39800 8576 39828
rect 6696 39788 6702 39800
rect 8570 39788 8576 39800
rect 8628 39828 8634 39840
rect 10962 39828 10968 39840
rect 8628 39800 10968 39828
rect 8628 39788 8634 39800
rect 10962 39788 10968 39800
rect 11020 39788 11026 39840
rect 11238 39788 11244 39840
rect 11296 39788 11302 39840
rect 11514 39788 11520 39840
rect 11572 39828 11578 39840
rect 13372 39828 13400 39868
rect 17678 39856 17684 39908
rect 17736 39896 17742 39908
rect 21545 39899 21603 39905
rect 21545 39896 21557 39899
rect 17736 39868 21557 39896
rect 17736 39856 17742 39868
rect 21545 39865 21557 39868
rect 21591 39896 21603 39899
rect 21591 39868 22094 39896
rect 21591 39865 21603 39868
rect 21545 39859 21603 39865
rect 11572 39800 13400 39828
rect 11572 39788 11578 39800
rect 13446 39788 13452 39840
rect 13504 39828 13510 39840
rect 14185 39831 14243 39837
rect 14185 39828 14197 39831
rect 13504 39800 14197 39828
rect 13504 39788 13510 39800
rect 14185 39797 14197 39800
rect 14231 39828 14243 39831
rect 14826 39828 14832 39840
rect 14231 39800 14832 39828
rect 14231 39797 14243 39800
rect 14185 39791 14243 39797
rect 14826 39788 14832 39800
rect 14884 39788 14890 39840
rect 14918 39788 14924 39840
rect 14976 39828 14982 39840
rect 16301 39831 16359 39837
rect 16301 39828 16313 39831
rect 14976 39800 16313 39828
rect 14976 39788 14982 39800
rect 16301 39797 16313 39800
rect 16347 39828 16359 39831
rect 16942 39828 16948 39840
rect 16347 39800 16948 39828
rect 16347 39797 16359 39800
rect 16301 39791 16359 39797
rect 16942 39788 16948 39800
rect 17000 39788 17006 39840
rect 20254 39788 20260 39840
rect 20312 39788 20318 39840
rect 22066 39828 22094 39868
rect 22186 39856 22192 39908
rect 22244 39856 22250 39908
rect 22296 39828 22324 39927
rect 25038 39924 25044 39976
rect 25096 39924 25102 39976
rect 22066 39800 22324 39828
rect 22554 39788 22560 39840
rect 22612 39828 22618 39840
rect 23109 39831 23167 39837
rect 23109 39828 23121 39831
rect 22612 39800 23121 39828
rect 22612 39788 22618 39800
rect 23109 39797 23121 39800
rect 23155 39828 23167 39831
rect 23566 39828 23572 39840
rect 23155 39800 23572 39828
rect 23155 39797 23167 39800
rect 23109 39791 23167 39797
rect 23566 39788 23572 39800
rect 23624 39788 23630 39840
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 7190 39584 7196 39636
rect 7248 39584 7254 39636
rect 7558 39584 7564 39636
rect 7616 39584 7622 39636
rect 9122 39584 9128 39636
rect 9180 39584 9186 39636
rect 10229 39627 10287 39633
rect 10229 39593 10241 39627
rect 10275 39624 10287 39627
rect 11238 39624 11244 39636
rect 10275 39596 11244 39624
rect 10275 39593 10287 39596
rect 10229 39587 10287 39593
rect 11238 39584 11244 39596
rect 11296 39584 11302 39636
rect 11517 39627 11575 39633
rect 11517 39593 11529 39627
rect 11563 39624 11575 39627
rect 12342 39624 12348 39636
rect 11563 39596 12348 39624
rect 11563 39593 11575 39596
rect 11517 39587 11575 39593
rect 12342 39584 12348 39596
rect 12400 39584 12406 39636
rect 15562 39624 15568 39636
rect 12636 39596 15568 39624
rect 11885 39559 11943 39565
rect 11885 39525 11897 39559
rect 11931 39556 11943 39559
rect 12434 39556 12440 39568
rect 11931 39528 12440 39556
rect 11931 39525 11943 39528
rect 11885 39519 11943 39525
rect 12434 39516 12440 39528
rect 12492 39516 12498 39568
rect 12636 39556 12664 39596
rect 15562 39584 15568 39596
rect 15620 39584 15626 39636
rect 17129 39627 17187 39633
rect 17129 39593 17141 39627
rect 17175 39624 17187 39627
rect 18598 39624 18604 39636
rect 17175 39596 18604 39624
rect 17175 39593 17187 39596
rect 17129 39587 17187 39593
rect 18598 39584 18604 39596
rect 18656 39584 18662 39636
rect 20254 39584 20260 39636
rect 20312 39584 20318 39636
rect 25038 39584 25044 39636
rect 25096 39624 25102 39636
rect 25317 39627 25375 39633
rect 25317 39624 25329 39627
rect 25096 39596 25329 39624
rect 25096 39584 25102 39596
rect 25317 39593 25329 39596
rect 25363 39593 25375 39627
rect 25317 39587 25375 39593
rect 12544 39528 12664 39556
rect 8294 39448 8300 39500
rect 8352 39488 8358 39500
rect 9677 39491 9735 39497
rect 9677 39488 9689 39491
rect 8352 39460 9689 39488
rect 8352 39448 8358 39460
rect 9677 39457 9689 39460
rect 9723 39457 9735 39491
rect 9677 39451 9735 39457
rect 10965 39491 11023 39497
rect 10965 39457 10977 39491
rect 11011 39488 11023 39491
rect 11514 39488 11520 39500
rect 11011 39460 11520 39488
rect 11011 39457 11023 39460
rect 10965 39451 11023 39457
rect 11514 39448 11520 39460
rect 11572 39448 11578 39500
rect 11974 39448 11980 39500
rect 12032 39488 12038 39500
rect 12544 39488 12572 39528
rect 12710 39516 12716 39568
rect 12768 39516 12774 39568
rect 14090 39516 14096 39568
rect 14148 39556 14154 39568
rect 15105 39559 15163 39565
rect 15105 39556 15117 39559
rect 14148 39528 15117 39556
rect 14148 39516 14154 39528
rect 15105 39525 15117 39528
rect 15151 39525 15163 39559
rect 15105 39519 15163 39525
rect 16666 39516 16672 39568
rect 16724 39556 16730 39568
rect 17862 39556 17868 39568
rect 16724 39528 17868 39556
rect 16724 39516 16730 39528
rect 17862 39516 17868 39528
rect 17920 39556 17926 39568
rect 18693 39559 18751 39565
rect 18693 39556 18705 39559
rect 17920 39528 18705 39556
rect 17920 39516 17926 39528
rect 18693 39525 18705 39528
rect 18739 39525 18751 39559
rect 20272 39556 20300 39584
rect 20272 39528 20484 39556
rect 18693 39519 18751 39525
rect 12032 39460 12572 39488
rect 12032 39448 12038 39460
rect 5442 39380 5448 39432
rect 5500 39380 5506 39432
rect 9582 39380 9588 39432
rect 9640 39380 9646 39432
rect 11146 39380 11152 39432
rect 11204 39380 11210 39432
rect 12728 39429 12756 39516
rect 12897 39491 12955 39497
rect 12897 39457 12909 39491
rect 12943 39488 12955 39491
rect 12986 39488 12992 39500
rect 12943 39460 12992 39488
rect 12943 39457 12955 39460
rect 12897 39451 12955 39457
rect 12986 39448 12992 39460
rect 13044 39448 13050 39500
rect 15749 39491 15807 39497
rect 15749 39457 15761 39491
rect 15795 39488 15807 39491
rect 16482 39488 16488 39500
rect 15795 39460 16488 39488
rect 15795 39457 15807 39460
rect 15749 39451 15807 39457
rect 16482 39448 16488 39460
rect 16540 39448 16546 39500
rect 16577 39491 16635 39497
rect 16577 39457 16589 39491
rect 16623 39488 16635 39491
rect 17126 39488 17132 39500
rect 16623 39460 17132 39488
rect 16623 39457 16635 39460
rect 16577 39451 16635 39457
rect 17126 39448 17132 39460
rect 17184 39448 17190 39500
rect 19426 39488 19432 39500
rect 17236 39460 19432 39488
rect 12713 39423 12771 39429
rect 12713 39389 12725 39423
rect 12759 39389 12771 39423
rect 12713 39383 12771 39389
rect 15562 39380 15568 39432
rect 15620 39420 15626 39432
rect 17236 39420 17264 39460
rect 19426 39448 19432 39460
rect 19484 39448 19490 39500
rect 20254 39448 20260 39500
rect 20312 39448 20318 39500
rect 20456 39497 20484 39528
rect 22278 39516 22284 39568
rect 22336 39556 22342 39568
rect 22646 39556 22652 39568
rect 22336 39528 22652 39556
rect 22336 39516 22342 39528
rect 22646 39516 22652 39528
rect 22704 39516 22710 39568
rect 20441 39491 20499 39497
rect 20441 39457 20453 39491
rect 20487 39457 20499 39491
rect 20441 39451 20499 39457
rect 23750 39448 23756 39500
rect 23808 39488 23814 39500
rect 24029 39491 24087 39497
rect 24029 39488 24041 39491
rect 23808 39460 24041 39488
rect 23808 39448 23814 39460
rect 24029 39457 24041 39460
rect 24075 39457 24087 39491
rect 24029 39451 24087 39457
rect 15620 39392 17264 39420
rect 15620 39380 15626 39392
rect 17402 39380 17408 39432
rect 17460 39420 17466 39432
rect 17773 39423 17831 39429
rect 17773 39420 17785 39423
rect 17460 39392 17785 39420
rect 17460 39380 17466 39392
rect 17773 39389 17785 39392
rect 17819 39389 17831 39423
rect 17773 39383 17831 39389
rect 20533 39423 20591 39429
rect 20533 39389 20545 39423
rect 20579 39420 20591 39423
rect 21174 39420 21180 39432
rect 20579 39392 21180 39420
rect 20579 39389 20591 39392
rect 20533 39383 20591 39389
rect 21174 39380 21180 39392
rect 21232 39380 21238 39432
rect 21634 39380 21640 39432
rect 21692 39380 21698 39432
rect 24670 39380 24676 39432
rect 24728 39380 24734 39432
rect 5350 39312 5356 39364
rect 5408 39352 5414 39364
rect 5721 39355 5779 39361
rect 5721 39352 5733 39355
rect 5408 39324 5733 39352
rect 5408 39312 5414 39324
rect 5721 39321 5733 39324
rect 5767 39321 5779 39355
rect 7558 39352 7564 39364
rect 6946 39324 7564 39352
rect 5721 39315 5779 39321
rect 7558 39312 7564 39324
rect 7616 39312 7622 39364
rect 9600 39352 9628 39380
rect 12621 39355 12679 39361
rect 9600 39324 12296 39352
rect 8573 39287 8631 39293
rect 8573 39253 8585 39287
rect 8619 39284 8631 39287
rect 8754 39284 8760 39296
rect 8619 39256 8760 39284
rect 8619 39253 8631 39256
rect 8573 39247 8631 39253
rect 8754 39244 8760 39256
rect 8812 39244 8818 39296
rect 9490 39244 9496 39296
rect 9548 39244 9554 39296
rect 9582 39244 9588 39296
rect 9640 39244 9646 39296
rect 10505 39287 10563 39293
rect 10505 39253 10517 39287
rect 10551 39284 10563 39287
rect 11057 39287 11115 39293
rect 11057 39284 11069 39287
rect 10551 39256 11069 39284
rect 10551 39253 10563 39256
rect 10505 39247 10563 39253
rect 11057 39253 11069 39256
rect 11103 39284 11115 39287
rect 11330 39284 11336 39296
rect 11103 39256 11336 39284
rect 11103 39253 11115 39256
rect 11057 39247 11115 39253
rect 11330 39244 11336 39256
rect 11388 39244 11394 39296
rect 12268 39293 12296 39324
rect 12621 39321 12633 39355
rect 12667 39352 12679 39355
rect 16761 39355 16819 39361
rect 12667 39324 12848 39352
rect 12667 39321 12679 39324
rect 12621 39315 12679 39321
rect 12253 39287 12311 39293
rect 12253 39253 12265 39287
rect 12299 39253 12311 39287
rect 12820 39284 12848 39324
rect 16761 39321 16773 39355
rect 16807 39352 16819 39355
rect 19429 39355 19487 39361
rect 19429 39352 19441 39355
rect 16807 39324 19441 39352
rect 16807 39321 16819 39324
rect 16761 39315 16819 39321
rect 19429 39321 19441 39324
rect 19475 39321 19487 39355
rect 21652 39352 21680 39380
rect 23753 39355 23811 39361
rect 19429 39315 19487 39321
rect 19536 39324 21680 39352
rect 23322 39324 23428 39352
rect 13262 39284 13268 39296
rect 12820 39256 13268 39284
rect 12253 39247 12311 39253
rect 13262 39244 13268 39256
rect 13320 39244 13326 39296
rect 15470 39244 15476 39296
rect 15528 39244 15534 39296
rect 15562 39244 15568 39296
rect 15620 39244 15626 39296
rect 16298 39244 16304 39296
rect 16356 39284 16362 39296
rect 16669 39287 16727 39293
rect 16669 39284 16681 39287
rect 16356 39256 16681 39284
rect 16356 39244 16362 39256
rect 16669 39253 16681 39256
rect 16715 39253 16727 39287
rect 16669 39247 16727 39253
rect 18414 39244 18420 39296
rect 18472 39244 18478 39296
rect 18598 39244 18604 39296
rect 18656 39284 18662 39296
rect 19536 39284 19564 39324
rect 18656 39256 19564 39284
rect 18656 39244 18662 39256
rect 20898 39244 20904 39296
rect 20956 39244 20962 39296
rect 21637 39287 21695 39293
rect 21637 39253 21649 39287
rect 21683 39284 21695 39287
rect 22186 39284 22192 39296
rect 21683 39256 22192 39284
rect 21683 39253 21695 39256
rect 21637 39247 21695 39253
rect 22186 39244 22192 39256
rect 22244 39244 22250 39296
rect 22278 39244 22284 39296
rect 22336 39244 22342 39296
rect 23400 39284 23428 39324
rect 23753 39321 23765 39355
rect 23799 39352 23811 39355
rect 25222 39352 25228 39364
rect 23799 39324 25228 39352
rect 23799 39321 23811 39324
rect 23753 39315 23811 39321
rect 25222 39312 25228 39324
rect 25280 39312 25286 39364
rect 24762 39284 24768 39296
rect 23400 39256 24768 39284
rect 24762 39244 24768 39256
rect 24820 39244 24826 39296
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 5350 39040 5356 39092
rect 5408 39040 5414 39092
rect 5902 39040 5908 39092
rect 5960 39080 5966 39092
rect 6549 39083 6607 39089
rect 6549 39080 6561 39083
rect 5960 39052 6561 39080
rect 5960 39040 5966 39052
rect 6549 39049 6561 39052
rect 6595 39049 6607 39083
rect 6549 39043 6607 39049
rect 7374 39040 7380 39092
rect 7432 39080 7438 39092
rect 8021 39083 8079 39089
rect 8021 39080 8033 39083
rect 7432 39052 8033 39080
rect 7432 39040 7438 39052
rect 8021 39049 8033 39052
rect 8067 39080 8079 39083
rect 8665 39083 8723 39089
rect 8665 39080 8677 39083
rect 8067 39052 8677 39080
rect 8067 39049 8079 39052
rect 8021 39043 8079 39049
rect 8665 39049 8677 39052
rect 8711 39049 8723 39083
rect 8665 39043 8723 39049
rect 8680 39012 8708 39043
rect 8754 39040 8760 39092
rect 8812 39040 8818 39092
rect 9125 39083 9183 39089
rect 9125 39049 9137 39083
rect 9171 39080 9183 39083
rect 9398 39080 9404 39092
rect 9171 39052 9404 39080
rect 9171 39049 9183 39052
rect 9125 39043 9183 39049
rect 9398 39040 9404 39052
rect 9456 39040 9462 39092
rect 9582 39040 9588 39092
rect 9640 39080 9646 39092
rect 10413 39083 10471 39089
rect 10413 39080 10425 39083
rect 9640 39052 10425 39080
rect 9640 39040 9646 39052
rect 10413 39049 10425 39052
rect 10459 39049 10471 39083
rect 12434 39080 12440 39092
rect 10413 39043 10471 39049
rect 10520 39052 12440 39080
rect 10520 39012 10548 39052
rect 12434 39040 12440 39052
rect 12492 39040 12498 39092
rect 17405 39083 17463 39089
rect 17405 39080 17417 39083
rect 12544 39052 17417 39080
rect 6012 38984 7144 39012
rect 8680 38984 10548 39012
rect 10781 39015 10839 39021
rect 6012 38956 6040 38984
rect 5994 38904 6000 38956
rect 6052 38904 6058 38956
rect 6086 38904 6092 38956
rect 6144 38944 6150 38956
rect 6917 38947 6975 38953
rect 6917 38944 6929 38947
rect 6144 38916 6929 38944
rect 6144 38904 6150 38916
rect 6917 38913 6929 38916
rect 6963 38913 6975 38947
rect 6917 38907 6975 38913
rect 7006 38836 7012 38888
rect 7064 38836 7070 38888
rect 7116 38885 7144 38984
rect 10781 38981 10793 39015
rect 10827 39012 10839 39015
rect 12544 39012 12572 39052
rect 17405 39049 17417 39052
rect 17451 39049 17463 39083
rect 17405 39043 17463 39049
rect 17862 39040 17868 39092
rect 17920 39080 17926 39092
rect 19245 39083 19303 39089
rect 19245 39080 19257 39083
rect 17920 39052 19257 39080
rect 17920 39040 17926 39052
rect 19245 39049 19257 39052
rect 19291 39049 19303 39083
rect 19245 39043 19303 39049
rect 20346 39040 20352 39092
rect 20404 39040 20410 39092
rect 23290 39040 23296 39092
rect 23348 39080 23354 39092
rect 23569 39083 23627 39089
rect 23569 39080 23581 39083
rect 23348 39052 23581 39080
rect 23348 39040 23354 39052
rect 23569 39049 23581 39052
rect 23615 39049 23627 39083
rect 23569 39043 23627 39049
rect 23658 39040 23664 39092
rect 23716 39080 23722 39092
rect 23716 39052 25360 39080
rect 23716 39040 23722 39052
rect 13814 39012 13820 39024
rect 10827 38984 12572 39012
rect 13478 38984 13820 39012
rect 10827 38981 10839 38984
rect 10781 38975 10839 38981
rect 13814 38972 13820 38984
rect 13872 38972 13878 39024
rect 13906 38972 13912 39024
rect 13964 38972 13970 39024
rect 15381 39015 15439 39021
rect 15381 38981 15393 39015
rect 15427 39012 15439 39015
rect 17310 39012 17316 39024
rect 15427 38984 17316 39012
rect 15427 38981 15439 38984
rect 15381 38975 15439 38981
rect 17310 38972 17316 38984
rect 17368 38972 17374 39024
rect 17773 39015 17831 39021
rect 17773 38981 17785 39015
rect 17819 39012 17831 39015
rect 18598 39012 18604 39024
rect 17819 38984 18604 39012
rect 17819 38981 17831 38984
rect 17773 38975 17831 38981
rect 18598 38972 18604 38984
rect 18656 38972 18662 39024
rect 20990 39012 20996 39024
rect 19076 38984 20996 39012
rect 10318 38904 10324 38956
rect 10376 38944 10382 38956
rect 10873 38947 10931 38953
rect 10873 38944 10885 38947
rect 10376 38916 10885 38944
rect 10376 38904 10382 38916
rect 10873 38913 10885 38916
rect 10919 38913 10931 38947
rect 10873 38907 10931 38913
rect 14182 38904 14188 38956
rect 14240 38904 14246 38956
rect 15473 38947 15531 38953
rect 15473 38913 15485 38947
rect 15519 38944 15531 38947
rect 15654 38944 15660 38956
rect 15519 38916 15660 38944
rect 15519 38913 15531 38916
rect 15473 38907 15531 38913
rect 15654 38904 15660 38916
rect 15712 38944 15718 38956
rect 16025 38947 16083 38953
rect 16025 38944 16037 38947
rect 15712 38916 16037 38944
rect 15712 38904 15718 38916
rect 16025 38913 16037 38916
rect 16071 38913 16083 38947
rect 16025 38907 16083 38913
rect 17865 38947 17923 38953
rect 17865 38913 17877 38947
rect 17911 38944 17923 38947
rect 18417 38947 18475 38953
rect 18417 38944 18429 38947
rect 17911 38916 18429 38944
rect 17911 38913 17923 38916
rect 17865 38907 17923 38913
rect 18417 38913 18429 38916
rect 18463 38913 18475 38947
rect 18417 38907 18475 38913
rect 7101 38879 7159 38885
rect 7101 38845 7113 38879
rect 7147 38845 7159 38879
rect 7101 38839 7159 38845
rect 8570 38836 8576 38888
rect 8628 38836 8634 38888
rect 9950 38836 9956 38888
rect 10008 38836 10014 38888
rect 10042 38836 10048 38888
rect 10100 38876 10106 38888
rect 10965 38879 11023 38885
rect 10965 38876 10977 38879
rect 10100 38848 10977 38876
rect 10100 38836 10106 38848
rect 10965 38845 10977 38848
rect 11011 38845 11023 38879
rect 10965 38839 11023 38845
rect 11698 38836 11704 38888
rect 11756 38836 11762 38888
rect 15565 38879 15623 38885
rect 12912 38848 14228 38876
rect 9030 38768 9036 38820
rect 9088 38808 9094 38820
rect 12342 38808 12348 38820
rect 9088 38780 12348 38808
rect 9088 38768 9094 38780
rect 12342 38768 12348 38780
rect 12400 38768 12406 38820
rect 12437 38811 12495 38817
rect 12437 38777 12449 38811
rect 12483 38808 12495 38811
rect 12618 38808 12624 38820
rect 12483 38780 12624 38808
rect 12483 38777 12495 38780
rect 12437 38771 12495 38777
rect 12618 38768 12624 38780
rect 12676 38768 12682 38820
rect 9674 38700 9680 38752
rect 9732 38740 9738 38752
rect 12912 38740 12940 38848
rect 14200 38820 14228 38848
rect 15565 38845 15577 38879
rect 15611 38876 15623 38879
rect 15838 38876 15844 38888
rect 15611 38848 15844 38876
rect 15611 38845 15623 38848
rect 15565 38839 15623 38845
rect 15838 38836 15844 38848
rect 15896 38836 15902 38888
rect 17957 38879 18015 38885
rect 17957 38845 17969 38879
rect 18003 38845 18015 38879
rect 17957 38839 18015 38845
rect 14182 38768 14188 38820
rect 14240 38808 14246 38820
rect 14240 38780 15148 38808
rect 14240 38768 14246 38780
rect 9732 38712 12940 38740
rect 9732 38700 9738 38712
rect 13262 38700 13268 38752
rect 13320 38740 13326 38752
rect 13446 38740 13452 38752
rect 13320 38712 13452 38740
rect 13320 38700 13326 38712
rect 13446 38700 13452 38712
rect 13504 38700 13510 38752
rect 13814 38700 13820 38752
rect 13872 38740 13878 38752
rect 14461 38743 14519 38749
rect 14461 38740 14473 38743
rect 13872 38712 14473 38740
rect 13872 38700 13878 38712
rect 14461 38709 14473 38712
rect 14507 38709 14519 38743
rect 14461 38703 14519 38709
rect 14550 38700 14556 38752
rect 14608 38740 14614 38752
rect 15013 38743 15071 38749
rect 15013 38740 15025 38743
rect 14608 38712 15025 38740
rect 14608 38700 14614 38712
rect 15013 38709 15025 38712
rect 15059 38709 15071 38743
rect 15120 38740 15148 38780
rect 15378 38768 15384 38820
rect 15436 38808 15442 38820
rect 17037 38811 17095 38817
rect 17037 38808 17049 38811
rect 15436 38780 17049 38808
rect 15436 38768 15442 38780
rect 17037 38777 17049 38780
rect 17083 38808 17095 38811
rect 17972 38808 18000 38839
rect 17083 38780 18000 38808
rect 17083 38777 17095 38780
rect 17037 38771 17095 38777
rect 16209 38743 16267 38749
rect 16209 38740 16221 38743
rect 15120 38712 16221 38740
rect 15013 38703 15071 38709
rect 16209 38709 16221 38712
rect 16255 38740 16267 38743
rect 16298 38740 16304 38752
rect 16255 38712 16304 38740
rect 16255 38709 16267 38712
rect 16209 38703 16267 38709
rect 16298 38700 16304 38712
rect 16356 38700 16362 38752
rect 16666 38700 16672 38752
rect 16724 38740 16730 38752
rect 17678 38740 17684 38752
rect 16724 38712 17684 38740
rect 16724 38700 16730 38712
rect 17678 38700 17684 38712
rect 17736 38700 17742 38752
rect 18432 38740 18460 38907
rect 19076 38885 19104 38984
rect 20990 38972 20996 38984
rect 21048 38972 21054 39024
rect 22373 39015 22431 39021
rect 22373 38981 22385 39015
rect 22419 39012 22431 39015
rect 22462 39012 22468 39024
rect 22419 38984 22468 39012
rect 22419 38981 22431 38984
rect 22373 38975 22431 38981
rect 22462 38972 22468 38984
rect 22520 38972 22526 39024
rect 23477 39015 23535 39021
rect 23477 38981 23489 39015
rect 23523 39012 23535 39015
rect 24578 39012 24584 39024
rect 23523 38984 24584 39012
rect 23523 38981 23535 38984
rect 23477 38975 23535 38981
rect 24578 38972 24584 38984
rect 24636 38972 24642 39024
rect 25332 39021 25360 39052
rect 25317 39015 25375 39021
rect 25317 38981 25329 39015
rect 25363 38981 25375 39015
rect 25317 38975 25375 38981
rect 19702 38904 19708 38956
rect 19760 38944 19766 38956
rect 20441 38947 20499 38953
rect 20441 38944 20453 38947
rect 19760 38916 20453 38944
rect 19760 38904 19766 38916
rect 20441 38913 20453 38916
rect 20487 38913 20499 38947
rect 20441 38907 20499 38913
rect 21453 38947 21511 38953
rect 21453 38913 21465 38947
rect 21499 38944 21511 38947
rect 22186 38944 22192 38956
rect 21499 38916 22192 38944
rect 21499 38913 21511 38916
rect 21453 38907 21511 38913
rect 22186 38904 22192 38916
rect 22244 38904 22250 38956
rect 24302 38944 24308 38956
rect 22664 38916 24308 38944
rect 19061 38879 19119 38885
rect 19061 38845 19073 38879
rect 19107 38845 19119 38879
rect 19061 38839 19119 38845
rect 19153 38879 19211 38885
rect 19153 38845 19165 38879
rect 19199 38845 19211 38879
rect 19153 38839 19211 38845
rect 18874 38768 18880 38820
rect 18932 38808 18938 38820
rect 19168 38808 19196 38839
rect 20162 38836 20168 38888
rect 20220 38836 20226 38888
rect 20714 38836 20720 38888
rect 20772 38876 20778 38888
rect 21818 38876 21824 38888
rect 20772 38848 21824 38876
rect 20772 38836 20778 38848
rect 21818 38836 21824 38848
rect 21876 38876 21882 38888
rect 22465 38879 22523 38885
rect 21876 38848 22094 38876
rect 21876 38836 21882 38848
rect 18932 38780 19196 38808
rect 19613 38811 19671 38817
rect 18932 38768 18938 38780
rect 19613 38777 19625 38811
rect 19659 38808 19671 38811
rect 21542 38808 21548 38820
rect 19659 38780 21548 38808
rect 19659 38777 19671 38780
rect 19613 38771 19671 38777
rect 21542 38768 21548 38780
rect 21600 38768 21606 38820
rect 22066 38808 22094 38848
rect 22465 38845 22477 38879
rect 22511 38876 22523 38879
rect 22554 38876 22560 38888
rect 22511 38848 22560 38876
rect 22511 38845 22523 38848
rect 22465 38839 22523 38845
rect 22554 38836 22560 38848
rect 22612 38836 22618 38888
rect 22664 38885 22692 38916
rect 24302 38904 24308 38916
rect 24360 38904 24366 38956
rect 22649 38879 22707 38885
rect 22649 38845 22661 38879
rect 22695 38845 22707 38879
rect 22649 38839 22707 38845
rect 23385 38879 23443 38885
rect 23385 38845 23397 38879
rect 23431 38876 23443 38879
rect 24026 38876 24032 38888
rect 23431 38848 24032 38876
rect 23431 38845 23443 38848
rect 23385 38839 23443 38845
rect 24026 38836 24032 38848
rect 24084 38836 24090 38888
rect 24581 38879 24639 38885
rect 24581 38845 24593 38879
rect 24627 38876 24639 38879
rect 24762 38876 24768 38888
rect 24627 38848 24768 38876
rect 24627 38845 24639 38848
rect 24581 38839 24639 38845
rect 24762 38836 24768 38848
rect 24820 38836 24826 38888
rect 25866 38808 25872 38820
rect 22066 38780 25872 38808
rect 25866 38768 25872 38780
rect 25924 38768 25930 38820
rect 20714 38740 20720 38752
rect 18432 38712 20720 38740
rect 20714 38700 20720 38712
rect 20772 38700 20778 38752
rect 20806 38700 20812 38752
rect 20864 38700 20870 38752
rect 20990 38700 20996 38752
rect 21048 38740 21054 38752
rect 21269 38743 21327 38749
rect 21269 38740 21281 38743
rect 21048 38712 21281 38740
rect 21048 38700 21054 38712
rect 21269 38709 21281 38712
rect 21315 38709 21327 38743
rect 21269 38703 21327 38709
rect 22002 38700 22008 38752
rect 22060 38700 22066 38752
rect 22462 38700 22468 38752
rect 22520 38740 22526 38752
rect 23566 38740 23572 38752
rect 22520 38712 23572 38740
rect 22520 38700 22526 38712
rect 23566 38700 23572 38712
rect 23624 38700 23630 38752
rect 23937 38743 23995 38749
rect 23937 38709 23949 38743
rect 23983 38740 23995 38743
rect 24302 38740 24308 38752
rect 23983 38712 24308 38740
rect 23983 38709 23995 38712
rect 23937 38703 23995 38709
rect 24302 38700 24308 38712
rect 24360 38700 24366 38752
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 10505 38539 10563 38545
rect 10505 38505 10517 38539
rect 10551 38536 10563 38539
rect 10686 38536 10692 38548
rect 10551 38508 10692 38536
rect 10551 38505 10563 38508
rect 10505 38499 10563 38505
rect 10686 38496 10692 38508
rect 10744 38496 10750 38548
rect 11701 38539 11759 38545
rect 11701 38505 11713 38539
rect 11747 38536 11759 38539
rect 11790 38536 11796 38548
rect 11747 38508 11796 38536
rect 11747 38505 11759 38508
rect 11701 38499 11759 38505
rect 11790 38496 11796 38508
rect 11848 38496 11854 38548
rect 18141 38539 18199 38545
rect 11900 38508 17724 38536
rect 8478 38428 8484 38480
rect 8536 38468 8542 38480
rect 8536 38440 11008 38468
rect 8536 38428 8542 38440
rect 5442 38360 5448 38412
rect 5500 38400 5506 38412
rect 5629 38403 5687 38409
rect 5629 38400 5641 38403
rect 5500 38372 5641 38400
rect 5500 38360 5506 38372
rect 5629 38369 5641 38372
rect 5675 38400 5687 38403
rect 6546 38400 6552 38412
rect 5675 38372 6552 38400
rect 5675 38369 5687 38372
rect 5629 38363 5687 38369
rect 6546 38360 6552 38372
rect 6604 38360 6610 38412
rect 6638 38360 6644 38412
rect 6696 38400 6702 38412
rect 7377 38403 7435 38409
rect 6696 38372 7236 38400
rect 6696 38360 6702 38372
rect 1302 38292 1308 38344
rect 1360 38332 1366 38344
rect 1581 38335 1639 38341
rect 1581 38332 1593 38335
rect 1360 38304 1593 38332
rect 1360 38292 1366 38304
rect 1581 38301 1593 38304
rect 1627 38332 1639 38335
rect 2041 38335 2099 38341
rect 2041 38332 2053 38335
rect 1627 38304 2053 38332
rect 1627 38301 1639 38304
rect 1581 38295 1639 38301
rect 2041 38301 2053 38304
rect 2087 38301 2099 38335
rect 2041 38295 2099 38301
rect 5905 38267 5963 38273
rect 5905 38233 5917 38267
rect 5951 38233 5963 38267
rect 5905 38227 5963 38233
rect 1765 38199 1823 38205
rect 1765 38165 1777 38199
rect 1811 38196 1823 38199
rect 4062 38196 4068 38208
rect 1811 38168 4068 38196
rect 1811 38165 1823 38168
rect 1765 38159 1823 38165
rect 4062 38156 4068 38168
rect 4120 38156 4126 38208
rect 5920 38196 5948 38227
rect 6362 38224 6368 38276
rect 6420 38224 6426 38276
rect 7208 38264 7236 38372
rect 7377 38369 7389 38403
rect 7423 38369 7435 38403
rect 7377 38363 7435 38369
rect 9861 38403 9919 38409
rect 9861 38369 9873 38403
rect 9907 38369 9919 38403
rect 9861 38363 9919 38369
rect 7392 38332 7420 38363
rect 7837 38335 7895 38341
rect 7837 38332 7849 38335
rect 7392 38304 7849 38332
rect 7837 38301 7849 38304
rect 7883 38332 7895 38335
rect 8294 38332 8300 38344
rect 7883 38304 8300 38332
rect 7883 38301 7895 38304
rect 7837 38295 7895 38301
rect 8294 38292 8300 38304
rect 8352 38292 8358 38344
rect 9493 38335 9551 38341
rect 9493 38301 9505 38335
rect 9539 38332 9551 38335
rect 9876 38332 9904 38363
rect 9539 38304 9904 38332
rect 9539 38301 9551 38304
rect 9493 38295 9551 38301
rect 9876 38264 9904 38304
rect 9950 38292 9956 38344
rect 10008 38332 10014 38344
rect 10137 38335 10195 38341
rect 10137 38332 10149 38335
rect 10008 38304 10149 38332
rect 10008 38292 10014 38304
rect 10137 38301 10149 38304
rect 10183 38301 10195 38335
rect 10980 38332 11008 38440
rect 11054 38360 11060 38412
rect 11112 38360 11118 38412
rect 11900 38400 11928 38508
rect 11974 38428 11980 38480
rect 12032 38468 12038 38480
rect 12713 38471 12771 38477
rect 12713 38468 12725 38471
rect 12032 38440 12725 38468
rect 12032 38428 12038 38440
rect 12713 38437 12725 38440
rect 12759 38437 12771 38471
rect 14737 38471 14795 38477
rect 14737 38468 14749 38471
rect 12713 38431 12771 38437
rect 13648 38440 14749 38468
rect 11256 38372 11928 38400
rect 11256 38332 11284 38372
rect 12434 38360 12440 38412
rect 12492 38400 12498 38412
rect 13265 38403 13323 38409
rect 13265 38400 13277 38403
rect 12492 38372 13277 38400
rect 12492 38360 12498 38372
rect 13265 38369 13277 38372
rect 13311 38369 13323 38403
rect 13265 38363 13323 38369
rect 10980 38304 11284 38332
rect 11333 38335 11391 38341
rect 10137 38295 10195 38301
rect 11333 38301 11345 38335
rect 11379 38332 11391 38335
rect 11698 38332 11704 38344
rect 11379 38304 11704 38332
rect 11379 38301 11391 38304
rect 11333 38295 11391 38301
rect 11698 38292 11704 38304
rect 11756 38292 11762 38344
rect 13648 38332 13676 38440
rect 14737 38437 14749 38440
rect 14783 38468 14795 38471
rect 16114 38468 16120 38480
rect 14783 38440 16120 38468
rect 14783 38437 14795 38440
rect 14737 38431 14795 38437
rect 16114 38428 16120 38440
rect 16172 38428 16178 38480
rect 16574 38468 16580 38480
rect 16316 38440 16580 38468
rect 13817 38403 13875 38409
rect 13817 38400 13829 38403
rect 11808 38304 13676 38332
rect 13740 38372 13829 38400
rect 11808 38264 11836 38304
rect 7208 38236 9352 38264
rect 9876 38236 11836 38264
rect 12437 38267 12495 38273
rect 7466 38196 7472 38208
rect 5920 38168 7472 38196
rect 7466 38156 7472 38168
rect 7524 38156 7530 38208
rect 8294 38156 8300 38208
rect 8352 38196 8358 38208
rect 9324 38205 9352 38236
rect 12437 38233 12449 38267
rect 12483 38264 12495 38267
rect 12802 38264 12808 38276
rect 12483 38236 12808 38264
rect 12483 38233 12495 38236
rect 12437 38227 12495 38233
rect 12802 38224 12808 38236
rect 12860 38264 12866 38276
rect 13173 38267 13231 38273
rect 13173 38264 13185 38267
rect 12860 38236 13185 38264
rect 12860 38224 12866 38236
rect 13173 38233 13185 38236
rect 13219 38233 13231 38267
rect 13173 38227 13231 38233
rect 8481 38199 8539 38205
rect 8481 38196 8493 38199
rect 8352 38168 8493 38196
rect 8352 38156 8358 38168
rect 8481 38165 8493 38168
rect 8527 38165 8539 38199
rect 8481 38159 8539 38165
rect 9309 38199 9367 38205
rect 9309 38165 9321 38199
rect 9355 38196 9367 38199
rect 9858 38196 9864 38208
rect 9355 38168 9864 38196
rect 9355 38165 9367 38168
rect 9309 38159 9367 38165
rect 9858 38156 9864 38168
rect 9916 38196 9922 38208
rect 10045 38199 10103 38205
rect 10045 38196 10057 38199
rect 9916 38168 10057 38196
rect 9916 38156 9922 38168
rect 10045 38165 10057 38168
rect 10091 38165 10103 38199
rect 10045 38159 10103 38165
rect 11238 38156 11244 38208
rect 11296 38156 11302 38208
rect 13081 38199 13139 38205
rect 13081 38165 13093 38199
rect 13127 38196 13139 38199
rect 13740 38196 13768 38372
rect 13817 38369 13829 38372
rect 13863 38400 13875 38403
rect 15378 38400 15384 38412
rect 13863 38372 15384 38400
rect 13863 38369 13875 38372
rect 13817 38363 13875 38369
rect 15378 38360 15384 38372
rect 15436 38360 15442 38412
rect 15654 38360 15660 38412
rect 15712 38400 15718 38412
rect 15838 38400 15844 38412
rect 15712 38372 15844 38400
rect 15712 38360 15718 38372
rect 15838 38360 15844 38372
rect 15896 38360 15902 38412
rect 16316 38409 16344 38440
rect 16574 38428 16580 38440
rect 16632 38428 16638 38480
rect 16301 38403 16359 38409
rect 16301 38369 16313 38403
rect 16347 38369 16359 38403
rect 16301 38363 16359 38369
rect 16390 38360 16396 38412
rect 16448 38400 16454 38412
rect 17696 38409 17724 38508
rect 18141 38505 18153 38539
rect 18187 38536 18199 38539
rect 18322 38536 18328 38548
rect 18187 38508 18328 38536
rect 18187 38505 18199 38508
rect 18141 38499 18199 38505
rect 18322 38496 18328 38508
rect 18380 38496 18386 38548
rect 19334 38496 19340 38548
rect 19392 38536 19398 38548
rect 19429 38539 19487 38545
rect 19429 38536 19441 38539
rect 19392 38508 19441 38536
rect 19392 38496 19398 38508
rect 19429 38505 19441 38508
rect 19475 38505 19487 38539
rect 19429 38499 19487 38505
rect 23566 38496 23572 38548
rect 23624 38536 23630 38548
rect 24029 38539 24087 38545
rect 24029 38536 24041 38539
rect 23624 38508 24041 38536
rect 23624 38496 23630 38508
rect 24029 38505 24041 38508
rect 24075 38505 24087 38539
rect 24029 38499 24087 38505
rect 24394 38496 24400 38548
rect 24452 38536 24458 38548
rect 24581 38539 24639 38545
rect 24581 38536 24593 38539
rect 24452 38508 24593 38536
rect 24452 38496 24458 38508
rect 24581 38505 24593 38508
rect 24627 38505 24639 38539
rect 24581 38499 24639 38505
rect 18598 38428 18604 38480
rect 18656 38468 18662 38480
rect 21177 38471 21235 38477
rect 21177 38468 21189 38471
rect 18656 38440 21189 38468
rect 18656 38428 18662 38440
rect 21177 38437 21189 38440
rect 21223 38437 21235 38471
rect 21177 38431 21235 38437
rect 21542 38428 21548 38480
rect 21600 38468 21606 38480
rect 22646 38468 22652 38480
rect 21600 38440 22652 38468
rect 21600 38428 21606 38440
rect 22646 38428 22652 38440
rect 22704 38468 22710 38480
rect 22704 38440 25268 38468
rect 22704 38428 22710 38440
rect 16485 38403 16543 38409
rect 16485 38400 16497 38403
rect 16448 38372 16497 38400
rect 16448 38360 16454 38372
rect 16485 38369 16497 38372
rect 16531 38369 16543 38403
rect 16485 38363 16543 38369
rect 17497 38403 17555 38409
rect 17497 38369 17509 38403
rect 17543 38369 17555 38403
rect 17497 38363 17555 38369
rect 17681 38403 17739 38409
rect 17681 38369 17693 38403
rect 17727 38400 17739 38403
rect 18417 38403 18475 38409
rect 18417 38400 18429 38403
rect 17727 38372 18429 38400
rect 17727 38369 17739 38372
rect 17681 38363 17739 38369
rect 18417 38369 18429 38372
rect 18463 38369 18475 38403
rect 18417 38363 18475 38369
rect 14918 38292 14924 38344
rect 14976 38332 14982 38344
rect 17402 38332 17408 38344
rect 14976 38304 17408 38332
rect 14976 38292 14982 38304
rect 17402 38292 17408 38304
rect 17460 38292 17466 38344
rect 13814 38224 13820 38276
rect 13872 38264 13878 38276
rect 16577 38267 16635 38273
rect 16577 38264 16589 38267
rect 13872 38236 16589 38264
rect 13872 38224 13878 38236
rect 16577 38233 16589 38236
rect 16623 38233 16635 38267
rect 17512 38264 17540 38363
rect 19610 38360 19616 38412
rect 19668 38400 19674 38412
rect 19981 38403 20039 38409
rect 19981 38400 19993 38403
rect 19668 38372 19993 38400
rect 19668 38360 19674 38372
rect 19981 38369 19993 38372
rect 20027 38369 20039 38403
rect 19981 38363 20039 38369
rect 20070 38360 20076 38412
rect 20128 38360 20134 38412
rect 21913 38403 21971 38409
rect 21913 38369 21925 38403
rect 21959 38369 21971 38403
rect 21913 38363 21971 38369
rect 17770 38292 17776 38344
rect 17828 38292 17834 38344
rect 18322 38292 18328 38344
rect 18380 38332 18386 38344
rect 18874 38332 18880 38344
rect 18380 38304 18880 38332
rect 18380 38292 18386 38304
rect 18874 38292 18880 38304
rect 18932 38332 18938 38344
rect 18969 38335 19027 38341
rect 18969 38332 18981 38335
rect 18932 38304 18981 38332
rect 18932 38292 18938 38304
rect 18969 38301 18981 38304
rect 19015 38301 19027 38335
rect 18969 38295 19027 38301
rect 19889 38335 19947 38341
rect 19889 38301 19901 38335
rect 19935 38332 19947 38335
rect 20088 38332 20116 38360
rect 19935 38304 20116 38332
rect 19935 38301 19947 38304
rect 19889 38295 19947 38301
rect 21358 38292 21364 38344
rect 21416 38292 21422 38344
rect 19150 38264 19156 38276
rect 17512 38236 19156 38264
rect 16577 38227 16635 38233
rect 19150 38224 19156 38236
rect 19208 38224 19214 38276
rect 19797 38267 19855 38273
rect 19797 38233 19809 38267
rect 19843 38264 19855 38267
rect 20070 38264 20076 38276
rect 19843 38236 20076 38264
rect 19843 38233 19855 38236
rect 19797 38227 19855 38233
rect 20070 38224 20076 38236
rect 20128 38224 20134 38276
rect 20901 38267 20959 38273
rect 20901 38233 20913 38267
rect 20947 38264 20959 38267
rect 21928 38264 21956 38363
rect 22094 38360 22100 38412
rect 22152 38360 22158 38412
rect 23201 38403 23259 38409
rect 23201 38369 23213 38403
rect 23247 38369 23259 38403
rect 23201 38363 23259 38369
rect 23293 38403 23351 38409
rect 23293 38369 23305 38403
rect 23339 38400 23351 38403
rect 23382 38400 23388 38412
rect 23339 38372 23388 38400
rect 23339 38369 23351 38372
rect 23293 38363 23351 38369
rect 22002 38292 22008 38344
rect 22060 38332 22066 38344
rect 22189 38335 22247 38341
rect 22189 38332 22201 38335
rect 22060 38304 22201 38332
rect 22060 38292 22066 38304
rect 22189 38301 22201 38304
rect 22235 38301 22247 38335
rect 23216 38332 23244 38363
rect 23382 38360 23388 38372
rect 23440 38360 23446 38412
rect 25240 38344 25268 38440
rect 24394 38332 24400 38344
rect 23216 38304 24400 38332
rect 22189 38295 22247 38301
rect 24394 38292 24400 38304
rect 24452 38292 24458 38344
rect 25222 38292 25228 38344
rect 25280 38292 25286 38344
rect 22094 38264 22100 38276
rect 20947 38236 21496 38264
rect 21928 38236 22100 38264
rect 20947 38233 20959 38236
rect 20901 38227 20959 38233
rect 13127 38168 13768 38196
rect 13127 38165 13139 38168
rect 13081 38159 13139 38165
rect 14734 38156 14740 38208
rect 14792 38196 14798 38208
rect 15013 38199 15071 38205
rect 15013 38196 15025 38199
rect 14792 38168 15025 38196
rect 14792 38156 14798 38168
rect 15013 38165 15025 38168
rect 15059 38165 15071 38199
rect 15013 38159 15071 38165
rect 15378 38156 15384 38208
rect 15436 38156 15442 38208
rect 15473 38199 15531 38205
rect 15473 38165 15485 38199
rect 15519 38196 15531 38199
rect 16758 38196 16764 38208
rect 15519 38168 16764 38196
rect 15519 38165 15531 38168
rect 15473 38159 15531 38165
rect 16758 38156 16764 38168
rect 16816 38156 16822 38208
rect 16945 38199 17003 38205
rect 16945 38165 16957 38199
rect 16991 38196 17003 38199
rect 17218 38196 17224 38208
rect 16991 38168 17224 38196
rect 16991 38165 17003 38168
rect 16945 38159 17003 38165
rect 17218 38156 17224 38168
rect 17276 38156 17282 38208
rect 17954 38156 17960 38208
rect 18012 38196 18018 38208
rect 18693 38199 18751 38205
rect 18693 38196 18705 38199
rect 18012 38168 18705 38196
rect 18012 38156 18018 38168
rect 18693 38165 18705 38168
rect 18739 38165 18751 38199
rect 18693 38159 18751 38165
rect 20533 38199 20591 38205
rect 20533 38165 20545 38199
rect 20579 38196 20591 38199
rect 20622 38196 20628 38208
rect 20579 38168 20628 38196
rect 20579 38165 20591 38168
rect 20533 38159 20591 38165
rect 20622 38156 20628 38168
rect 20680 38156 20686 38208
rect 21468 38196 21496 38236
rect 22094 38224 22100 38236
rect 22152 38264 22158 38276
rect 22278 38264 22284 38276
rect 22152 38236 22284 38264
rect 22152 38224 22158 38236
rect 22278 38224 22284 38236
rect 22336 38224 22342 38276
rect 22370 38196 22376 38208
rect 21468 38168 22376 38196
rect 22370 38156 22376 38168
rect 22428 38156 22434 38208
rect 22554 38156 22560 38208
rect 22612 38156 22618 38208
rect 23382 38156 23388 38208
rect 23440 38156 23446 38208
rect 23753 38199 23811 38205
rect 23753 38165 23765 38199
rect 23799 38196 23811 38199
rect 23842 38196 23848 38208
rect 23799 38168 23848 38196
rect 23799 38165 23811 38168
rect 23753 38159 23811 38165
rect 23842 38156 23848 38168
rect 23900 38156 23906 38208
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 5442 37992 5448 38004
rect 4264 37964 5448 37992
rect 4264 37865 4292 37964
rect 5442 37952 5448 37964
rect 5500 37952 5506 38004
rect 5994 37952 6000 38004
rect 6052 37952 6058 38004
rect 8846 37992 8852 38004
rect 8220 37964 8852 37992
rect 6362 37924 6368 37936
rect 5750 37896 6368 37924
rect 6362 37884 6368 37896
rect 6420 37884 6426 37936
rect 8220 37924 8248 37964
rect 8846 37952 8852 37964
rect 8904 37952 8910 38004
rect 9953 37995 10011 38001
rect 9953 37961 9965 37995
rect 9999 37992 10011 37995
rect 10410 37992 10416 38004
rect 9999 37964 10416 37992
rect 9999 37961 10011 37964
rect 9953 37955 10011 37961
rect 10410 37952 10416 37964
rect 10468 37952 10474 38004
rect 10594 37952 10600 38004
rect 10652 37952 10658 38004
rect 12069 37995 12127 38001
rect 11164 37964 12020 37992
rect 7866 37896 8248 37924
rect 8294 37884 8300 37936
rect 8352 37884 8358 37936
rect 4249 37859 4307 37865
rect 4249 37825 4261 37859
rect 4295 37825 4307 37859
rect 4249 37819 4307 37825
rect 8662 37816 8668 37868
rect 8720 37816 8726 37868
rect 9861 37859 9919 37865
rect 9861 37825 9873 37859
rect 9907 37856 9919 37859
rect 11164 37856 11192 37964
rect 9907 37828 11192 37856
rect 11992 37856 12020 37964
rect 12069 37961 12081 37995
rect 12115 37992 12127 37995
rect 14734 37992 14740 38004
rect 12115 37964 14740 37992
rect 12115 37961 12127 37964
rect 12069 37955 12127 37961
rect 14734 37952 14740 37964
rect 14792 37952 14798 38004
rect 15378 37952 15384 38004
rect 15436 37992 15442 38004
rect 16117 37995 16175 38001
rect 16117 37992 16129 37995
rect 15436 37964 16129 37992
rect 15436 37952 15442 37964
rect 16117 37961 16129 37964
rect 16163 37961 16175 37995
rect 16117 37955 16175 37961
rect 16482 37952 16488 38004
rect 16540 37992 16546 38004
rect 16850 37992 16856 38004
rect 16540 37964 16856 37992
rect 16540 37952 16546 37964
rect 16850 37952 16856 37964
rect 16908 37952 16914 38004
rect 19061 37995 19119 38001
rect 19061 37992 19073 37995
rect 17052 37964 19073 37992
rect 12161 37927 12219 37933
rect 12161 37893 12173 37927
rect 12207 37924 12219 37927
rect 14550 37924 14556 37936
rect 12207 37896 14556 37924
rect 12207 37893 12219 37896
rect 12161 37887 12219 37893
rect 14550 37884 14556 37896
rect 14608 37884 14614 37936
rect 15028 37896 15424 37924
rect 13541 37859 13599 37865
rect 11992 37828 12434 37856
rect 9907 37825 9919 37828
rect 9861 37819 9919 37825
rect 4525 37791 4583 37797
rect 4525 37757 4537 37791
rect 4571 37788 4583 37791
rect 5534 37788 5540 37800
rect 4571 37760 5540 37788
rect 4571 37757 4583 37760
rect 4525 37751 4583 37757
rect 5534 37748 5540 37760
rect 5592 37748 5598 37800
rect 6549 37791 6607 37797
rect 6549 37757 6561 37791
rect 6595 37788 6607 37791
rect 7098 37788 7104 37800
rect 6595 37760 7104 37788
rect 6595 37757 6607 37760
rect 6549 37751 6607 37757
rect 7098 37748 7104 37760
rect 7156 37748 7162 37800
rect 8570 37748 8576 37800
rect 8628 37748 8634 37800
rect 8680 37720 8708 37816
rect 9582 37748 9588 37800
rect 9640 37788 9646 37800
rect 10045 37791 10103 37797
rect 10045 37788 10057 37791
rect 9640 37760 10057 37788
rect 9640 37748 9646 37760
rect 10045 37757 10057 37760
rect 10091 37757 10103 37791
rect 12253 37791 12311 37797
rect 12253 37788 12265 37791
rect 10045 37751 10103 37757
rect 11256 37760 12265 37788
rect 11256 37729 11284 37760
rect 12253 37757 12265 37760
rect 12299 37757 12311 37791
rect 12406 37788 12434 37828
rect 13541 37825 13553 37859
rect 13587 37856 13599 37859
rect 15028 37856 15056 37896
rect 13587 37828 15056 37856
rect 13587 37825 13599 37828
rect 13541 37819 13599 37825
rect 15194 37816 15200 37868
rect 15252 37856 15258 37868
rect 15289 37859 15347 37865
rect 15289 37856 15301 37859
rect 15252 37828 15301 37856
rect 15252 37816 15258 37828
rect 15289 37825 15301 37828
rect 15335 37825 15347 37859
rect 15396 37856 15424 37896
rect 15562 37884 15568 37936
rect 15620 37924 15626 37936
rect 17052 37924 17080 37964
rect 19061 37961 19073 37964
rect 19107 37961 19119 37995
rect 19061 37955 19119 37961
rect 19518 37952 19524 38004
rect 19576 37952 19582 38004
rect 20622 37952 20628 38004
rect 20680 37952 20686 38004
rect 20993 37995 21051 38001
rect 20993 37961 21005 37995
rect 21039 37961 21051 37995
rect 20993 37955 21051 37961
rect 15620 37896 17080 37924
rect 18325 37927 18383 37933
rect 15620 37884 15626 37896
rect 18325 37893 18337 37927
rect 18371 37924 18383 37927
rect 18414 37924 18420 37936
rect 18371 37896 18420 37924
rect 18371 37893 18383 37896
rect 18325 37887 18383 37893
rect 18414 37884 18420 37896
rect 18472 37884 18478 37936
rect 18874 37884 18880 37936
rect 18932 37924 18938 37936
rect 20533 37927 20591 37933
rect 20533 37924 20545 37927
rect 18932 37896 20545 37924
rect 18932 37884 18938 37896
rect 20533 37893 20545 37896
rect 20579 37924 20591 37927
rect 21008 37924 21036 37955
rect 21266 37952 21272 38004
rect 21324 37952 21330 38004
rect 22186 37992 22192 38004
rect 22066 37964 22192 37992
rect 21726 37924 21732 37936
rect 20579 37896 20760 37924
rect 21008 37896 21732 37924
rect 20579 37893 20591 37896
rect 20533 37887 20591 37893
rect 15654 37856 15660 37868
rect 15396 37828 15660 37856
rect 15289 37819 15347 37825
rect 15654 37816 15660 37828
rect 15712 37816 15718 37868
rect 16114 37816 16120 37868
rect 16172 37816 16178 37868
rect 16942 37816 16948 37868
rect 17000 37856 17006 37868
rect 19429 37859 19487 37865
rect 17000 37842 17250 37856
rect 17000 37828 17264 37842
rect 17000 37816 17006 37828
rect 12406 37760 13952 37788
rect 12253 37751 12311 37757
rect 11241 37723 11299 37729
rect 11241 37720 11253 37723
rect 8680 37692 11253 37720
rect 11241 37689 11253 37692
rect 11287 37689 11299 37723
rect 11241 37683 11299 37689
rect 11422 37680 11428 37732
rect 11480 37720 11486 37732
rect 12897 37723 12955 37729
rect 12897 37720 12909 37723
rect 11480 37692 12909 37720
rect 11480 37680 11486 37692
rect 12897 37689 12909 37692
rect 12943 37689 12955 37723
rect 13924 37720 13952 37760
rect 13998 37748 14004 37800
rect 14056 37748 14062 37800
rect 14274 37748 14280 37800
rect 14332 37788 14338 37800
rect 14645 37791 14703 37797
rect 14645 37788 14657 37791
rect 14332 37760 14657 37788
rect 14332 37748 14338 37760
rect 14645 37757 14657 37760
rect 14691 37788 14703 37791
rect 15212 37788 15240 37816
rect 14691 37760 15240 37788
rect 14691 37757 14703 37760
rect 14645 37751 14703 37757
rect 15378 37748 15384 37800
rect 15436 37748 15442 37800
rect 15565 37791 15623 37797
rect 15565 37757 15577 37791
rect 15611 37788 15623 37791
rect 16132 37788 16160 37816
rect 15611 37760 16160 37788
rect 17236 37788 17264 37828
rect 19429 37825 19441 37859
rect 19475 37856 19487 37859
rect 20346 37856 20352 37868
rect 19475 37828 20352 37856
rect 19475 37825 19487 37828
rect 19429 37819 19487 37825
rect 20346 37816 20352 37828
rect 20404 37816 20410 37868
rect 20732 37856 20760 37896
rect 21726 37884 21732 37896
rect 21784 37884 21790 37936
rect 21453 37859 21511 37865
rect 21453 37856 21465 37859
rect 20732 37828 21465 37856
rect 21453 37825 21465 37828
rect 21499 37856 21511 37859
rect 22066 37856 22094 37964
rect 22186 37952 22192 37964
rect 22244 37952 22250 38004
rect 23750 37992 23756 38004
rect 22664 37964 23756 37992
rect 21499 37828 22094 37856
rect 22189 37859 22247 37865
rect 21499 37825 21511 37828
rect 21453 37819 21511 37825
rect 22189 37825 22201 37859
rect 22235 37856 22247 37859
rect 22370 37856 22376 37868
rect 22235 37828 22376 37856
rect 22235 37825 22247 37828
rect 22189 37819 22247 37825
rect 22370 37816 22376 37828
rect 22428 37816 22434 37868
rect 17770 37788 17776 37800
rect 17236 37760 17776 37788
rect 15611 37757 15623 37760
rect 15565 37751 15623 37757
rect 17770 37748 17776 37760
rect 17828 37748 17834 37800
rect 18601 37791 18659 37797
rect 18601 37757 18613 37791
rect 18647 37788 18659 37791
rect 19613 37791 19671 37797
rect 18647 37760 19334 37788
rect 18647 37757 18659 37760
rect 18601 37751 18659 37757
rect 16114 37720 16120 37732
rect 13924 37692 16120 37720
rect 12897 37683 12955 37689
rect 16114 37680 16120 37692
rect 16172 37680 16178 37732
rect 19306 37720 19334 37760
rect 19613 37757 19625 37791
rect 19659 37757 19671 37791
rect 19613 37751 19671 37757
rect 20441 37791 20499 37797
rect 20441 37757 20453 37791
rect 20487 37788 20499 37791
rect 21542 37788 21548 37800
rect 20487 37760 21548 37788
rect 20487 37757 20499 37760
rect 20441 37751 20499 37757
rect 19426 37720 19432 37732
rect 19306 37692 19432 37720
rect 19426 37680 19432 37692
rect 19484 37680 19490 37732
rect 8938 37612 8944 37664
rect 8996 37652 9002 37664
rect 9493 37655 9551 37661
rect 9493 37652 9505 37655
rect 8996 37624 9505 37652
rect 8996 37612 9002 37624
rect 9493 37621 9505 37624
rect 9539 37621 9551 37655
rect 9493 37615 9551 37621
rect 11606 37612 11612 37664
rect 11664 37652 11670 37664
rect 11701 37655 11759 37661
rect 11701 37652 11713 37655
rect 11664 37624 11713 37652
rect 11664 37612 11670 37624
rect 11701 37621 11713 37624
rect 11747 37621 11759 37655
rect 11701 37615 11759 37621
rect 13722 37612 13728 37664
rect 13780 37652 13786 37664
rect 14921 37655 14979 37661
rect 14921 37652 14933 37655
rect 13780 37624 14933 37652
rect 13780 37612 13786 37624
rect 14921 37621 14933 37624
rect 14967 37621 14979 37655
rect 14921 37615 14979 37621
rect 17310 37612 17316 37664
rect 17368 37652 17374 37664
rect 19628 37652 19656 37751
rect 21542 37748 21548 37760
rect 21600 37748 21606 37800
rect 22278 37748 22284 37800
rect 22336 37788 22342 37800
rect 22664 37797 22692 37964
rect 23750 37952 23756 37964
rect 23808 37952 23814 38004
rect 24394 37952 24400 38004
rect 24452 37952 24458 38004
rect 23658 37884 23664 37936
rect 23716 37884 23722 37936
rect 24210 37816 24216 37868
rect 24268 37856 24274 37868
rect 24762 37856 24768 37868
rect 24268 37828 24768 37856
rect 24268 37816 24274 37828
rect 24762 37816 24768 37828
rect 24820 37856 24826 37868
rect 25317 37859 25375 37865
rect 25317 37856 25329 37859
rect 24820 37828 25329 37856
rect 24820 37816 24826 37828
rect 25317 37825 25329 37828
rect 25363 37825 25375 37859
rect 25317 37819 25375 37825
rect 22649 37791 22707 37797
rect 22649 37788 22661 37791
rect 22336 37760 22661 37788
rect 22336 37748 22342 37760
rect 22649 37757 22661 37760
rect 22695 37757 22707 37791
rect 22925 37791 22983 37797
rect 22925 37788 22937 37791
rect 22649 37751 22707 37757
rect 22756 37760 22937 37788
rect 22462 37680 22468 37732
rect 22520 37720 22526 37732
rect 22756 37720 22784 37760
rect 22925 37757 22937 37760
rect 22971 37757 22983 37791
rect 22925 37751 22983 37757
rect 23658 37748 23664 37800
rect 23716 37788 23722 37800
rect 24673 37791 24731 37797
rect 24673 37788 24685 37791
rect 23716 37760 24685 37788
rect 23716 37748 23722 37760
rect 24673 37757 24685 37760
rect 24719 37757 24731 37791
rect 24673 37751 24731 37757
rect 22520 37692 22784 37720
rect 22520 37680 22526 37692
rect 17368 37624 19656 37652
rect 17368 37612 17374 37624
rect 21542 37612 21548 37664
rect 21600 37652 21606 37664
rect 22005 37655 22063 37661
rect 22005 37652 22017 37655
rect 21600 37624 22017 37652
rect 21600 37612 21606 37624
rect 22005 37621 22017 37624
rect 22051 37621 22063 37655
rect 22005 37615 22063 37621
rect 25133 37655 25191 37661
rect 25133 37621 25145 37655
rect 25179 37652 25191 37655
rect 25498 37652 25504 37664
rect 25179 37624 25504 37652
rect 25179 37621 25191 37624
rect 25133 37615 25191 37621
rect 25498 37612 25504 37624
rect 25556 37612 25562 37664
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 7650 37408 7656 37460
rect 7708 37448 7714 37460
rect 8205 37451 8263 37457
rect 8205 37448 8217 37451
rect 7708 37420 8217 37448
rect 7708 37408 7714 37420
rect 8205 37417 8217 37420
rect 8251 37417 8263 37451
rect 8205 37411 8263 37417
rect 11054 37408 11060 37460
rect 11112 37448 11118 37460
rect 11974 37448 11980 37460
rect 11112 37420 11980 37448
rect 11112 37408 11118 37420
rect 11974 37408 11980 37420
rect 12032 37408 12038 37460
rect 14458 37408 14464 37460
rect 14516 37408 14522 37460
rect 16114 37408 16120 37460
rect 16172 37408 16178 37460
rect 18874 37408 18880 37460
rect 18932 37448 18938 37460
rect 19058 37448 19064 37460
rect 18932 37420 19064 37448
rect 18932 37408 18938 37420
rect 19058 37408 19064 37420
rect 19116 37448 19122 37460
rect 20809 37451 20867 37457
rect 20809 37448 20821 37451
rect 19116 37420 20821 37448
rect 19116 37408 19122 37420
rect 20809 37417 20821 37420
rect 20855 37417 20867 37451
rect 20809 37411 20867 37417
rect 21085 37451 21143 37457
rect 21085 37417 21097 37451
rect 21131 37448 21143 37451
rect 21266 37448 21272 37460
rect 21131 37420 21272 37448
rect 21131 37417 21143 37420
rect 21085 37411 21143 37417
rect 21266 37408 21272 37420
rect 21324 37408 21330 37460
rect 23658 37408 23664 37460
rect 23716 37448 23722 37460
rect 23937 37451 23995 37457
rect 23937 37448 23949 37451
rect 23716 37420 23949 37448
rect 23716 37408 23722 37420
rect 23937 37417 23949 37420
rect 23983 37417 23995 37451
rect 23937 37411 23995 37417
rect 24118 37408 24124 37460
rect 24176 37408 24182 37460
rect 24210 37408 24216 37460
rect 24268 37408 24274 37460
rect 6546 37340 6552 37392
rect 6604 37380 6610 37392
rect 8570 37380 8576 37392
rect 6604 37352 8576 37380
rect 6604 37340 6610 37352
rect 8570 37340 8576 37352
rect 8628 37380 8634 37392
rect 14366 37380 14372 37392
rect 8628 37352 9260 37380
rect 8628 37340 8634 37352
rect 9232 37324 9260 37352
rect 13188 37352 14372 37380
rect 5994 37272 6000 37324
rect 6052 37312 6058 37324
rect 7561 37315 7619 37321
rect 7561 37312 7573 37315
rect 6052 37284 7573 37312
rect 6052 37272 6058 37284
rect 7561 37281 7573 37284
rect 7607 37281 7619 37315
rect 7561 37275 7619 37281
rect 9214 37272 9220 37324
rect 9272 37272 9278 37324
rect 9306 37272 9312 37324
rect 9364 37312 9370 37324
rect 11057 37315 11115 37321
rect 11057 37312 11069 37315
rect 9364 37284 11069 37312
rect 9364 37272 9370 37284
rect 11057 37281 11069 37284
rect 11103 37281 11115 37315
rect 11330 37312 11336 37324
rect 11057 37275 11115 37281
rect 11164 37284 11336 37312
rect 7745 37247 7803 37253
rect 7745 37213 7757 37247
rect 7791 37244 7803 37247
rect 8938 37244 8944 37256
rect 7791 37216 8944 37244
rect 7791 37213 7803 37216
rect 7745 37207 7803 37213
rect 8938 37204 8944 37216
rect 8996 37204 9002 37256
rect 10045 37247 10103 37253
rect 10045 37213 10057 37247
rect 10091 37244 10103 37247
rect 10594 37244 10600 37256
rect 10091 37216 10600 37244
rect 10091 37213 10103 37216
rect 10045 37207 10103 37213
rect 10594 37204 10600 37216
rect 10652 37204 10658 37256
rect 11164 37244 11192 37284
rect 11330 37272 11336 37284
rect 11388 37312 11394 37324
rect 13188 37321 13216 37352
rect 14366 37340 14372 37352
rect 14424 37340 14430 37392
rect 13173 37315 13231 37321
rect 11388 37284 13032 37312
rect 11388 37272 11394 37284
rect 10704 37216 11192 37244
rect 12529 37247 12587 37253
rect 8662 37136 8668 37188
rect 8720 37176 8726 37188
rect 10704 37176 10732 37216
rect 12529 37213 12541 37247
rect 12575 37244 12587 37247
rect 12618 37244 12624 37256
rect 12575 37216 12624 37244
rect 12575 37213 12587 37216
rect 12529 37207 12587 37213
rect 12618 37204 12624 37216
rect 12676 37204 12682 37256
rect 13004 37244 13032 37284
rect 13173 37281 13185 37315
rect 13219 37281 13231 37315
rect 14093 37315 14151 37321
rect 14093 37312 14105 37315
rect 13173 37275 13231 37281
rect 13280 37284 14105 37312
rect 13280 37253 13308 37284
rect 14093 37281 14105 37284
rect 14139 37281 14151 37315
rect 14476 37312 14504 37408
rect 15841 37383 15899 37389
rect 15841 37380 15853 37383
rect 15396 37352 15853 37380
rect 14476 37284 14780 37312
rect 14093 37275 14151 37281
rect 13265 37247 13323 37253
rect 13265 37244 13277 37247
rect 13004 37216 13277 37244
rect 13265 37213 13277 37216
rect 13311 37213 13323 37247
rect 13265 37207 13323 37213
rect 13357 37247 13415 37253
rect 13357 37213 13369 37247
rect 13403 37244 13415 37247
rect 13998 37244 14004 37256
rect 13403 37216 14004 37244
rect 13403 37213 13415 37216
rect 13357 37207 13415 37213
rect 13998 37204 14004 37216
rect 14056 37204 14062 37256
rect 8720 37148 10732 37176
rect 10965 37179 11023 37185
rect 8720 37136 8726 37148
rect 10965 37145 10977 37179
rect 11011 37176 11023 37179
rect 13630 37176 13636 37188
rect 11011 37148 13636 37176
rect 11011 37145 11023 37148
rect 10965 37139 11023 37145
rect 13630 37136 13636 37148
rect 13688 37136 13694 37188
rect 14752 37176 14780 37284
rect 14826 37272 14832 37324
rect 14884 37312 14890 37324
rect 15289 37315 15347 37321
rect 15289 37312 15301 37315
rect 14884 37284 15301 37312
rect 14884 37272 14890 37284
rect 15289 37281 15301 37284
rect 15335 37281 15347 37315
rect 15289 37275 15347 37281
rect 15105 37247 15163 37253
rect 15105 37213 15117 37247
rect 15151 37244 15163 37247
rect 15396 37244 15424 37352
rect 15841 37349 15853 37352
rect 15887 37380 15899 37383
rect 23290 37380 23296 37392
rect 15887 37352 23296 37380
rect 15887 37349 15899 37352
rect 15841 37343 15899 37349
rect 23290 37340 23296 37352
rect 23348 37340 23354 37392
rect 15930 37272 15936 37324
rect 15988 37312 15994 37324
rect 16669 37315 16727 37321
rect 16669 37312 16681 37315
rect 15988 37284 16681 37312
rect 15988 37272 15994 37284
rect 16669 37281 16681 37284
rect 16715 37281 16727 37315
rect 16669 37275 16727 37281
rect 17218 37272 17224 37324
rect 17276 37312 17282 37324
rect 17862 37312 17868 37324
rect 17276 37284 17868 37312
rect 17276 37272 17282 37284
rect 17862 37272 17868 37284
rect 17920 37272 17926 37324
rect 18601 37315 18659 37321
rect 18601 37312 18613 37315
rect 17972 37284 18613 37312
rect 15151 37216 15424 37244
rect 15151 37213 15163 37216
rect 15105 37207 15163 37213
rect 17310 37204 17316 37256
rect 17368 37244 17374 37256
rect 17972 37244 18000 37284
rect 18601 37281 18613 37284
rect 18647 37281 18659 37315
rect 20717 37315 20775 37321
rect 20717 37312 20729 37315
rect 18601 37275 18659 37281
rect 18800 37284 20729 37312
rect 18800 37256 18828 37284
rect 20717 37281 20729 37284
rect 20763 37281 20775 37315
rect 24136 37312 24164 37408
rect 20717 37275 20775 37281
rect 24044 37284 24164 37312
rect 24044 37256 24072 37284
rect 17368 37216 18000 37244
rect 18417 37247 18475 37253
rect 17368 37204 17374 37216
rect 18417 37213 18429 37247
rect 18463 37244 18475 37247
rect 18782 37244 18788 37256
rect 18463 37216 18788 37244
rect 18463 37213 18475 37216
rect 18417 37207 18475 37213
rect 18782 37204 18788 37216
rect 18840 37204 18846 37256
rect 20349 37247 20407 37253
rect 20349 37213 20361 37247
rect 20395 37244 20407 37247
rect 21266 37244 21272 37256
rect 20395 37216 21272 37244
rect 20395 37213 20407 37216
rect 20349 37207 20407 37213
rect 21266 37204 21272 37216
rect 21324 37244 21330 37256
rect 21453 37247 21511 37253
rect 21453 37244 21465 37247
rect 21324 37216 21465 37244
rect 21324 37204 21330 37216
rect 21453 37213 21465 37216
rect 21499 37213 21511 37247
rect 21453 37207 21511 37213
rect 22094 37204 22100 37256
rect 22152 37244 22158 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22152 37216 22845 37244
rect 22152 37204 22158 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 22833 37207 22891 37213
rect 24026 37204 24032 37256
rect 24084 37204 24090 37256
rect 24118 37204 24124 37256
rect 24176 37244 24182 37256
rect 24394 37244 24400 37256
rect 24176 37216 24400 37244
rect 24176 37204 24182 37216
rect 24394 37204 24400 37216
rect 24452 37244 24458 37256
rect 24581 37247 24639 37253
rect 24581 37244 24593 37247
rect 24452 37216 24593 37244
rect 24452 37204 24458 37216
rect 24581 37213 24593 37216
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 15197 37179 15255 37185
rect 15197 37176 15209 37179
rect 14752 37148 15209 37176
rect 15197 37145 15209 37148
rect 15243 37145 15255 37179
rect 15197 37139 15255 37145
rect 16485 37179 16543 37185
rect 16485 37145 16497 37179
rect 16531 37176 16543 37179
rect 18598 37176 18604 37188
rect 16531 37148 18604 37176
rect 16531 37145 16543 37148
rect 16485 37139 16543 37145
rect 18598 37136 18604 37148
rect 18656 37136 18662 37188
rect 19334 37136 19340 37188
rect 19392 37176 19398 37188
rect 19521 37179 19579 37185
rect 19521 37176 19533 37179
rect 19392 37148 19533 37176
rect 19392 37136 19398 37148
rect 19521 37145 19533 37148
rect 19567 37145 19579 37179
rect 19521 37139 19579 37145
rect 22278 37136 22284 37188
rect 22336 37136 22342 37188
rect 25958 37176 25964 37188
rect 22388 37148 25964 37176
rect 7837 37111 7895 37117
rect 7837 37077 7849 37111
rect 7883 37108 7895 37111
rect 9122 37108 9128 37120
rect 7883 37080 9128 37108
rect 7883 37077 7895 37080
rect 7837 37071 7895 37077
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 10226 37068 10232 37120
rect 10284 37108 10290 37120
rect 10505 37111 10563 37117
rect 10505 37108 10517 37111
rect 10284 37080 10517 37108
rect 10284 37068 10290 37080
rect 10505 37077 10517 37080
rect 10551 37077 10563 37111
rect 10505 37071 10563 37077
rect 10870 37068 10876 37120
rect 10928 37068 10934 37120
rect 11885 37111 11943 37117
rect 11885 37077 11897 37111
rect 11931 37108 11943 37111
rect 11974 37108 11980 37120
rect 11931 37080 11980 37108
rect 11931 37077 11943 37080
rect 11885 37071 11943 37077
rect 11974 37068 11980 37080
rect 12032 37068 12038 37120
rect 13725 37111 13783 37117
rect 13725 37077 13737 37111
rect 13771 37108 13783 37111
rect 13814 37108 13820 37120
rect 13771 37080 13820 37108
rect 13771 37077 13783 37080
rect 13725 37071 13783 37077
rect 13814 37068 13820 37080
rect 13872 37068 13878 37120
rect 14734 37068 14740 37120
rect 14792 37068 14798 37120
rect 15286 37068 15292 37120
rect 15344 37108 15350 37120
rect 15930 37108 15936 37120
rect 15344 37080 15936 37108
rect 15344 37068 15350 37080
rect 15930 37068 15936 37080
rect 15988 37068 15994 37120
rect 16574 37068 16580 37120
rect 16632 37068 16638 37120
rect 17218 37068 17224 37120
rect 17276 37108 17282 37120
rect 17313 37111 17371 37117
rect 17313 37108 17325 37111
rect 17276 37080 17325 37108
rect 17276 37068 17282 37080
rect 17313 37077 17325 37080
rect 17359 37077 17371 37111
rect 17313 37071 17371 37077
rect 17402 37068 17408 37120
rect 17460 37108 17466 37120
rect 18049 37111 18107 37117
rect 18049 37108 18061 37111
rect 17460 37080 18061 37108
rect 17460 37068 17466 37080
rect 18049 37077 18061 37080
rect 18095 37077 18107 37111
rect 18049 37071 18107 37077
rect 18509 37111 18567 37117
rect 18509 37077 18521 37111
rect 18555 37108 18567 37111
rect 18874 37108 18880 37120
rect 18555 37080 18880 37108
rect 18555 37077 18567 37080
rect 18509 37071 18567 37077
rect 18874 37068 18880 37080
rect 18932 37068 18938 37120
rect 19610 37068 19616 37120
rect 19668 37108 19674 37120
rect 20622 37108 20628 37120
rect 19668 37080 20628 37108
rect 19668 37068 19674 37080
rect 20622 37068 20628 37080
rect 20680 37108 20686 37120
rect 22388 37108 22416 37148
rect 25958 37136 25964 37148
rect 26016 37136 26022 37188
rect 20680 37080 22416 37108
rect 20680 37068 20686 37080
rect 22646 37068 22652 37120
rect 22704 37108 22710 37120
rect 23477 37111 23535 37117
rect 23477 37108 23489 37111
rect 22704 37080 23489 37108
rect 22704 37068 22710 37080
rect 23477 37077 23489 37080
rect 23523 37077 23535 37111
rect 23477 37071 23535 37077
rect 25038 37068 25044 37120
rect 25096 37108 25102 37120
rect 25225 37111 25283 37117
rect 25225 37108 25237 37111
rect 25096 37080 25237 37108
rect 25096 37068 25102 37080
rect 25225 37077 25237 37080
rect 25271 37077 25283 37111
rect 25225 37071 25283 37077
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 7466 36864 7472 36916
rect 7524 36904 7530 36916
rect 10042 36904 10048 36916
rect 7524 36876 10048 36904
rect 7524 36864 7530 36876
rect 10042 36864 10048 36876
rect 10100 36864 10106 36916
rect 10594 36864 10600 36916
rect 10652 36904 10658 36916
rect 11517 36907 11575 36913
rect 11517 36904 11529 36907
rect 10652 36876 11529 36904
rect 10652 36864 10658 36876
rect 6362 36796 6368 36848
rect 6420 36836 6426 36848
rect 7650 36836 7656 36848
rect 6420 36808 7656 36836
rect 6420 36796 6426 36808
rect 7650 36796 7656 36808
rect 7708 36836 7714 36848
rect 8941 36839 8999 36845
rect 7708 36808 7774 36836
rect 7708 36796 7714 36808
rect 8941 36805 8953 36839
rect 8987 36836 8999 36839
rect 9030 36836 9036 36848
rect 8987 36808 9036 36836
rect 8987 36805 8999 36808
rect 8941 36799 8999 36805
rect 9030 36796 9036 36808
rect 9088 36836 9094 36848
rect 11164 36845 11192 36876
rect 11517 36873 11529 36876
rect 11563 36904 11575 36907
rect 15286 36904 15292 36916
rect 11563 36876 15292 36904
rect 11563 36873 11575 36876
rect 11517 36867 11575 36873
rect 15286 36864 15292 36876
rect 15344 36864 15350 36916
rect 15930 36864 15936 36916
rect 15988 36864 15994 36916
rect 16390 36864 16396 36916
rect 16448 36904 16454 36916
rect 17129 36907 17187 36913
rect 17129 36904 17141 36907
rect 16448 36876 17141 36904
rect 16448 36864 16454 36876
rect 17129 36873 17141 36876
rect 17175 36873 17187 36907
rect 17129 36867 17187 36873
rect 17218 36864 17224 36916
rect 17276 36864 17282 36916
rect 17589 36907 17647 36913
rect 17589 36873 17601 36907
rect 17635 36904 17647 36907
rect 19702 36904 19708 36916
rect 17635 36876 19708 36904
rect 17635 36873 17647 36876
rect 17589 36867 17647 36873
rect 19702 36864 19708 36876
rect 19760 36864 19766 36916
rect 20162 36864 20168 36916
rect 20220 36904 20226 36916
rect 20625 36907 20683 36913
rect 20625 36904 20637 36907
rect 20220 36876 20637 36904
rect 20220 36864 20226 36876
rect 20625 36873 20637 36876
rect 20671 36873 20683 36907
rect 20625 36867 20683 36873
rect 21358 36864 21364 36916
rect 21416 36904 21422 36916
rect 21453 36907 21511 36913
rect 21453 36904 21465 36907
rect 21416 36876 21465 36904
rect 21416 36864 21422 36876
rect 21453 36873 21465 36876
rect 21499 36873 21511 36907
rect 21453 36867 21511 36873
rect 21634 36864 21640 36916
rect 21692 36904 21698 36916
rect 22186 36904 22192 36916
rect 21692 36876 22192 36904
rect 21692 36864 21698 36876
rect 22186 36864 22192 36876
rect 22244 36904 22250 36916
rect 22281 36907 22339 36913
rect 22281 36904 22293 36907
rect 22244 36876 22293 36904
rect 22244 36864 22250 36876
rect 22281 36873 22293 36876
rect 22327 36904 22339 36907
rect 22741 36907 22799 36913
rect 22327 36876 22600 36904
rect 22327 36873 22339 36876
rect 22281 36867 22339 36873
rect 9493 36839 9551 36845
rect 9493 36836 9505 36839
rect 9088 36808 9505 36836
rect 9088 36796 9094 36808
rect 9493 36805 9505 36808
rect 9539 36805 9551 36839
rect 9493 36799 9551 36805
rect 11149 36839 11207 36845
rect 11149 36805 11161 36839
rect 11195 36836 11207 36839
rect 11195 36808 11229 36836
rect 11195 36805 11207 36808
rect 11149 36799 11207 36805
rect 12618 36796 12624 36848
rect 12676 36836 12682 36848
rect 13722 36836 13728 36848
rect 12676 36808 13728 36836
rect 12676 36796 12682 36808
rect 13722 36796 13728 36808
rect 13780 36796 13786 36848
rect 15102 36796 15108 36848
rect 15160 36796 15166 36848
rect 19610 36836 19616 36848
rect 18892 36808 19616 36836
rect 9214 36728 9220 36780
rect 9272 36728 9278 36780
rect 9398 36728 9404 36780
rect 9456 36768 9462 36780
rect 12989 36771 13047 36777
rect 9456 36740 12020 36768
rect 9456 36728 9462 36740
rect 10318 36660 10324 36712
rect 10376 36660 10382 36712
rect 11992 36709 12020 36740
rect 12989 36737 13001 36771
rect 13035 36768 13047 36771
rect 13633 36771 13691 36777
rect 13633 36768 13645 36771
rect 13035 36740 13645 36768
rect 13035 36737 13047 36740
rect 12989 36731 13047 36737
rect 13633 36737 13645 36740
rect 13679 36737 13691 36771
rect 13633 36731 13691 36737
rect 15013 36771 15071 36777
rect 15013 36737 15025 36771
rect 15059 36768 15071 36771
rect 15930 36768 15936 36780
rect 15059 36740 15936 36768
rect 15059 36737 15071 36740
rect 15013 36731 15071 36737
rect 11977 36703 12035 36709
rect 11977 36669 11989 36703
rect 12023 36700 12035 36703
rect 13081 36703 13139 36709
rect 13081 36700 13093 36703
rect 12023 36672 13093 36700
rect 12023 36669 12035 36672
rect 11977 36663 12035 36669
rect 13081 36669 13093 36672
rect 13127 36669 13139 36703
rect 13081 36663 13139 36669
rect 13173 36703 13231 36709
rect 13173 36669 13185 36703
rect 13219 36669 13231 36703
rect 13173 36663 13231 36669
rect 12710 36592 12716 36644
rect 12768 36632 12774 36644
rect 13188 36632 13216 36663
rect 12768 36604 13216 36632
rect 13648 36632 13676 36731
rect 15930 36728 15936 36740
rect 15988 36728 15994 36780
rect 13722 36660 13728 36712
rect 13780 36700 13786 36712
rect 15197 36703 15255 36709
rect 15197 36700 15209 36703
rect 13780 36672 15209 36700
rect 13780 36660 13786 36672
rect 15197 36669 15209 36672
rect 15243 36669 15255 36703
rect 15197 36663 15255 36669
rect 17037 36703 17095 36709
rect 17037 36669 17049 36703
rect 17083 36700 17095 36703
rect 17494 36700 17500 36712
rect 17083 36672 17500 36700
rect 17083 36669 17095 36672
rect 17037 36663 17095 36669
rect 17494 36660 17500 36672
rect 17552 36660 17558 36712
rect 18892 36632 18920 36808
rect 19610 36796 19616 36808
rect 19668 36796 19674 36848
rect 20530 36796 20536 36848
rect 20588 36836 20594 36848
rect 20717 36839 20775 36845
rect 20717 36836 20729 36839
rect 20588 36808 20729 36836
rect 20588 36796 20594 36808
rect 20717 36805 20729 36808
rect 20763 36836 20775 36839
rect 21269 36839 21327 36845
rect 21269 36836 21281 36839
rect 20763 36808 21281 36836
rect 20763 36805 20775 36808
rect 20717 36799 20775 36805
rect 21269 36805 21281 36808
rect 21315 36805 21327 36839
rect 22462 36836 22468 36848
rect 21269 36799 21327 36805
rect 22112 36808 22468 36836
rect 19337 36771 19395 36777
rect 19337 36737 19349 36771
rect 19383 36768 19395 36771
rect 19978 36768 19984 36780
rect 19383 36740 19984 36768
rect 19383 36737 19395 36740
rect 19337 36731 19395 36737
rect 19978 36728 19984 36740
rect 20036 36728 20042 36780
rect 19429 36703 19487 36709
rect 19429 36669 19441 36703
rect 19475 36669 19487 36703
rect 19429 36663 19487 36669
rect 13648 36604 18920 36632
rect 12768 36592 12774 36604
rect 18966 36592 18972 36644
rect 19024 36592 19030 36644
rect 19444 36632 19472 36663
rect 19518 36660 19524 36712
rect 19576 36660 19582 36712
rect 20438 36660 20444 36712
rect 20496 36700 20502 36712
rect 22112 36709 22140 36808
rect 22462 36796 22468 36808
rect 22520 36796 22526 36848
rect 22572 36836 22600 36876
rect 22741 36873 22753 36907
rect 22787 36904 22799 36907
rect 23382 36904 23388 36916
rect 22787 36876 23388 36904
rect 22787 36873 22799 36876
rect 22741 36867 22799 36873
rect 23382 36864 23388 36876
rect 23440 36864 23446 36916
rect 23569 36907 23627 36913
rect 23569 36873 23581 36907
rect 23615 36904 23627 36907
rect 24670 36904 24676 36916
rect 23615 36876 24676 36904
rect 23615 36873 23627 36876
rect 23569 36867 23627 36873
rect 24670 36864 24676 36876
rect 24728 36864 24734 36916
rect 23017 36839 23075 36845
rect 23017 36836 23029 36839
rect 22572 36808 23029 36836
rect 23017 36805 23029 36808
rect 23063 36805 23075 36839
rect 23017 36799 23075 36805
rect 23658 36796 23664 36848
rect 23716 36836 23722 36848
rect 23716 36822 23874 36836
rect 23716 36808 23888 36822
rect 23716 36796 23722 36808
rect 22373 36771 22431 36777
rect 22373 36737 22385 36771
rect 22419 36768 22431 36771
rect 22419 36740 23244 36768
rect 22419 36737 22431 36740
rect 22373 36731 22431 36737
rect 20809 36703 20867 36709
rect 20809 36700 20821 36703
rect 20496 36672 20821 36700
rect 20496 36660 20502 36672
rect 20809 36669 20821 36672
rect 20855 36669 20867 36703
rect 20809 36663 20867 36669
rect 22097 36703 22155 36709
rect 22097 36669 22109 36703
rect 22143 36669 22155 36703
rect 22097 36663 22155 36669
rect 20990 36632 20996 36644
rect 19444 36604 20996 36632
rect 20990 36592 20996 36604
rect 21048 36592 21054 36644
rect 21358 36592 21364 36644
rect 21416 36632 21422 36644
rect 22186 36632 22192 36644
rect 21416 36604 22192 36632
rect 21416 36592 21422 36604
rect 22186 36592 22192 36604
rect 22244 36592 22250 36644
rect 6822 36524 6828 36576
rect 6880 36564 6886 36576
rect 12158 36564 12164 36576
rect 6880 36536 12164 36564
rect 6880 36524 6886 36536
rect 12158 36524 12164 36536
rect 12216 36524 12222 36576
rect 12250 36524 12256 36576
rect 12308 36524 12314 36576
rect 12342 36524 12348 36576
rect 12400 36564 12406 36576
rect 12621 36567 12679 36573
rect 12621 36564 12633 36567
rect 12400 36536 12633 36564
rect 12400 36524 12406 36536
rect 12621 36533 12633 36536
rect 12667 36533 12679 36567
rect 12621 36527 12679 36533
rect 14366 36524 14372 36576
rect 14424 36564 14430 36576
rect 14645 36567 14703 36573
rect 14645 36564 14657 36567
rect 14424 36536 14657 36564
rect 14424 36524 14430 36536
rect 14645 36533 14657 36536
rect 14691 36533 14703 36567
rect 14645 36527 14703 36533
rect 15749 36567 15807 36573
rect 15749 36533 15761 36567
rect 15795 36564 15807 36567
rect 15930 36564 15936 36576
rect 15795 36536 15936 36564
rect 15795 36533 15807 36536
rect 15749 36527 15807 36533
rect 15930 36524 15936 36536
rect 15988 36524 15994 36576
rect 19518 36524 19524 36576
rect 19576 36564 19582 36576
rect 23216 36573 23244 36740
rect 23860 36700 23888 36808
rect 25038 36796 25044 36848
rect 25096 36796 25102 36848
rect 25038 36700 25044 36712
rect 23860 36672 25044 36700
rect 25038 36660 25044 36672
rect 25096 36660 25102 36712
rect 25317 36703 25375 36709
rect 25317 36700 25329 36703
rect 25240 36672 25329 36700
rect 20257 36567 20315 36573
rect 20257 36564 20269 36567
rect 19576 36536 20269 36564
rect 19576 36524 19582 36536
rect 20257 36533 20269 36536
rect 20303 36533 20315 36567
rect 20257 36527 20315 36533
rect 23201 36567 23259 36573
rect 23201 36533 23213 36567
rect 23247 36564 23259 36567
rect 23382 36564 23388 36576
rect 23247 36536 23388 36564
rect 23247 36533 23259 36536
rect 23201 36527 23259 36533
rect 23382 36524 23388 36536
rect 23440 36564 23446 36576
rect 24854 36564 24860 36576
rect 23440 36536 24860 36564
rect 23440 36524 23446 36536
rect 24854 36524 24860 36536
rect 24912 36524 24918 36576
rect 24946 36524 24952 36576
rect 25004 36564 25010 36576
rect 25240 36564 25268 36672
rect 25317 36669 25329 36672
rect 25363 36669 25375 36703
rect 25317 36663 25375 36669
rect 25004 36536 25268 36564
rect 25004 36524 25010 36536
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 7006 36320 7012 36372
rect 7064 36360 7070 36372
rect 9493 36363 9551 36369
rect 9493 36360 9505 36363
rect 7064 36332 9505 36360
rect 7064 36320 7070 36332
rect 9493 36329 9505 36332
rect 9539 36329 9551 36363
rect 9493 36323 9551 36329
rect 13173 36363 13231 36369
rect 13173 36329 13185 36363
rect 13219 36360 13231 36363
rect 13354 36360 13360 36372
rect 13219 36332 13360 36360
rect 13219 36329 13231 36332
rect 13173 36323 13231 36329
rect 13354 36320 13360 36332
rect 13412 36320 13418 36372
rect 15013 36363 15071 36369
rect 15013 36329 15025 36363
rect 15059 36360 15071 36363
rect 15470 36360 15476 36372
rect 15059 36332 15476 36360
rect 15059 36329 15071 36332
rect 15013 36323 15071 36329
rect 15470 36320 15476 36332
rect 15528 36320 15534 36372
rect 16574 36320 16580 36372
rect 16632 36360 16638 36372
rect 16945 36363 17003 36369
rect 16945 36360 16957 36363
rect 16632 36332 16957 36360
rect 16632 36320 16638 36332
rect 16945 36329 16957 36332
rect 16991 36360 17003 36363
rect 17770 36360 17776 36372
rect 16991 36332 17776 36360
rect 16991 36329 17003 36332
rect 16945 36323 17003 36329
rect 17770 36320 17776 36332
rect 17828 36320 17834 36372
rect 25038 36360 25044 36372
rect 22066 36332 25044 36360
rect 17310 36252 17316 36304
rect 17368 36292 17374 36304
rect 17368 36264 20024 36292
rect 17368 36252 17374 36264
rect 5534 36184 5540 36236
rect 5592 36224 5598 36236
rect 8389 36227 8447 36233
rect 8389 36224 8401 36227
rect 5592 36196 8401 36224
rect 5592 36184 5598 36196
rect 8389 36193 8401 36196
rect 8435 36224 8447 36227
rect 10045 36227 10103 36233
rect 10045 36224 10057 36227
rect 8435 36196 10057 36224
rect 8435 36193 8447 36196
rect 8389 36187 8447 36193
rect 10045 36193 10057 36196
rect 10091 36193 10103 36227
rect 10045 36187 10103 36193
rect 12526 36184 12532 36236
rect 12584 36184 12590 36236
rect 14461 36227 14519 36233
rect 14461 36193 14473 36227
rect 14507 36224 14519 36227
rect 14918 36224 14924 36236
rect 14507 36196 14924 36224
rect 14507 36193 14519 36196
rect 14461 36187 14519 36193
rect 14918 36184 14924 36196
rect 14976 36184 14982 36236
rect 19794 36184 19800 36236
rect 19852 36224 19858 36236
rect 19996 36233 20024 36264
rect 21174 36252 21180 36304
rect 21232 36292 21238 36304
rect 21232 36264 21404 36292
rect 21232 36252 21238 36264
rect 19889 36227 19947 36233
rect 19889 36224 19901 36227
rect 19852 36196 19901 36224
rect 19852 36184 19858 36196
rect 19889 36193 19901 36196
rect 19935 36193 19947 36227
rect 19889 36187 19947 36193
rect 19981 36227 20039 36233
rect 19981 36193 19993 36227
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 20898 36184 20904 36236
rect 20956 36224 20962 36236
rect 21376 36233 21404 36264
rect 21269 36227 21327 36233
rect 21269 36224 21281 36227
rect 20956 36196 21281 36224
rect 20956 36184 20962 36196
rect 21269 36193 21281 36196
rect 21315 36193 21327 36227
rect 21269 36187 21327 36193
rect 21361 36227 21419 36233
rect 21361 36193 21373 36227
rect 21407 36193 21419 36227
rect 21361 36187 21419 36193
rect 1578 36116 1584 36168
rect 1636 36156 1642 36168
rect 2041 36159 2099 36165
rect 2041 36156 2053 36159
rect 1636 36128 2053 36156
rect 1636 36116 1642 36128
rect 2041 36125 2053 36128
rect 2087 36125 2099 36159
rect 2041 36119 2099 36125
rect 6546 36116 6552 36168
rect 6604 36156 6610 36168
rect 6641 36159 6699 36165
rect 6641 36156 6653 36159
rect 6604 36128 6653 36156
rect 6604 36116 6610 36128
rect 6641 36125 6653 36128
rect 6687 36125 6699 36159
rect 6641 36119 6699 36125
rect 9953 36159 10011 36165
rect 9953 36125 9965 36159
rect 9999 36156 10011 36159
rect 11054 36156 11060 36168
rect 9999 36128 11060 36156
rect 9999 36125 10011 36128
rect 9953 36119 10011 36125
rect 11054 36116 11060 36128
rect 11112 36116 11118 36168
rect 11698 36116 11704 36168
rect 11756 36156 11762 36168
rect 11977 36159 12035 36165
rect 11977 36156 11989 36159
rect 11756 36128 11989 36156
rect 11756 36116 11762 36128
rect 11977 36125 11989 36128
rect 12023 36156 12035 36159
rect 12066 36156 12072 36168
rect 12023 36128 12072 36156
rect 12023 36125 12035 36128
rect 11977 36119 12035 36125
rect 12066 36116 12072 36128
rect 12124 36116 12130 36168
rect 12158 36116 12164 36168
rect 12216 36156 12222 36168
rect 12805 36159 12863 36165
rect 12805 36156 12817 36159
rect 12216 36128 12817 36156
rect 12216 36116 12222 36128
rect 12805 36125 12817 36128
rect 12851 36125 12863 36159
rect 12805 36119 12863 36125
rect 15378 36116 15384 36168
rect 15436 36156 15442 36168
rect 15436 36128 16804 36156
rect 15436 36116 15442 36128
rect 6914 36048 6920 36100
rect 6972 36048 6978 36100
rect 7650 36048 7656 36100
rect 7708 36048 7714 36100
rect 9861 36091 9919 36097
rect 9861 36057 9873 36091
rect 9907 36088 9919 36091
rect 14274 36088 14280 36100
rect 9907 36060 14280 36088
rect 9907 36057 9919 36060
rect 9861 36051 9919 36057
rect 14274 36048 14280 36060
rect 14332 36048 14338 36100
rect 14645 36091 14703 36097
rect 14645 36057 14657 36091
rect 14691 36088 14703 36091
rect 15473 36091 15531 36097
rect 15473 36088 15485 36091
rect 14691 36060 15485 36088
rect 14691 36057 14703 36060
rect 14645 36051 14703 36057
rect 15473 36057 15485 36060
rect 15519 36057 15531 36091
rect 16776 36088 16804 36128
rect 16850 36116 16856 36168
rect 16908 36156 16914 36168
rect 17497 36159 17555 36165
rect 17497 36156 17509 36159
rect 16908 36128 17509 36156
rect 16908 36116 16914 36128
rect 17497 36125 17509 36128
rect 17543 36125 17555 36159
rect 17497 36119 17555 36125
rect 21082 36116 21088 36168
rect 21140 36156 21146 36168
rect 21177 36159 21235 36165
rect 21177 36156 21189 36159
rect 21140 36128 21189 36156
rect 21140 36116 21146 36128
rect 21177 36125 21189 36128
rect 21223 36125 21235 36159
rect 21177 36119 21235 36125
rect 19797 36091 19855 36097
rect 19797 36088 19809 36091
rect 16776 36060 19809 36088
rect 15473 36051 15531 36057
rect 19797 36057 19809 36060
rect 19843 36088 19855 36091
rect 22066 36088 22094 36332
rect 25038 36320 25044 36332
rect 25096 36320 25102 36372
rect 24670 36252 24676 36304
rect 24728 36292 24734 36304
rect 24728 36264 25176 36292
rect 24728 36252 24734 36264
rect 22278 36184 22284 36236
rect 22336 36224 22342 36236
rect 24946 36224 24952 36236
rect 22336 36196 24952 36224
rect 22336 36184 22342 36196
rect 24946 36184 24952 36196
rect 25004 36184 25010 36236
rect 25148 36233 25176 36264
rect 25133 36227 25191 36233
rect 25133 36193 25145 36227
rect 25179 36193 25191 36227
rect 25133 36187 25191 36193
rect 23842 36116 23848 36168
rect 23900 36156 23906 36168
rect 25041 36159 25099 36165
rect 25041 36156 25053 36159
rect 23900 36128 25053 36156
rect 23900 36116 23906 36128
rect 25041 36125 25053 36128
rect 25087 36125 25099 36159
rect 25041 36119 25099 36125
rect 19843 36060 22094 36088
rect 22557 36091 22615 36097
rect 19843 36057 19855 36060
rect 19797 36051 19855 36057
rect 22557 36057 22569 36091
rect 22603 36088 22615 36091
rect 22646 36088 22652 36100
rect 22603 36060 22652 36088
rect 22603 36057 22615 36060
rect 22557 36051 22615 36057
rect 22646 36048 22652 36060
rect 22704 36048 22710 36100
rect 23566 36048 23572 36100
rect 23624 36048 23630 36100
rect 23934 36048 23940 36100
rect 23992 36088 23998 36100
rect 24949 36091 25007 36097
rect 24949 36088 24961 36091
rect 23992 36060 24961 36088
rect 23992 36048 23998 36060
rect 24949 36057 24961 36060
rect 24995 36057 25007 36091
rect 24949 36051 25007 36057
rect 1765 36023 1823 36029
rect 1765 35989 1777 36023
rect 1811 36020 1823 36023
rect 4154 36020 4160 36032
rect 1811 35992 4160 36020
rect 1811 35989 1823 35992
rect 1765 35983 1823 35989
rect 4154 35980 4160 35992
rect 4212 35980 4218 36032
rect 11333 36023 11391 36029
rect 11333 35989 11345 36023
rect 11379 36020 11391 36023
rect 11790 36020 11796 36032
rect 11379 35992 11796 36020
rect 11379 35989 11391 35992
rect 11333 35983 11391 35989
rect 11790 35980 11796 35992
rect 11848 35980 11854 36032
rect 12250 35980 12256 36032
rect 12308 36020 12314 36032
rect 12710 36020 12716 36032
rect 12308 35992 12716 36020
rect 12308 35980 12314 35992
rect 12710 35980 12716 35992
rect 12768 35980 12774 36032
rect 12894 35980 12900 36032
rect 12952 36020 12958 36032
rect 13909 36023 13967 36029
rect 13909 36020 13921 36023
rect 12952 35992 13921 36020
rect 12952 35980 12958 35992
rect 13909 35989 13921 35992
rect 13955 36020 13967 36023
rect 14553 36023 14611 36029
rect 14553 36020 14565 36023
rect 13955 35992 14565 36020
rect 13955 35989 13967 35992
rect 13909 35983 13967 35989
rect 14553 35989 14565 35992
rect 14599 35989 14611 36023
rect 14553 35983 14611 35989
rect 15194 35980 15200 36032
rect 15252 36020 15258 36032
rect 15378 36020 15384 36032
rect 15252 35992 15384 36020
rect 15252 35980 15258 35992
rect 15378 35980 15384 35992
rect 15436 35980 15442 36032
rect 18141 36023 18199 36029
rect 18141 35989 18153 36023
rect 18187 36020 18199 36023
rect 18414 36020 18420 36032
rect 18187 35992 18420 36020
rect 18187 35989 18199 35992
rect 18141 35983 18199 35989
rect 18414 35980 18420 35992
rect 18472 35980 18478 36032
rect 19429 36023 19487 36029
rect 19429 35989 19441 36023
rect 19475 36020 19487 36023
rect 19610 36020 19616 36032
rect 19475 35992 19616 36020
rect 19475 35989 19487 35992
rect 19429 35983 19487 35989
rect 19610 35980 19616 35992
rect 19668 35980 19674 36032
rect 20809 36023 20867 36029
rect 20809 35989 20821 36023
rect 20855 36020 20867 36023
rect 20898 36020 20904 36032
rect 20855 35992 20904 36020
rect 20855 35989 20867 35992
rect 20809 35983 20867 35989
rect 20898 35980 20904 35992
rect 20956 35980 20962 36032
rect 24029 36023 24087 36029
rect 24029 35989 24041 36023
rect 24075 36020 24087 36023
rect 24486 36020 24492 36032
rect 24075 35992 24492 36020
rect 24075 35989 24087 35992
rect 24029 35983 24087 35989
rect 24486 35980 24492 35992
rect 24544 35980 24550 36032
rect 24578 35980 24584 36032
rect 24636 35980 24642 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 6546 35816 6552 35828
rect 4264 35788 6552 35816
rect 4264 35689 4292 35788
rect 6546 35776 6552 35788
rect 6604 35776 6610 35828
rect 6914 35776 6920 35828
rect 6972 35816 6978 35828
rect 7377 35819 7435 35825
rect 7377 35816 7389 35819
rect 6972 35788 7389 35816
rect 6972 35776 6978 35788
rect 7377 35785 7389 35788
rect 7423 35785 7435 35819
rect 10318 35816 10324 35828
rect 7377 35779 7435 35785
rect 8496 35788 10324 35816
rect 5902 35748 5908 35760
rect 5750 35720 5908 35748
rect 5902 35708 5908 35720
rect 5960 35748 5966 35760
rect 6457 35751 6515 35757
rect 6457 35748 6469 35751
rect 5960 35720 6469 35748
rect 5960 35708 5966 35720
rect 6457 35717 6469 35720
rect 6503 35748 6515 35751
rect 8294 35748 8300 35760
rect 6503 35720 8300 35748
rect 6503 35717 6515 35720
rect 6457 35711 6515 35717
rect 8294 35708 8300 35720
rect 8352 35708 8358 35760
rect 8496 35689 8524 35788
rect 10318 35776 10324 35788
rect 10376 35776 10382 35828
rect 11698 35776 11704 35828
rect 11756 35776 11762 35828
rect 13817 35819 13875 35825
rect 13817 35816 13829 35819
rect 12084 35788 13829 35816
rect 9766 35708 9772 35760
rect 9824 35708 9830 35760
rect 12084 35692 12112 35788
rect 13817 35785 13829 35788
rect 13863 35816 13875 35819
rect 13906 35816 13912 35828
rect 13863 35788 13912 35816
rect 13863 35785 13875 35788
rect 13817 35779 13875 35785
rect 13906 35776 13912 35788
rect 13964 35776 13970 35828
rect 19426 35816 19432 35828
rect 17880 35788 19432 35816
rect 13446 35708 13452 35760
rect 13504 35748 13510 35760
rect 17494 35748 17500 35760
rect 13504 35720 17500 35748
rect 13504 35708 13510 35720
rect 17494 35708 17500 35720
rect 17552 35708 17558 35760
rect 4249 35683 4307 35689
rect 4249 35649 4261 35683
rect 4295 35649 4307 35683
rect 4249 35643 4307 35649
rect 8021 35683 8079 35689
rect 8021 35649 8033 35683
rect 8067 35649 8079 35683
rect 8021 35643 8079 35649
rect 8481 35683 8539 35689
rect 8481 35649 8493 35683
rect 8527 35649 8539 35683
rect 8481 35643 8539 35649
rect 4522 35572 4528 35624
rect 4580 35572 4586 35624
rect 5994 35572 6000 35624
rect 6052 35572 6058 35624
rect 7006 35436 7012 35488
rect 7064 35436 7070 35488
rect 8036 35476 8064 35643
rect 10686 35640 10692 35692
rect 10744 35680 10750 35692
rect 12066 35680 12072 35692
rect 10744 35652 12072 35680
rect 10744 35640 10750 35652
rect 12066 35640 12072 35652
rect 12124 35640 12130 35692
rect 17218 35640 17224 35692
rect 17276 35680 17282 35692
rect 17880 35689 17908 35788
rect 19426 35776 19432 35788
rect 19484 35776 19490 35828
rect 23658 35776 23664 35828
rect 23716 35816 23722 35828
rect 23716 35788 24348 35816
rect 23716 35776 23722 35788
rect 18141 35751 18199 35757
rect 18141 35717 18153 35751
rect 18187 35748 18199 35751
rect 18414 35748 18420 35760
rect 18187 35720 18420 35748
rect 18187 35717 18199 35720
rect 18141 35711 18199 35717
rect 18414 35708 18420 35720
rect 18472 35708 18478 35760
rect 24320 35748 24348 35788
rect 24394 35748 24400 35760
rect 24242 35720 24400 35748
rect 24394 35708 24400 35720
rect 24452 35708 24458 35760
rect 17865 35683 17923 35689
rect 17865 35680 17877 35683
rect 17276 35652 17877 35680
rect 17276 35640 17282 35652
rect 17865 35649 17877 35652
rect 17911 35649 17923 35683
rect 17865 35643 17923 35649
rect 19242 35640 19248 35692
rect 19300 35640 19306 35692
rect 8754 35572 8760 35624
rect 8812 35572 8818 35624
rect 8846 35572 8852 35624
rect 8904 35612 8910 35624
rect 12526 35612 12532 35624
rect 8904 35584 12532 35612
rect 8904 35572 8910 35584
rect 12526 35572 12532 35584
rect 12584 35572 12590 35624
rect 13173 35615 13231 35621
rect 13173 35581 13185 35615
rect 13219 35612 13231 35615
rect 13219 35584 13400 35612
rect 13219 35581 13231 35584
rect 13173 35575 13231 35581
rect 10244 35516 11836 35544
rect 10244 35485 10272 35516
rect 10229 35479 10287 35485
rect 10229 35476 10241 35479
rect 8036 35448 10241 35476
rect 10229 35445 10241 35448
rect 10275 35445 10287 35479
rect 11808 35476 11836 35516
rect 13372 35488 13400 35584
rect 13446 35572 13452 35624
rect 13504 35572 13510 35624
rect 17770 35572 17776 35624
rect 17828 35612 17834 35624
rect 17828 35584 22094 35612
rect 17828 35572 17834 35584
rect 22066 35544 22094 35584
rect 22646 35572 22652 35624
rect 22704 35572 22710 35624
rect 24026 35612 24032 35624
rect 22756 35584 24032 35612
rect 22756 35544 22784 35584
rect 24026 35572 24032 35584
rect 24084 35572 24090 35624
rect 24670 35572 24676 35624
rect 24728 35572 24734 35624
rect 24946 35572 24952 35624
rect 25004 35572 25010 35624
rect 25130 35572 25136 35624
rect 25188 35612 25194 35624
rect 25317 35615 25375 35621
rect 25317 35612 25329 35615
rect 25188 35584 25329 35612
rect 25188 35572 25194 35584
rect 25317 35581 25329 35584
rect 25363 35612 25375 35615
rect 25590 35612 25596 35624
rect 25363 35584 25596 35612
rect 25363 35581 25375 35584
rect 25317 35575 25375 35581
rect 25590 35572 25596 35584
rect 25648 35572 25654 35624
rect 22066 35516 22784 35544
rect 12434 35476 12440 35488
rect 11808 35448 12440 35476
rect 10229 35439 10287 35445
rect 12434 35436 12440 35448
rect 12492 35436 12498 35488
rect 13354 35436 13360 35488
rect 13412 35436 13418 35488
rect 16298 35436 16304 35488
rect 16356 35476 16362 35488
rect 18322 35476 18328 35488
rect 16356 35448 18328 35476
rect 16356 35436 16362 35448
rect 18322 35436 18328 35448
rect 18380 35436 18386 35488
rect 19613 35479 19671 35485
rect 19613 35445 19625 35479
rect 19659 35476 19671 35479
rect 22002 35476 22008 35488
rect 19659 35448 22008 35476
rect 19659 35445 19671 35448
rect 19613 35439 19671 35445
rect 22002 35436 22008 35448
rect 22060 35436 22066 35488
rect 22462 35436 22468 35488
rect 22520 35476 22526 35488
rect 23201 35479 23259 35485
rect 23201 35476 23213 35479
rect 22520 35448 23213 35476
rect 22520 35436 22526 35448
rect 23201 35445 23213 35448
rect 23247 35445 23259 35479
rect 23201 35439 23259 35445
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 4522 35232 4528 35284
rect 4580 35272 4586 35284
rect 5537 35275 5595 35281
rect 5537 35272 5549 35275
rect 4580 35244 5549 35272
rect 4580 35232 4586 35244
rect 5537 35241 5549 35244
rect 5583 35272 5595 35275
rect 5583 35244 7512 35272
rect 5583 35241 5595 35244
rect 5537 35235 5595 35241
rect 7484 35204 7512 35244
rect 7742 35232 7748 35284
rect 7800 35272 7806 35284
rect 7837 35275 7895 35281
rect 7837 35272 7849 35275
rect 7800 35244 7849 35272
rect 7800 35232 7806 35244
rect 7837 35241 7849 35244
rect 7883 35241 7895 35275
rect 7837 35235 7895 35241
rect 8294 35232 8300 35284
rect 8352 35272 8358 35284
rect 8938 35272 8944 35284
rect 8352 35244 8944 35272
rect 8352 35232 8358 35244
rect 8938 35232 8944 35244
rect 8996 35232 9002 35284
rect 9309 35275 9367 35281
rect 9309 35241 9321 35275
rect 9355 35272 9367 35275
rect 9490 35272 9496 35284
rect 9355 35244 9496 35272
rect 9355 35241 9367 35244
rect 9309 35235 9367 35241
rect 9490 35232 9496 35244
rect 9548 35232 9554 35284
rect 12618 35272 12624 35284
rect 9784 35244 12624 35272
rect 9582 35204 9588 35216
rect 7484 35176 9588 35204
rect 9582 35164 9588 35176
rect 9640 35164 9646 35216
rect 6546 35096 6552 35148
rect 6604 35136 6610 35148
rect 7285 35139 7343 35145
rect 7285 35136 7297 35139
rect 6604 35108 7297 35136
rect 6604 35096 6610 35108
rect 7285 35105 7297 35108
rect 7331 35105 7343 35139
rect 7285 35099 7343 35105
rect 7558 35096 7564 35148
rect 7616 35136 7622 35148
rect 9784 35145 9812 35244
rect 12618 35232 12624 35244
rect 12676 35232 12682 35284
rect 13081 35275 13139 35281
rect 13081 35241 13093 35275
rect 13127 35272 13139 35275
rect 13354 35272 13360 35284
rect 13127 35244 13360 35272
rect 13127 35241 13139 35244
rect 13081 35235 13139 35241
rect 13354 35232 13360 35244
rect 13412 35232 13418 35284
rect 15473 35275 15531 35281
rect 15473 35241 15485 35275
rect 15519 35272 15531 35275
rect 15654 35272 15660 35284
rect 15519 35244 15660 35272
rect 15519 35241 15531 35244
rect 15473 35235 15531 35241
rect 15654 35232 15660 35244
rect 15712 35232 15718 35284
rect 17494 35232 17500 35284
rect 17552 35272 17558 35284
rect 19150 35272 19156 35284
rect 17552 35244 19156 35272
rect 17552 35232 17558 35244
rect 19150 35232 19156 35244
rect 19208 35232 19214 35284
rect 19242 35232 19248 35284
rect 19300 35272 19306 35284
rect 19300 35244 20852 35272
rect 19300 35232 19306 35244
rect 20824 35204 20852 35244
rect 23934 35232 23940 35284
rect 23992 35232 23998 35284
rect 24670 35232 24676 35284
rect 24728 35272 24734 35284
rect 25225 35275 25283 35281
rect 25225 35272 25237 35275
rect 24728 35244 25237 35272
rect 24728 35232 24734 35244
rect 25225 35241 25237 35244
rect 25271 35241 25283 35275
rect 25225 35235 25283 35241
rect 23566 35204 23572 35216
rect 20824 35176 23572 35204
rect 8389 35139 8447 35145
rect 8389 35136 8401 35139
rect 7616 35108 8401 35136
rect 7616 35096 7622 35108
rect 8389 35105 8401 35108
rect 8435 35105 8447 35139
rect 8389 35099 8447 35105
rect 9769 35139 9827 35145
rect 9769 35105 9781 35139
rect 9815 35105 9827 35139
rect 9769 35099 9827 35105
rect 9953 35139 10011 35145
rect 9953 35105 9965 35139
rect 9999 35136 10011 35139
rect 10042 35136 10048 35148
rect 9999 35108 10048 35136
rect 9999 35105 10011 35108
rect 9953 35099 10011 35105
rect 10042 35096 10048 35108
rect 10100 35096 10106 35148
rect 10318 35096 10324 35148
rect 10376 35136 10382 35148
rect 12345 35139 12403 35145
rect 12345 35136 12357 35139
rect 10376 35108 12357 35136
rect 10376 35096 10382 35108
rect 12345 35105 12357 35108
rect 12391 35136 12403 35139
rect 13446 35136 13452 35148
rect 12391 35108 13452 35136
rect 12391 35105 12403 35108
rect 12345 35099 12403 35105
rect 13446 35096 13452 35108
rect 13504 35096 13510 35148
rect 15654 35096 15660 35148
rect 15712 35136 15718 35148
rect 17218 35136 17224 35148
rect 15712 35108 17224 35136
rect 15712 35096 15718 35108
rect 17218 35096 17224 35108
rect 17276 35096 17282 35148
rect 18414 35136 18420 35148
rect 18248 35108 18420 35136
rect 5902 35028 5908 35080
rect 5960 35028 5966 35080
rect 8297 35071 8355 35077
rect 8297 35037 8309 35071
rect 8343 35068 8355 35071
rect 10778 35068 10784 35080
rect 8343 35040 10784 35068
rect 8343 35037 8355 35040
rect 8297 35031 8355 35037
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 18248 35077 18276 35108
rect 18414 35096 18420 35108
rect 18472 35136 18478 35148
rect 20254 35136 20260 35148
rect 18472 35108 20260 35136
rect 18472 35096 18478 35108
rect 20254 35096 20260 35108
rect 20312 35096 20318 35148
rect 13725 35071 13783 35077
rect 13725 35037 13737 35071
rect 13771 35037 13783 35071
rect 13725 35031 13783 35037
rect 18233 35071 18291 35077
rect 18233 35037 18245 35071
rect 18279 35037 18291 35071
rect 18233 35031 18291 35037
rect 7006 34960 7012 35012
rect 7064 34960 7070 35012
rect 8205 35003 8263 35009
rect 8205 34969 8217 35003
rect 8251 34969 8263 35003
rect 8205 34963 8263 34969
rect 8220 34932 8248 34963
rect 8938 34960 8944 35012
rect 8996 35000 9002 35012
rect 10686 35000 10692 35012
rect 8996 34972 10692 35000
rect 8996 34960 9002 34972
rect 10686 34960 10692 34972
rect 10744 35000 10750 35012
rect 10744 34972 10902 35000
rect 10744 34960 10750 34972
rect 11790 34960 11796 35012
rect 11848 35000 11854 35012
rect 12069 35003 12127 35009
rect 12069 35000 12081 35003
rect 11848 34972 12081 35000
rect 11848 34960 11854 34972
rect 12069 34969 12081 34972
rect 12115 34969 12127 35003
rect 12069 34963 12127 34969
rect 13446 34960 13452 35012
rect 13504 35000 13510 35012
rect 13740 35000 13768 35031
rect 19334 35028 19340 35080
rect 19392 35068 19398 35080
rect 19429 35071 19487 35077
rect 19429 35068 19441 35071
rect 19392 35040 19441 35068
rect 19392 35028 19398 35040
rect 19429 35037 19441 35040
rect 19475 35037 19487 35071
rect 20824 35054 20852 35176
rect 23566 35164 23572 35176
rect 23624 35164 23630 35216
rect 22186 35096 22192 35148
rect 22244 35096 22250 35148
rect 23385 35139 23443 35145
rect 23385 35105 23397 35139
rect 23431 35136 23443 35139
rect 24118 35136 24124 35148
rect 23431 35108 24124 35136
rect 23431 35105 23443 35108
rect 23385 35099 23443 35105
rect 24118 35096 24124 35108
rect 24176 35096 24182 35148
rect 19429 35031 19487 35037
rect 20990 35028 20996 35080
rect 21048 35068 21054 35080
rect 22373 35071 22431 35077
rect 22373 35068 22385 35071
rect 21048 35040 22385 35068
rect 21048 35028 21054 35040
rect 22373 35037 22385 35040
rect 22419 35037 22431 35071
rect 22373 35031 22431 35037
rect 22646 35028 22652 35080
rect 22704 35068 22710 35080
rect 23569 35071 23627 35077
rect 23569 35068 23581 35071
rect 22704 35040 23581 35068
rect 22704 35028 22710 35040
rect 23569 35037 23581 35040
rect 23615 35037 23627 35071
rect 23569 35031 23627 35037
rect 24026 35028 24032 35080
rect 24084 35068 24090 35080
rect 24486 35068 24492 35080
rect 24084 35040 24492 35068
rect 24084 35028 24090 35040
rect 24486 35028 24492 35040
rect 24544 35068 24550 35080
rect 24581 35071 24639 35077
rect 24581 35068 24593 35071
rect 24544 35040 24593 35068
rect 24544 35028 24550 35040
rect 24581 35037 24593 35040
rect 24627 35037 24639 35071
rect 24581 35031 24639 35037
rect 16945 35003 17003 35009
rect 13504 34972 13768 35000
rect 16514 34972 16896 35000
rect 13504 34960 13510 34972
rect 8294 34932 8300 34944
rect 8220 34904 8300 34932
rect 8294 34892 8300 34904
rect 8352 34892 8358 34944
rect 9674 34892 9680 34944
rect 9732 34892 9738 34944
rect 10597 34935 10655 34941
rect 10597 34901 10609 34935
rect 10643 34932 10655 34935
rect 11698 34932 11704 34944
rect 10643 34904 11704 34932
rect 10643 34901 10655 34904
rect 10597 34895 10655 34901
rect 11698 34892 11704 34904
rect 11756 34892 11762 34944
rect 12710 34892 12716 34944
rect 12768 34932 12774 34944
rect 14093 34935 14151 34941
rect 14093 34932 14105 34935
rect 12768 34904 14105 34932
rect 12768 34892 12774 34904
rect 14093 34901 14105 34904
rect 14139 34901 14151 34935
rect 16868 34932 16896 34972
rect 16945 34969 16957 35003
rect 16991 35000 17003 35003
rect 17218 35000 17224 35012
rect 16991 34972 17224 35000
rect 16991 34969 17003 34972
rect 16945 34963 17003 34969
rect 17218 34960 17224 34972
rect 17276 34960 17282 35012
rect 18877 35003 18935 35009
rect 18877 34969 18889 35003
rect 18923 35000 18935 35003
rect 19705 35003 19763 35009
rect 19705 35000 19717 35003
rect 18923 34972 19717 35000
rect 18923 34969 18935 34972
rect 18877 34963 18935 34969
rect 19705 34969 19717 34972
rect 19751 34969 19763 35003
rect 19705 34963 19763 34969
rect 21082 34960 21088 35012
rect 21140 35000 21146 35012
rect 23477 35003 23535 35009
rect 23477 35000 23489 35003
rect 21140 34972 23489 35000
rect 21140 34960 21146 34972
rect 23477 34969 23489 34972
rect 23523 34969 23535 35003
rect 23477 34963 23535 34969
rect 19242 34932 19248 34944
rect 16868 34904 19248 34932
rect 14093 34895 14151 34901
rect 19242 34892 19248 34904
rect 19300 34892 19306 34944
rect 21174 34892 21180 34944
rect 21232 34892 21238 34944
rect 22281 34935 22339 34941
rect 22281 34901 22293 34935
rect 22327 34932 22339 34935
rect 22646 34932 22652 34944
rect 22327 34904 22652 34932
rect 22327 34901 22339 34904
rect 22281 34895 22339 34901
rect 22646 34892 22652 34904
rect 22704 34892 22710 34944
rect 22738 34892 22744 34944
rect 22796 34892 22802 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 4890 34688 4896 34740
rect 4948 34728 4954 34740
rect 5537 34731 5595 34737
rect 5537 34728 5549 34731
rect 4948 34700 5549 34728
rect 4948 34688 4954 34700
rect 5537 34697 5549 34700
rect 5583 34697 5595 34731
rect 5537 34691 5595 34697
rect 5997 34731 6055 34737
rect 5997 34697 6009 34731
rect 6043 34728 6055 34731
rect 6086 34728 6092 34740
rect 6043 34700 6092 34728
rect 6043 34697 6055 34700
rect 5997 34691 6055 34697
rect 5552 34660 5580 34691
rect 6086 34688 6092 34700
rect 6144 34688 6150 34740
rect 7650 34688 7656 34740
rect 7708 34728 7714 34740
rect 7708 34700 7972 34728
rect 7708 34688 7714 34700
rect 6730 34660 6736 34672
rect 5552 34632 6736 34660
rect 6730 34620 6736 34632
rect 6788 34620 6794 34672
rect 5626 34552 5632 34604
rect 5684 34552 5690 34604
rect 7944 34592 7972 34700
rect 8570 34688 8576 34740
rect 8628 34728 8634 34740
rect 8849 34731 8907 34737
rect 8849 34728 8861 34731
rect 8628 34700 8861 34728
rect 8628 34688 8634 34700
rect 8849 34697 8861 34700
rect 8895 34728 8907 34731
rect 9306 34728 9312 34740
rect 8895 34700 9312 34728
rect 8895 34697 8907 34700
rect 8849 34691 8907 34697
rect 9306 34688 9312 34700
rect 9364 34688 9370 34740
rect 10965 34731 11023 34737
rect 10965 34697 10977 34731
rect 11011 34728 11023 34731
rect 11054 34728 11060 34740
rect 11011 34700 11060 34728
rect 11011 34697 11023 34700
rect 10965 34691 11023 34697
rect 11054 34688 11060 34700
rect 11112 34688 11118 34740
rect 11146 34688 11152 34740
rect 11204 34728 11210 34740
rect 11241 34731 11299 34737
rect 11241 34728 11253 34731
rect 11204 34700 11253 34728
rect 11204 34688 11210 34700
rect 11241 34697 11253 34700
rect 11287 34728 11299 34731
rect 11422 34728 11428 34740
rect 11287 34700 11428 34728
rect 11287 34697 11299 34700
rect 11241 34691 11299 34697
rect 11422 34688 11428 34700
rect 11480 34688 11486 34740
rect 12066 34688 12072 34740
rect 12124 34728 12130 34740
rect 12710 34728 12716 34740
rect 12124 34700 12716 34728
rect 12124 34688 12130 34700
rect 10318 34620 10324 34672
rect 10376 34660 10382 34672
rect 11072 34660 11100 34688
rect 11514 34660 11520 34672
rect 10376 34632 10640 34660
rect 11072 34632 11520 34660
rect 10376 34620 10382 34632
rect 10612 34601 10640 34632
rect 11514 34620 11520 34632
rect 11572 34620 11578 34672
rect 11974 34620 11980 34672
rect 12032 34620 12038 34672
rect 12406 34660 12434 34700
rect 12710 34688 12716 34700
rect 12768 34688 12774 34740
rect 13630 34688 13636 34740
rect 13688 34728 13694 34740
rect 13909 34731 13967 34737
rect 13909 34728 13921 34731
rect 13688 34700 13921 34728
rect 13688 34688 13694 34700
rect 13909 34697 13921 34700
rect 13955 34697 13967 34731
rect 13909 34691 13967 34697
rect 14369 34731 14427 34737
rect 14369 34697 14381 34731
rect 14415 34728 14427 34731
rect 14734 34728 14740 34740
rect 14415 34700 14740 34728
rect 14415 34697 14427 34700
rect 14369 34691 14427 34697
rect 14734 34688 14740 34700
rect 14792 34688 14798 34740
rect 17218 34688 17224 34740
rect 17276 34688 17282 34740
rect 18325 34731 18383 34737
rect 18325 34697 18337 34731
rect 18371 34697 18383 34731
rect 18325 34691 18383 34697
rect 12406 34632 12466 34660
rect 17034 34620 17040 34672
rect 17092 34660 17098 34672
rect 18340 34660 18368 34691
rect 18598 34688 18604 34740
rect 18656 34728 18662 34740
rect 18693 34731 18751 34737
rect 18693 34728 18705 34731
rect 18656 34700 18705 34728
rect 18656 34688 18662 34700
rect 18693 34697 18705 34700
rect 18739 34697 18751 34731
rect 18693 34691 18751 34697
rect 20625 34731 20683 34737
rect 20625 34697 20637 34731
rect 20671 34728 20683 34731
rect 22465 34731 22523 34737
rect 20671 34700 22094 34728
rect 20671 34697 20683 34700
rect 20625 34691 20683 34697
rect 17092 34632 18368 34660
rect 17092 34620 17098 34632
rect 21818 34620 21824 34672
rect 21876 34620 21882 34672
rect 22066 34660 22094 34700
rect 22465 34697 22477 34731
rect 22511 34728 22523 34731
rect 22554 34728 22560 34740
rect 22511 34700 22560 34728
rect 22511 34697 22523 34700
rect 22465 34691 22523 34697
rect 22554 34688 22560 34700
rect 22612 34688 22618 34740
rect 22646 34688 22652 34740
rect 22704 34728 22710 34740
rect 22830 34728 22836 34740
rect 22704 34700 22836 34728
rect 22704 34688 22710 34700
rect 22830 34688 22836 34700
rect 22888 34728 22894 34740
rect 23201 34731 23259 34737
rect 23201 34728 23213 34731
rect 22888 34700 23213 34728
rect 22888 34688 22894 34700
rect 23201 34697 23213 34700
rect 23247 34697 23259 34731
rect 23201 34691 23259 34697
rect 23937 34731 23995 34737
rect 23937 34697 23949 34731
rect 23983 34728 23995 34731
rect 24394 34728 24400 34740
rect 23983 34700 24400 34728
rect 23983 34697 23995 34700
rect 23937 34691 23995 34697
rect 24394 34688 24400 34700
rect 24452 34688 24458 34740
rect 24581 34731 24639 34737
rect 24581 34697 24593 34731
rect 24627 34728 24639 34731
rect 24762 34728 24768 34740
rect 24627 34700 24768 34728
rect 24627 34697 24639 34700
rect 24581 34691 24639 34697
rect 24762 34688 24768 34700
rect 24820 34688 24826 34740
rect 22066 34632 22600 34660
rect 10597 34595 10655 34601
rect 7944 34578 9246 34592
rect 7958 34564 9260 34578
rect 5445 34527 5503 34533
rect 5445 34493 5457 34527
rect 5491 34524 5503 34527
rect 5491 34496 5580 34524
rect 5491 34493 5503 34496
rect 5445 34487 5503 34493
rect 5552 34468 5580 34496
rect 5810 34484 5816 34536
rect 5868 34524 5874 34536
rect 6546 34524 6552 34536
rect 5868 34496 6552 34524
rect 5868 34484 5874 34496
rect 6546 34484 6552 34496
rect 6604 34484 6610 34536
rect 6822 34484 6828 34536
rect 6880 34484 6886 34536
rect 8297 34527 8355 34533
rect 8297 34493 8309 34527
rect 8343 34524 8355 34527
rect 8846 34524 8852 34536
rect 8343 34496 8852 34524
rect 8343 34493 8355 34496
rect 8297 34487 8355 34493
rect 8846 34484 8852 34496
rect 8904 34484 8910 34536
rect 9232 34524 9260 34564
rect 10597 34561 10609 34595
rect 10643 34592 10655 34595
rect 11701 34595 11759 34601
rect 11701 34592 11713 34595
rect 10643 34564 11713 34592
rect 10643 34561 10655 34564
rect 10597 34555 10655 34561
rect 11701 34561 11713 34564
rect 11747 34561 11759 34595
rect 13630 34592 13636 34604
rect 11701 34555 11759 34561
rect 13188 34564 13636 34592
rect 9766 34524 9772 34536
rect 9232 34496 9772 34524
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 10321 34527 10379 34533
rect 10321 34493 10333 34527
rect 10367 34524 10379 34527
rect 10367 34496 10548 34524
rect 10367 34493 10379 34496
rect 10321 34487 10379 34493
rect 5534 34416 5540 34468
rect 5592 34416 5598 34468
rect 10520 34456 10548 34496
rect 11146 34484 11152 34536
rect 11204 34524 11210 34536
rect 12342 34524 12348 34536
rect 11204 34496 12348 34524
rect 11204 34484 11210 34496
rect 12342 34484 12348 34496
rect 12400 34484 12406 34536
rect 12526 34484 12532 34536
rect 12584 34524 12590 34536
rect 13188 34524 13216 34564
rect 13630 34552 13636 34564
rect 13688 34552 13694 34604
rect 14277 34595 14335 34601
rect 14277 34561 14289 34595
rect 14323 34592 14335 34595
rect 17865 34595 17923 34601
rect 14323 34564 17632 34592
rect 14323 34561 14335 34564
rect 14277 34555 14335 34561
rect 12584 34496 13216 34524
rect 12584 34484 12590 34496
rect 13446 34484 13452 34536
rect 13504 34484 13510 34536
rect 14461 34527 14519 34533
rect 14461 34493 14473 34527
rect 14507 34493 14519 34527
rect 14461 34487 14519 34493
rect 11054 34456 11060 34468
rect 10520 34428 11060 34456
rect 11054 34416 11060 34428
rect 11112 34456 11118 34468
rect 14476 34456 14504 34487
rect 11112 34428 11376 34456
rect 11112 34416 11118 34428
rect 11348 34388 11376 34428
rect 13372 34428 14504 34456
rect 17604 34456 17632 34564
rect 17865 34561 17877 34595
rect 17911 34592 17923 34595
rect 18322 34592 18328 34604
rect 17911 34564 18328 34592
rect 17911 34561 17923 34564
rect 17865 34555 17923 34561
rect 18322 34552 18328 34564
rect 18380 34552 18386 34604
rect 19337 34595 19395 34601
rect 19337 34592 19349 34595
rect 18800 34564 19349 34592
rect 17770 34484 17776 34536
rect 17828 34524 17834 34536
rect 18800 34533 18828 34564
rect 19337 34561 19349 34564
rect 19383 34561 19395 34595
rect 19337 34555 19395 34561
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19521 34595 19579 34601
rect 19521 34592 19533 34595
rect 19484 34564 19533 34592
rect 19484 34552 19490 34564
rect 19521 34561 19533 34564
rect 19567 34592 19579 34595
rect 20165 34595 20223 34601
rect 20165 34592 20177 34595
rect 19567 34564 20177 34592
rect 19567 34561 19579 34564
rect 19521 34555 19579 34561
rect 20165 34561 20177 34564
rect 20211 34561 20223 34595
rect 20165 34555 20223 34561
rect 20254 34552 20260 34604
rect 20312 34552 20318 34604
rect 20806 34552 20812 34604
rect 20864 34592 20870 34604
rect 22370 34592 22376 34604
rect 20864 34564 22376 34592
rect 20864 34552 20870 34564
rect 22370 34552 22376 34564
rect 22428 34552 22434 34604
rect 22572 34601 22600 34632
rect 22557 34595 22615 34601
rect 22557 34561 22569 34595
rect 22603 34561 22615 34595
rect 22557 34555 22615 34561
rect 23753 34595 23811 34601
rect 23753 34561 23765 34595
rect 23799 34592 23811 34595
rect 24210 34592 24216 34604
rect 23799 34564 24216 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 24210 34552 24216 34564
rect 24268 34552 24274 34604
rect 24302 34552 24308 34604
rect 24360 34592 24366 34604
rect 24397 34595 24455 34601
rect 24397 34592 24409 34595
rect 24360 34564 24409 34592
rect 24360 34552 24366 34564
rect 24397 34561 24409 34564
rect 24443 34561 24455 34595
rect 24397 34555 24455 34561
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 18785 34527 18843 34533
rect 18785 34524 18797 34527
rect 17828 34496 18797 34524
rect 17828 34484 17834 34496
rect 18785 34493 18797 34496
rect 18831 34493 18843 34527
rect 18785 34487 18843 34493
rect 18877 34527 18935 34533
rect 18877 34493 18889 34527
rect 18923 34493 18935 34527
rect 18877 34487 18935 34493
rect 20073 34527 20131 34533
rect 20073 34493 20085 34527
rect 20119 34493 20131 34527
rect 20073 34487 20131 34493
rect 18598 34456 18604 34468
rect 17604 34428 18604 34456
rect 13372 34388 13400 34428
rect 18598 34416 18604 34428
rect 18656 34416 18662 34468
rect 18690 34416 18696 34468
rect 18748 34456 18754 34468
rect 18892 34456 18920 34487
rect 18748 34428 18920 34456
rect 20088 34456 20116 34487
rect 20714 34484 20720 34536
rect 20772 34524 20778 34536
rect 20901 34527 20959 34533
rect 20901 34524 20913 34527
rect 20772 34496 20913 34524
rect 20772 34484 20778 34496
rect 20901 34493 20913 34496
rect 20947 34493 20959 34527
rect 20901 34487 20959 34493
rect 22281 34527 22339 34533
rect 22281 34493 22293 34527
rect 22327 34493 22339 34527
rect 23658 34524 23664 34536
rect 22281 34487 22339 34493
rect 22940 34496 23664 34524
rect 22094 34456 22100 34468
rect 20088 34428 22100 34456
rect 18748 34416 18754 34428
rect 22094 34416 22100 34428
rect 22152 34416 22158 34468
rect 11348 34360 13400 34388
rect 22296 34388 22324 34487
rect 22940 34465 22968 34496
rect 23658 34484 23664 34496
rect 23716 34484 23722 34536
rect 22925 34459 22983 34465
rect 22925 34425 22937 34459
rect 22971 34425 22983 34459
rect 22925 34419 22983 34425
rect 24026 34388 24032 34400
rect 22296 34360 24032 34388
rect 24026 34348 24032 34360
rect 24084 34348 24090 34400
rect 25130 34348 25136 34400
rect 25188 34348 25194 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 6822 34144 6828 34196
rect 6880 34184 6886 34196
rect 7101 34187 7159 34193
rect 7101 34184 7113 34187
rect 6880 34156 7113 34184
rect 6880 34144 6886 34156
rect 7101 34153 7113 34156
rect 7147 34153 7159 34187
rect 7101 34147 7159 34153
rect 7929 34187 7987 34193
rect 7929 34153 7941 34187
rect 7975 34184 7987 34187
rect 8754 34184 8760 34196
rect 7975 34156 8760 34184
rect 7975 34153 7987 34156
rect 7929 34147 7987 34153
rect 8754 34144 8760 34156
rect 8812 34144 8818 34196
rect 9122 34144 9128 34196
rect 9180 34144 9186 34196
rect 9766 34144 9772 34196
rect 9824 34184 9830 34196
rect 10413 34187 10471 34193
rect 10413 34184 10425 34187
rect 9824 34156 10425 34184
rect 9824 34144 9830 34156
rect 10413 34153 10425 34156
rect 10459 34153 10471 34187
rect 10413 34147 10471 34153
rect 11057 34187 11115 34193
rect 11057 34153 11069 34187
rect 11103 34184 11115 34187
rect 11238 34184 11244 34196
rect 11103 34156 11244 34184
rect 11103 34153 11115 34156
rect 11057 34147 11115 34153
rect 11238 34144 11244 34156
rect 11296 34144 11302 34196
rect 11514 34144 11520 34196
rect 11572 34184 11578 34196
rect 14182 34184 14188 34196
rect 11572 34156 14188 34184
rect 11572 34144 11578 34156
rect 14182 34144 14188 34156
rect 14240 34144 14246 34196
rect 14274 34144 14280 34196
rect 14332 34144 14338 34196
rect 17313 34187 17371 34193
rect 17313 34153 17325 34187
rect 17359 34184 17371 34187
rect 18414 34184 18420 34196
rect 17359 34156 18420 34184
rect 17359 34153 17371 34156
rect 17313 34147 17371 34153
rect 18414 34144 18420 34156
rect 18472 34144 18478 34196
rect 20349 34187 20407 34193
rect 20349 34153 20361 34187
rect 20395 34184 20407 34187
rect 21082 34184 21088 34196
rect 20395 34156 21088 34184
rect 20395 34153 20407 34156
rect 20349 34147 20407 34153
rect 21082 34144 21088 34156
rect 21140 34144 21146 34196
rect 21358 34144 21364 34196
rect 21416 34184 21422 34196
rect 23845 34187 23903 34193
rect 23845 34184 23857 34187
rect 21416 34156 23857 34184
rect 21416 34144 21422 34156
rect 23845 34153 23857 34156
rect 23891 34153 23903 34187
rect 23845 34147 23903 34153
rect 24489 34187 24547 34193
rect 24489 34153 24501 34187
rect 24535 34184 24547 34187
rect 24854 34184 24860 34196
rect 24535 34156 24860 34184
rect 24535 34153 24547 34156
rect 24489 34147 24547 34153
rect 11882 34116 11888 34128
rect 11624 34088 11888 34116
rect 5626 34008 5632 34060
rect 5684 34048 5690 34060
rect 5813 34051 5871 34057
rect 5813 34048 5825 34051
rect 5684 34020 5825 34048
rect 5684 34008 5690 34020
rect 5813 34017 5825 34020
rect 5859 34017 5871 34051
rect 5813 34011 5871 34017
rect 9582 34008 9588 34060
rect 9640 34048 9646 34060
rect 9677 34051 9735 34057
rect 9677 34048 9689 34051
rect 9640 34020 9689 34048
rect 9640 34008 9646 34020
rect 9677 34017 9689 34020
rect 9723 34017 9735 34051
rect 9677 34011 9735 34017
rect 11514 34008 11520 34060
rect 11572 34008 11578 34060
rect 11624 34057 11652 34088
rect 11882 34076 11888 34088
rect 11940 34076 11946 34128
rect 12434 34076 12440 34128
rect 12492 34116 12498 34128
rect 12492 34088 14872 34116
rect 12492 34076 12498 34088
rect 11609 34051 11667 34057
rect 11609 34017 11621 34051
rect 11655 34017 11667 34051
rect 11609 34011 11667 34017
rect 11698 34008 11704 34060
rect 11756 34048 11762 34060
rect 14844 34057 14872 34088
rect 16850 34076 16856 34128
rect 16908 34116 16914 34128
rect 19702 34116 19708 34128
rect 16908 34088 19708 34116
rect 16908 34076 16914 34088
rect 19702 34076 19708 34088
rect 19760 34076 19766 34128
rect 22462 34116 22468 34128
rect 19812 34088 22468 34116
rect 13541 34051 13599 34057
rect 13541 34048 13553 34051
rect 11756 34020 13553 34048
rect 11756 34008 11762 34020
rect 13541 34017 13553 34020
rect 13587 34017 13599 34051
rect 13541 34011 13599 34017
rect 14829 34051 14887 34057
rect 14829 34017 14841 34051
rect 14875 34017 14887 34051
rect 19242 34048 19248 34060
rect 14829 34011 14887 34017
rect 16960 34020 19248 34048
rect 5994 33940 6000 33992
rect 6052 33980 6058 33992
rect 6457 33983 6515 33989
rect 6457 33980 6469 33983
rect 6052 33952 6469 33980
rect 6052 33940 6058 33952
rect 6457 33949 6469 33952
rect 6503 33949 6515 33983
rect 6457 33943 6515 33949
rect 8570 33940 8576 33992
rect 8628 33940 8634 33992
rect 10597 33983 10655 33989
rect 10597 33949 10609 33983
rect 10643 33980 10655 33983
rect 11146 33980 11152 33992
rect 10643 33952 11152 33980
rect 10643 33949 10655 33952
rect 10597 33943 10655 33949
rect 11146 33940 11152 33952
rect 11204 33940 11210 33992
rect 11238 33940 11244 33992
rect 11296 33980 11302 33992
rect 11716 33980 11744 34008
rect 11296 33952 11744 33980
rect 11296 33940 11302 33952
rect 15562 33940 15568 33992
rect 15620 33940 15626 33992
rect 16850 33940 16856 33992
rect 16908 33980 16914 33992
rect 16960 33980 16988 34020
rect 19242 34008 19248 34020
rect 19300 34008 19306 34060
rect 19812 34057 19840 34088
rect 22462 34076 22468 34088
rect 22520 34076 22526 34128
rect 19797 34051 19855 34057
rect 19797 34017 19809 34051
rect 19843 34017 19855 34051
rect 21358 34048 21364 34060
rect 19797 34011 19855 34017
rect 21192 34020 21364 34048
rect 20990 33980 20996 33992
rect 16908 33966 16988 33980
rect 16908 33952 16974 33966
rect 17696 33952 20996 33980
rect 16908 33940 16914 33952
rect 9585 33915 9643 33921
rect 9585 33881 9597 33915
rect 9631 33912 9643 33915
rect 12158 33912 12164 33924
rect 9631 33884 12164 33912
rect 9631 33881 9643 33884
rect 9585 33875 9643 33881
rect 12158 33872 12164 33884
rect 12216 33872 12222 33924
rect 13449 33915 13507 33921
rect 13449 33881 13461 33915
rect 13495 33912 13507 33915
rect 13538 33912 13544 33924
rect 13495 33884 13544 33912
rect 13495 33881 13507 33884
rect 13449 33875 13507 33881
rect 13538 33872 13544 33884
rect 13596 33872 13602 33924
rect 15102 33872 15108 33924
rect 15160 33912 15166 33924
rect 15841 33915 15899 33921
rect 15841 33912 15853 33915
rect 15160 33884 15853 33912
rect 15160 33872 15166 33884
rect 15841 33881 15853 33884
rect 15887 33881 15899 33915
rect 15841 33875 15899 33881
rect 7834 33804 7840 33856
rect 7892 33844 7898 33856
rect 9493 33847 9551 33853
rect 9493 33844 9505 33847
rect 7892 33816 9505 33844
rect 7892 33804 7898 33816
rect 9493 33813 9505 33816
rect 9539 33813 9551 33847
rect 9493 33807 9551 33813
rect 11422 33804 11428 33856
rect 11480 33804 11486 33856
rect 12710 33804 12716 33856
rect 12768 33844 12774 33856
rect 12989 33847 13047 33853
rect 12989 33844 13001 33847
rect 12768 33816 13001 33844
rect 12768 33804 12774 33816
rect 12989 33813 13001 33816
rect 13035 33813 13047 33847
rect 12989 33807 13047 33813
rect 13354 33804 13360 33856
rect 13412 33804 13418 33856
rect 14090 33804 14096 33856
rect 14148 33844 14154 33856
rect 14645 33847 14703 33853
rect 14645 33844 14657 33847
rect 14148 33816 14657 33844
rect 14148 33804 14154 33816
rect 14645 33813 14657 33816
rect 14691 33813 14703 33847
rect 14645 33807 14703 33813
rect 14737 33847 14795 33853
rect 14737 33813 14749 33847
rect 14783 33844 14795 33847
rect 17696 33844 17724 33952
rect 20990 33940 20996 33952
rect 21048 33980 21054 33992
rect 21192 33980 21220 34020
rect 21358 34008 21364 34020
rect 21416 34008 21422 34060
rect 21450 34008 21456 34060
rect 21508 34008 21514 34060
rect 21048 33952 21220 33980
rect 21269 33983 21327 33989
rect 21048 33940 21054 33952
rect 21269 33949 21281 33983
rect 21315 33980 21327 33983
rect 21818 33980 21824 33992
rect 21315 33952 21824 33980
rect 21315 33949 21327 33952
rect 21269 33943 21327 33949
rect 21818 33940 21824 33952
rect 21876 33940 21882 33992
rect 22002 33940 22008 33992
rect 22060 33940 22066 33992
rect 24029 33983 24087 33989
rect 24029 33949 24041 33983
rect 24075 33980 24087 33983
rect 24504 33980 24532 34147
rect 24854 34144 24860 34156
rect 24912 34144 24918 34196
rect 24075 33952 24532 33980
rect 24857 33983 24915 33989
rect 24075 33949 24087 33952
rect 24029 33943 24087 33949
rect 24857 33949 24869 33983
rect 24903 33980 24915 33983
rect 25317 33983 25375 33989
rect 25317 33980 25329 33983
rect 24903 33952 25329 33980
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 25317 33949 25329 33952
rect 25363 33980 25375 33983
rect 25406 33980 25412 33992
rect 25363 33952 25412 33980
rect 25363 33949 25375 33952
rect 25317 33943 25375 33949
rect 25406 33940 25412 33952
rect 25464 33940 25470 33992
rect 19981 33915 20039 33921
rect 19981 33912 19993 33915
rect 19352 33884 19993 33912
rect 14783 33816 17724 33844
rect 14783 33813 14795 33816
rect 14737 33807 14795 33813
rect 17770 33804 17776 33856
rect 17828 33844 17834 33856
rect 19352 33853 19380 33884
rect 19981 33881 19993 33884
rect 20027 33881 20039 33915
rect 19981 33875 20039 33881
rect 21177 33915 21235 33921
rect 21177 33881 21189 33915
rect 21223 33912 21235 33915
rect 21726 33912 21732 33924
rect 21223 33884 21732 33912
rect 21223 33881 21235 33884
rect 21177 33875 21235 33881
rect 21726 33872 21732 33884
rect 21784 33872 21790 33924
rect 22462 33872 22468 33924
rect 22520 33912 22526 33924
rect 22520 33884 25176 33912
rect 22520 33872 22526 33884
rect 19337 33847 19395 33853
rect 19337 33844 19349 33847
rect 17828 33816 19349 33844
rect 17828 33804 17834 33816
rect 19337 33813 19349 33816
rect 19383 33813 19395 33847
rect 19337 33807 19395 33813
rect 19886 33804 19892 33856
rect 19944 33844 19950 33856
rect 20714 33844 20720 33856
rect 19944 33816 20720 33844
rect 19944 33804 19950 33816
rect 20714 33804 20720 33816
rect 20772 33804 20778 33856
rect 20806 33804 20812 33856
rect 20864 33804 20870 33856
rect 22646 33804 22652 33856
rect 22704 33804 22710 33856
rect 23106 33804 23112 33856
rect 23164 33804 23170 33856
rect 23198 33804 23204 33856
rect 23256 33844 23262 33856
rect 23474 33844 23480 33856
rect 23256 33816 23480 33844
rect 23256 33804 23262 33816
rect 23474 33804 23480 33816
rect 23532 33804 23538 33856
rect 25148 33853 25176 33884
rect 25133 33847 25191 33853
rect 25133 33813 25145 33847
rect 25179 33813 25191 33847
rect 25133 33807 25191 33813
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 6178 33600 6184 33652
rect 6236 33640 6242 33652
rect 7650 33640 7656 33652
rect 6236 33612 7656 33640
rect 6236 33600 6242 33612
rect 7650 33600 7656 33612
rect 7708 33640 7714 33652
rect 8297 33643 8355 33649
rect 8297 33640 8309 33643
rect 7708 33612 8309 33640
rect 7708 33600 7714 33612
rect 8297 33609 8309 33612
rect 8343 33609 8355 33643
rect 8297 33603 8355 33609
rect 8757 33643 8815 33649
rect 8757 33609 8769 33643
rect 8803 33640 8815 33643
rect 9674 33640 9680 33652
rect 8803 33612 9680 33640
rect 8803 33609 8815 33612
rect 8757 33603 8815 33609
rect 9674 33600 9680 33612
rect 9732 33600 9738 33652
rect 10505 33643 10563 33649
rect 10505 33609 10517 33643
rect 10551 33640 10563 33643
rect 10870 33640 10876 33652
rect 10551 33612 10876 33640
rect 10551 33609 10563 33612
rect 10505 33603 10563 33609
rect 10870 33600 10876 33612
rect 10928 33600 10934 33652
rect 11701 33643 11759 33649
rect 11701 33609 11713 33643
rect 11747 33609 11759 33643
rect 11701 33603 11759 33609
rect 12161 33643 12219 33649
rect 12161 33609 12173 33643
rect 12207 33640 12219 33643
rect 12250 33640 12256 33652
rect 12207 33612 12256 33640
rect 12207 33609 12219 33612
rect 12161 33603 12219 33609
rect 10778 33532 10784 33584
rect 10836 33572 10842 33584
rect 11716 33572 11744 33603
rect 12250 33600 12256 33612
rect 12308 33600 12314 33652
rect 15102 33600 15108 33652
rect 15160 33600 15166 33652
rect 16025 33643 16083 33649
rect 16025 33609 16037 33643
rect 16071 33640 16083 33643
rect 17402 33640 17408 33652
rect 16071 33612 17408 33640
rect 16071 33609 16083 33612
rect 16025 33603 16083 33609
rect 17402 33600 17408 33612
rect 17460 33600 17466 33652
rect 19610 33640 19616 33652
rect 17696 33612 19616 33640
rect 10836 33544 11744 33572
rect 15933 33575 15991 33581
rect 10836 33532 10842 33544
rect 15933 33541 15945 33575
rect 15979 33572 15991 33575
rect 17696 33572 17724 33612
rect 19610 33600 19616 33612
rect 19668 33600 19674 33652
rect 19702 33600 19708 33652
rect 19760 33640 19766 33652
rect 22373 33643 22431 33649
rect 19760 33612 22324 33640
rect 19760 33600 19766 33612
rect 19242 33572 19248 33584
rect 15979 33544 17724 33572
rect 19090 33544 19248 33572
rect 15979 33541 15991 33544
rect 15933 33535 15991 33541
rect 19242 33532 19248 33544
rect 19300 33532 19306 33584
rect 19521 33575 19579 33581
rect 19521 33541 19533 33575
rect 19567 33572 19579 33575
rect 20441 33575 20499 33581
rect 20441 33572 20453 33575
rect 19567 33544 20453 33572
rect 19567 33541 19579 33544
rect 19521 33535 19579 33541
rect 20441 33541 20453 33544
rect 20487 33541 20499 33575
rect 22296 33572 22324 33612
rect 22373 33609 22385 33643
rect 22419 33640 22431 33643
rect 23106 33640 23112 33652
rect 22419 33612 23112 33640
rect 22419 33609 22431 33612
rect 22373 33603 22431 33609
rect 23106 33600 23112 33612
rect 23164 33600 23170 33652
rect 25222 33600 25228 33652
rect 25280 33600 25286 33652
rect 23842 33572 23848 33584
rect 22296 33544 23848 33572
rect 20441 33535 20499 33541
rect 23842 33532 23848 33544
rect 23900 33532 23906 33584
rect 24486 33532 24492 33584
rect 24544 33532 24550 33584
rect 1210 33464 1216 33516
rect 1268 33504 1274 33516
rect 1581 33507 1639 33513
rect 1581 33504 1593 33507
rect 1268 33476 1593 33504
rect 1268 33464 1274 33476
rect 1581 33473 1593 33476
rect 1627 33504 1639 33507
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1627 33476 2053 33504
rect 1627 33473 1639 33476
rect 1581 33467 1639 33473
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 8386 33464 8392 33516
rect 8444 33464 8450 33516
rect 10137 33507 10195 33513
rect 10137 33473 10149 33507
rect 10183 33504 10195 33507
rect 10965 33507 11023 33513
rect 10965 33504 10977 33507
rect 10183 33476 10977 33504
rect 10183 33473 10195 33476
rect 10137 33467 10195 33473
rect 10965 33473 10977 33476
rect 11011 33473 11023 33507
rect 10965 33467 11023 33473
rect 11422 33464 11428 33516
rect 11480 33504 11486 33516
rect 11790 33504 11796 33516
rect 11480 33476 11796 33504
rect 11480 33464 11486 33476
rect 11790 33464 11796 33476
rect 11848 33464 11854 33516
rect 12069 33507 12127 33513
rect 12069 33473 12081 33507
rect 12115 33504 12127 33507
rect 14274 33504 14280 33516
rect 12115 33476 14280 33504
rect 12115 33473 12127 33476
rect 12069 33467 12127 33473
rect 14274 33464 14280 33476
rect 14332 33464 14338 33516
rect 14458 33464 14464 33516
rect 14516 33464 14522 33516
rect 16942 33504 16948 33516
rect 15212 33476 16948 33504
rect 15212 33448 15240 33476
rect 16942 33464 16948 33476
rect 17000 33464 17006 33516
rect 21085 33507 21143 33513
rect 21085 33473 21097 33507
rect 21131 33504 21143 33507
rect 21174 33504 21180 33516
rect 21131 33476 21180 33504
rect 21131 33473 21143 33476
rect 21085 33467 21143 33473
rect 21174 33464 21180 33476
rect 21232 33504 21238 33516
rect 21232 33476 22600 33504
rect 21232 33464 21238 33476
rect 8205 33439 8263 33445
rect 8205 33405 8217 33439
rect 8251 33436 8263 33439
rect 9030 33436 9036 33448
rect 8251 33408 9036 33436
rect 8251 33405 8263 33408
rect 8205 33399 8263 33405
rect 9030 33396 9036 33408
rect 9088 33396 9094 33448
rect 9861 33439 9919 33445
rect 9861 33405 9873 33439
rect 9907 33405 9919 33439
rect 9861 33399 9919 33405
rect 7098 33328 7104 33380
rect 7156 33368 7162 33380
rect 9876 33368 9904 33399
rect 9950 33396 9956 33448
rect 10008 33436 10014 33448
rect 10045 33439 10103 33445
rect 10045 33436 10057 33439
rect 10008 33408 10057 33436
rect 10008 33396 10014 33408
rect 10045 33405 10057 33408
rect 10091 33405 10103 33439
rect 10045 33399 10103 33405
rect 12253 33439 12311 33445
rect 12253 33405 12265 33439
rect 12299 33405 12311 33439
rect 12253 33399 12311 33405
rect 11054 33368 11060 33380
rect 7156 33340 9168 33368
rect 9876 33340 11060 33368
rect 7156 33328 7162 33340
rect 1765 33303 1823 33309
rect 1765 33269 1777 33303
rect 1811 33300 1823 33303
rect 3878 33300 3884 33312
rect 1811 33272 3884 33300
rect 1811 33269 1823 33272
rect 1765 33263 1823 33269
rect 3878 33260 3884 33272
rect 3936 33260 3942 33312
rect 9030 33260 9036 33312
rect 9088 33260 9094 33312
rect 9140 33300 9168 33340
rect 11054 33328 11060 33340
rect 11112 33328 11118 33380
rect 12268 33300 12296 33399
rect 12342 33396 12348 33448
rect 12400 33436 12406 33448
rect 15194 33436 15200 33448
rect 12400 33408 15200 33436
rect 12400 33396 12406 33408
rect 15194 33396 15200 33408
rect 15252 33396 15258 33448
rect 16114 33396 16120 33448
rect 16172 33396 16178 33448
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 19797 33439 19855 33445
rect 19797 33436 19809 33439
rect 19484 33408 19809 33436
rect 19484 33396 19490 33408
rect 19797 33405 19809 33408
rect 19843 33405 19855 33439
rect 19797 33399 19855 33405
rect 20346 33396 20352 33448
rect 20404 33436 20410 33448
rect 22462 33436 22468 33448
rect 20404 33408 22468 33436
rect 20404 33396 20410 33408
rect 22462 33396 22468 33408
rect 22520 33396 22526 33448
rect 22572 33445 22600 33476
rect 22557 33439 22615 33445
rect 22557 33405 22569 33439
rect 22603 33405 22615 33439
rect 22557 33399 22615 33405
rect 23290 33396 23296 33448
rect 23348 33436 23354 33448
rect 23477 33439 23535 33445
rect 23477 33436 23489 33439
rect 23348 33408 23489 33436
rect 23348 33396 23354 33408
rect 23477 33405 23489 33408
rect 23523 33405 23535 33439
rect 23477 33399 23535 33405
rect 13354 33328 13360 33380
rect 13412 33368 13418 33380
rect 13909 33371 13967 33377
rect 13909 33368 13921 33371
rect 13412 33340 13921 33368
rect 13412 33328 13418 33340
rect 13909 33337 13921 33340
rect 13955 33368 13967 33371
rect 17678 33368 17684 33380
rect 13955 33340 17684 33368
rect 13955 33337 13967 33340
rect 13909 33331 13967 33337
rect 17678 33328 17684 33340
rect 17736 33328 17742 33380
rect 21818 33328 21824 33380
rect 21876 33368 21882 33380
rect 23017 33371 23075 33377
rect 23017 33368 23029 33371
rect 21876 33340 23029 33368
rect 21876 33328 21882 33340
rect 23017 33337 23029 33340
rect 23063 33368 23075 33371
rect 23198 33368 23204 33380
rect 23063 33340 23204 33368
rect 23063 33337 23075 33340
rect 23017 33331 23075 33337
rect 23198 33328 23204 33340
rect 23256 33328 23262 33380
rect 9140 33272 12296 33300
rect 14090 33260 14096 33312
rect 14148 33260 14154 33312
rect 15562 33260 15568 33312
rect 15620 33260 15626 33312
rect 15930 33260 15936 33312
rect 15988 33300 15994 33312
rect 16390 33300 16396 33312
rect 15988 33272 16396 33300
rect 15988 33260 15994 33272
rect 16390 33260 16396 33272
rect 16448 33260 16454 33312
rect 18049 33303 18107 33309
rect 18049 33269 18061 33303
rect 18095 33300 18107 33303
rect 18322 33300 18328 33312
rect 18095 33272 18328 33300
rect 18095 33269 18107 33272
rect 18049 33263 18107 33269
rect 18322 33260 18328 33272
rect 18380 33300 18386 33312
rect 18966 33300 18972 33312
rect 18380 33272 18972 33300
rect 18380 33260 18386 33272
rect 18966 33260 18972 33272
rect 19024 33260 19030 33312
rect 20714 33260 20720 33312
rect 20772 33300 20778 33312
rect 22005 33303 22063 33309
rect 22005 33300 22017 33303
rect 20772 33272 22017 33300
rect 20772 33260 20778 33272
rect 22005 33269 22017 33272
rect 22051 33269 22063 33303
rect 22005 33263 22063 33269
rect 22278 33260 22284 33312
rect 22336 33300 22342 33312
rect 22554 33300 22560 33312
rect 22336 33272 22560 33300
rect 22336 33260 22342 33272
rect 22554 33260 22560 33272
rect 22612 33260 22618 33312
rect 23492 33300 23520 33399
rect 23750 33396 23756 33448
rect 23808 33396 23814 33448
rect 24946 33300 24952 33312
rect 23492 33272 24952 33300
rect 24946 33260 24952 33272
rect 25004 33260 25010 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 7558 33056 7564 33108
rect 7616 33056 7622 33108
rect 7929 33099 7987 33105
rect 7929 33065 7941 33099
rect 7975 33096 7987 33099
rect 8938 33096 8944 33108
rect 7975 33068 8944 33096
rect 7975 33065 7987 33068
rect 7929 33059 7987 33065
rect 6089 32963 6147 32969
rect 6089 32929 6101 32963
rect 6135 32960 6147 32963
rect 7098 32960 7104 32972
rect 6135 32932 7104 32960
rect 6135 32929 6147 32932
rect 6089 32923 6147 32929
rect 7098 32920 7104 32932
rect 7156 32920 7162 32972
rect 7944 32960 7972 33059
rect 8938 33056 8944 33068
rect 8996 33096 9002 33108
rect 9674 33096 9680 33108
rect 8996 33068 9680 33096
rect 8996 33056 9002 33068
rect 9674 33056 9680 33068
rect 9732 33056 9738 33108
rect 16206 33056 16212 33108
rect 16264 33096 16270 33108
rect 16393 33099 16451 33105
rect 16393 33096 16405 33099
rect 16264 33068 16405 33096
rect 16264 33056 16270 33068
rect 16393 33065 16405 33068
rect 16439 33096 16451 33099
rect 16439 33068 17172 33096
rect 16439 33065 16451 33068
rect 16393 33059 16451 33065
rect 7208 32932 7972 32960
rect 5810 32852 5816 32904
rect 5868 32852 5874 32904
rect 7208 32878 7236 32932
rect 8386 32920 8392 32972
rect 8444 32920 8450 32972
rect 15654 32920 15660 32972
rect 15712 32960 15718 32972
rect 16945 32963 17003 32969
rect 15712 32932 16068 32960
rect 15712 32920 15718 32932
rect 7558 32852 7564 32904
rect 7616 32892 7622 32904
rect 16040 32901 16068 32932
rect 16945 32929 16957 32963
rect 16991 32960 17003 32963
rect 16991 32932 17080 32960
rect 16991 32929 17003 32932
rect 16945 32923 17003 32929
rect 9125 32895 9183 32901
rect 9125 32892 9137 32895
rect 7616 32864 9137 32892
rect 7616 32852 7622 32864
rect 9125 32861 9137 32864
rect 9171 32861 9183 32895
rect 9125 32855 9183 32861
rect 16025 32895 16083 32901
rect 16025 32861 16037 32895
rect 16071 32892 16083 32895
rect 16666 32892 16672 32904
rect 16071 32864 16672 32892
rect 16071 32861 16083 32864
rect 16025 32855 16083 32861
rect 16666 32852 16672 32864
rect 16724 32852 16730 32904
rect 10962 32784 10968 32836
rect 11020 32824 11026 32836
rect 12802 32824 12808 32836
rect 11020 32796 12808 32824
rect 11020 32784 11026 32796
rect 12802 32784 12808 32796
rect 12860 32784 12866 32836
rect 15318 32796 15608 32824
rect 8294 32716 8300 32768
rect 8352 32756 8358 32768
rect 9769 32759 9827 32765
rect 9769 32756 9781 32759
rect 8352 32728 9781 32756
rect 8352 32716 8358 32728
rect 9769 32725 9781 32728
rect 9815 32725 9827 32759
rect 9769 32719 9827 32725
rect 14182 32716 14188 32768
rect 14240 32756 14246 32768
rect 14277 32759 14335 32765
rect 14277 32756 14289 32759
rect 14240 32728 14289 32756
rect 14240 32716 14246 32728
rect 14277 32725 14289 32728
rect 14323 32725 14335 32759
rect 14277 32719 14335 32725
rect 14826 32716 14832 32768
rect 14884 32756 14890 32768
rect 15102 32756 15108 32768
rect 14884 32728 15108 32756
rect 14884 32716 14890 32728
rect 15102 32716 15108 32728
rect 15160 32716 15166 32768
rect 15580 32756 15608 32796
rect 15654 32784 15660 32836
rect 15712 32824 15718 32836
rect 15749 32827 15807 32833
rect 15749 32824 15761 32827
rect 15712 32796 15761 32824
rect 15712 32784 15718 32796
rect 15749 32793 15761 32796
rect 15795 32793 15807 32827
rect 17052 32824 17080 32932
rect 17144 32901 17172 33068
rect 17218 33056 17224 33108
rect 17276 33096 17282 33108
rect 17678 33096 17684 33108
rect 17276 33068 17684 33096
rect 17276 33056 17282 33068
rect 17678 33056 17684 33068
rect 17736 33096 17742 33108
rect 17773 33099 17831 33105
rect 17773 33096 17785 33099
rect 17736 33068 17785 33096
rect 17736 33056 17742 33068
rect 17773 33065 17785 33068
rect 17819 33065 17831 33099
rect 17773 33059 17831 33065
rect 18506 33056 18512 33108
rect 18564 33096 18570 33108
rect 18874 33096 18880 33108
rect 18564 33068 18880 33096
rect 18564 33056 18570 33068
rect 18874 33056 18880 33068
rect 18932 33056 18938 33108
rect 23474 33056 23480 33108
rect 23532 33056 23538 33108
rect 23842 33056 23848 33108
rect 23900 33056 23906 33108
rect 25038 33056 25044 33108
rect 25096 33096 25102 33108
rect 25133 33099 25191 33105
rect 25133 33096 25145 33099
rect 25096 33068 25145 33096
rect 25096 33056 25102 33068
rect 25133 33065 25145 33068
rect 25179 33065 25191 33099
rect 25133 33059 25191 33065
rect 17402 32988 17408 33040
rect 17460 33028 17466 33040
rect 19886 33028 19892 33040
rect 17460 33000 19892 33028
rect 17460 32988 17466 33000
rect 19886 32988 19892 33000
rect 19944 33028 19950 33040
rect 20625 33031 20683 33037
rect 19944 33000 20576 33028
rect 19944 32988 19950 33000
rect 17494 32920 17500 32972
rect 17552 32960 17558 32972
rect 19610 32960 19616 32972
rect 17552 32932 19616 32960
rect 17552 32920 17558 32932
rect 19610 32920 19616 32932
rect 19668 32920 19674 32972
rect 19981 32963 20039 32969
rect 19981 32929 19993 32963
rect 20027 32960 20039 32963
rect 20254 32960 20260 32972
rect 20027 32932 20260 32960
rect 20027 32929 20039 32932
rect 19981 32923 20039 32929
rect 20254 32920 20260 32932
rect 20312 32920 20318 32972
rect 17129 32895 17187 32901
rect 17129 32861 17141 32895
rect 17175 32861 17187 32895
rect 17129 32855 17187 32861
rect 17586 32852 17592 32904
rect 17644 32892 17650 32904
rect 20441 32895 20499 32901
rect 20441 32892 20453 32895
rect 17644 32864 20453 32892
rect 17644 32852 17650 32864
rect 20441 32861 20453 32864
rect 20487 32861 20499 32895
rect 20441 32855 20499 32861
rect 20346 32824 20352 32836
rect 17052 32796 20352 32824
rect 15749 32787 15807 32793
rect 20346 32784 20352 32796
rect 20404 32784 20410 32836
rect 20548 32824 20576 33000
rect 20625 32997 20637 33031
rect 20671 33028 20683 33031
rect 22094 33028 22100 33040
rect 20671 33000 22100 33028
rect 20671 32997 20683 33000
rect 20625 32991 20683 32997
rect 22094 32988 22100 33000
rect 22152 32988 22158 33040
rect 22278 32988 22284 33040
rect 22336 33028 22342 33040
rect 23017 33031 23075 33037
rect 23017 33028 23029 33031
rect 22336 33000 23029 33028
rect 22336 32988 22342 33000
rect 23017 32997 23029 33000
rect 23063 32997 23075 33031
rect 23017 32991 23075 32997
rect 21082 32920 21088 32972
rect 21140 32960 21146 32972
rect 21361 32963 21419 32969
rect 21361 32960 21373 32963
rect 21140 32932 21373 32960
rect 21140 32920 21146 32932
rect 21361 32929 21373 32932
rect 21407 32960 21419 32963
rect 22002 32960 22008 32972
rect 21407 32932 22008 32960
rect 21407 32929 21419 32932
rect 21361 32923 21419 32929
rect 22002 32920 22008 32932
rect 22060 32920 22066 32972
rect 23492 32960 23520 33056
rect 22112 32932 23520 32960
rect 21453 32895 21511 32901
rect 21453 32861 21465 32895
rect 21499 32892 21511 32895
rect 21726 32892 21732 32904
rect 21499 32864 21732 32892
rect 21499 32861 21511 32864
rect 21453 32855 21511 32861
rect 21726 32852 21732 32864
rect 21784 32892 21790 32904
rect 22112 32892 22140 32932
rect 21784 32864 22140 32892
rect 21784 32852 21790 32864
rect 22370 32852 22376 32904
rect 22428 32852 22434 32904
rect 22830 32852 22836 32904
rect 22888 32892 22894 32904
rect 23201 32895 23259 32901
rect 23201 32892 23213 32895
rect 22888 32864 23213 32892
rect 22888 32852 22894 32864
rect 23201 32861 23213 32864
rect 23247 32861 23259 32895
rect 23201 32855 23259 32861
rect 24029 32895 24087 32901
rect 24029 32861 24041 32895
rect 24075 32892 24087 32895
rect 24857 32895 24915 32901
rect 24075 32864 24532 32892
rect 24075 32861 24087 32864
rect 24029 32855 24087 32861
rect 21545 32827 21603 32833
rect 21545 32824 21557 32827
rect 20548 32796 21557 32824
rect 21545 32793 21557 32796
rect 21591 32824 21603 32827
rect 21818 32824 21824 32836
rect 21591 32796 21824 32824
rect 21591 32793 21603 32796
rect 21545 32787 21603 32793
rect 21818 32784 21824 32796
rect 21876 32784 21882 32836
rect 24118 32824 24124 32836
rect 22572 32796 24124 32824
rect 16574 32756 16580 32768
rect 15580 32728 16580 32756
rect 16574 32716 16580 32728
rect 16632 32716 16638 32768
rect 17037 32759 17095 32765
rect 17037 32725 17049 32759
rect 17083 32756 17095 32759
rect 17218 32756 17224 32768
rect 17083 32728 17224 32756
rect 17083 32725 17095 32728
rect 17037 32719 17095 32725
rect 17218 32716 17224 32728
rect 17276 32716 17282 32768
rect 17494 32716 17500 32768
rect 17552 32716 17558 32768
rect 19334 32716 19340 32768
rect 19392 32756 19398 32768
rect 19794 32756 19800 32768
rect 19392 32728 19800 32756
rect 19392 32716 19398 32728
rect 19794 32716 19800 32728
rect 19852 32716 19858 32768
rect 21913 32759 21971 32765
rect 21913 32725 21925 32759
rect 21959 32756 21971 32759
rect 22370 32756 22376 32768
rect 21959 32728 22376 32756
rect 21959 32725 21971 32728
rect 21913 32719 21971 32725
rect 22370 32716 22376 32728
rect 22428 32716 22434 32768
rect 22572 32765 22600 32796
rect 24118 32784 24124 32796
rect 24176 32784 24182 32836
rect 24504 32833 24532 32864
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 25314 32892 25320 32904
rect 24903 32864 25320 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 24489 32827 24547 32833
rect 24489 32793 24501 32827
rect 24535 32824 24547 32827
rect 24946 32824 24952 32836
rect 24535 32796 24952 32824
rect 24535 32793 24547 32796
rect 24489 32787 24547 32793
rect 24946 32784 24952 32796
rect 25004 32784 25010 32836
rect 22557 32759 22615 32765
rect 22557 32725 22569 32759
rect 22603 32725 22615 32759
rect 22557 32719 22615 32725
rect 24670 32716 24676 32768
rect 24728 32716 24734 32768
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 12069 32555 12127 32561
rect 12069 32521 12081 32555
rect 12115 32552 12127 32555
rect 12621 32555 12679 32561
rect 12621 32552 12633 32555
rect 12115 32524 12633 32552
rect 12115 32521 12127 32524
rect 12069 32515 12127 32521
rect 12621 32521 12633 32524
rect 12667 32552 12679 32555
rect 12802 32552 12808 32564
rect 12667 32524 12808 32552
rect 12667 32521 12679 32524
rect 12621 32515 12679 32521
rect 12802 32512 12808 32524
rect 12860 32512 12866 32564
rect 13081 32555 13139 32561
rect 13081 32521 13093 32555
rect 13127 32552 13139 32555
rect 14461 32555 14519 32561
rect 14461 32552 14473 32555
rect 13127 32524 14473 32552
rect 13127 32521 13139 32524
rect 13081 32515 13139 32521
rect 14461 32521 14473 32524
rect 14507 32521 14519 32555
rect 14461 32515 14519 32521
rect 15654 32512 15660 32564
rect 15712 32552 15718 32564
rect 17310 32552 17316 32564
rect 15712 32524 17316 32552
rect 15712 32512 15718 32524
rect 17310 32512 17316 32524
rect 17368 32512 17374 32564
rect 17494 32512 17500 32564
rect 17552 32552 17558 32564
rect 18049 32555 18107 32561
rect 18049 32552 18061 32555
rect 17552 32524 18061 32552
rect 17552 32512 17558 32524
rect 18049 32521 18061 32524
rect 18095 32521 18107 32555
rect 18049 32515 18107 32521
rect 18782 32512 18788 32564
rect 18840 32552 18846 32564
rect 20441 32555 20499 32561
rect 18840 32524 20208 32552
rect 18840 32512 18846 32524
rect 8294 32444 8300 32496
rect 8352 32444 8358 32496
rect 9674 32484 9680 32496
rect 9522 32456 9680 32484
rect 9674 32444 9680 32456
rect 9732 32484 9738 32496
rect 10229 32487 10287 32493
rect 10229 32484 10241 32487
rect 9732 32456 10241 32484
rect 9732 32444 9738 32456
rect 10229 32453 10241 32456
rect 10275 32484 10287 32487
rect 10594 32484 10600 32496
rect 10275 32456 10600 32484
rect 10275 32453 10287 32456
rect 10229 32447 10287 32453
rect 10594 32444 10600 32456
rect 10652 32444 10658 32496
rect 14182 32444 14188 32496
rect 14240 32444 14246 32496
rect 14366 32444 14372 32496
rect 14424 32444 14430 32496
rect 14642 32444 14648 32496
rect 14700 32484 14706 32496
rect 17770 32484 17776 32496
rect 14700 32456 17776 32484
rect 14700 32444 14706 32456
rect 17770 32444 17776 32456
rect 17828 32444 17834 32496
rect 17957 32487 18015 32493
rect 17957 32453 17969 32487
rect 18003 32484 18015 32487
rect 19518 32484 19524 32496
rect 18003 32456 19524 32484
rect 18003 32453 18015 32456
rect 17957 32447 18015 32453
rect 19518 32444 19524 32456
rect 19576 32444 19582 32496
rect 5810 32376 5816 32428
rect 5868 32416 5874 32428
rect 12713 32419 12771 32425
rect 5868 32388 8064 32416
rect 5868 32376 5874 32388
rect 8036 32360 8064 32388
rect 12713 32385 12725 32419
rect 12759 32416 12771 32419
rect 12802 32416 12808 32428
rect 12759 32388 12808 32416
rect 12759 32385 12771 32388
rect 12713 32379 12771 32385
rect 12802 32376 12808 32388
rect 12860 32376 12866 32428
rect 13722 32416 13728 32428
rect 13372 32388 13728 32416
rect 7561 32351 7619 32357
rect 7561 32317 7573 32351
rect 7607 32348 7619 32351
rect 7742 32348 7748 32360
rect 7607 32320 7748 32348
rect 7607 32317 7619 32320
rect 7561 32311 7619 32317
rect 7742 32308 7748 32320
rect 7800 32308 7806 32360
rect 8018 32308 8024 32360
rect 8076 32308 8082 32360
rect 9030 32308 9036 32360
rect 9088 32348 9094 32360
rect 11698 32348 11704 32360
rect 9088 32320 11704 32348
rect 9088 32308 9094 32320
rect 11698 32308 11704 32320
rect 11756 32308 11762 32360
rect 12529 32351 12587 32357
rect 12529 32317 12541 32351
rect 12575 32348 12587 32351
rect 13372 32348 13400 32388
rect 13722 32376 13728 32388
rect 13780 32376 13786 32428
rect 14200 32416 14228 32444
rect 15933 32419 15991 32425
rect 15933 32416 15945 32419
rect 14200 32388 15945 32416
rect 15933 32385 15945 32388
rect 15979 32416 15991 32419
rect 16114 32416 16120 32428
rect 15979 32388 16120 32416
rect 15979 32385 15991 32388
rect 15933 32379 15991 32385
rect 16114 32376 16120 32388
rect 16172 32376 16178 32428
rect 16942 32376 16948 32428
rect 17000 32416 17006 32428
rect 17402 32416 17408 32428
rect 17000 32388 17408 32416
rect 17000 32376 17006 32388
rect 17402 32376 17408 32388
rect 17460 32376 17466 32428
rect 19150 32376 19156 32428
rect 19208 32416 19214 32428
rect 19794 32416 19800 32428
rect 19208 32388 19800 32416
rect 19208 32376 19214 32388
rect 19794 32376 19800 32388
rect 19852 32376 19858 32428
rect 20180 32416 20208 32524
rect 20441 32521 20453 32555
rect 20487 32552 20499 32555
rect 20622 32552 20628 32564
rect 20487 32524 20628 32552
rect 20487 32521 20499 32524
rect 20441 32515 20499 32521
rect 20622 32512 20628 32524
rect 20680 32512 20686 32564
rect 21453 32555 21511 32561
rect 21453 32521 21465 32555
rect 21499 32552 21511 32555
rect 21499 32524 22094 32552
rect 21499 32521 21511 32524
rect 21453 32515 21511 32521
rect 20346 32444 20352 32496
rect 20404 32484 20410 32496
rect 21542 32484 21548 32496
rect 20404 32456 21548 32484
rect 20404 32444 20410 32456
rect 21542 32444 21548 32456
rect 21600 32444 21606 32496
rect 22066 32484 22094 32524
rect 22186 32512 22192 32564
rect 22244 32552 22250 32564
rect 22370 32552 22376 32564
rect 22244 32524 22376 32552
rect 22244 32512 22250 32524
rect 22370 32512 22376 32524
rect 22428 32512 22434 32564
rect 22462 32512 22468 32564
rect 22520 32512 22526 32564
rect 23750 32512 23756 32564
rect 23808 32552 23814 32564
rect 24121 32555 24179 32561
rect 24121 32552 24133 32555
rect 23808 32524 24133 32552
rect 23808 32512 23814 32524
rect 24121 32521 24133 32524
rect 24167 32521 24179 32555
rect 24121 32515 24179 32521
rect 23566 32484 23572 32496
rect 22066 32456 23572 32484
rect 23566 32444 23572 32456
rect 23624 32444 23630 32496
rect 21269 32419 21327 32425
rect 21269 32416 21281 32419
rect 20180 32388 21281 32416
rect 21269 32385 21281 32388
rect 21315 32385 21327 32419
rect 21269 32379 21327 32385
rect 22066 32388 22508 32416
rect 12575 32320 13400 32348
rect 12575 32317 12587 32320
rect 12529 32311 12587 32317
rect 13446 32308 13452 32360
rect 13504 32348 13510 32360
rect 14185 32351 14243 32357
rect 14185 32348 14197 32351
rect 13504 32320 14197 32348
rect 13504 32308 13510 32320
rect 14185 32317 14197 32320
rect 14231 32317 14243 32351
rect 14185 32311 14243 32317
rect 17126 32308 17132 32360
rect 17184 32348 17190 32360
rect 18141 32351 18199 32357
rect 18141 32348 18153 32351
rect 17184 32320 18153 32348
rect 17184 32308 17190 32320
rect 18141 32317 18153 32320
rect 18187 32317 18199 32351
rect 18141 32311 18199 32317
rect 19245 32351 19303 32357
rect 19245 32317 19257 32351
rect 19291 32348 19303 32351
rect 19334 32348 19340 32360
rect 19291 32320 19340 32348
rect 19291 32317 19303 32320
rect 19245 32311 19303 32317
rect 19334 32308 19340 32320
rect 19392 32308 19398 32360
rect 19429 32351 19487 32357
rect 19429 32317 19441 32351
rect 19475 32317 19487 32351
rect 19429 32311 19487 32317
rect 9582 32240 9588 32292
rect 9640 32280 9646 32292
rect 9769 32283 9827 32289
rect 9769 32280 9781 32283
rect 9640 32252 9781 32280
rect 9640 32240 9646 32252
rect 9769 32249 9781 32252
rect 9815 32280 9827 32283
rect 15102 32280 15108 32292
rect 9815 32252 15108 32280
rect 9815 32249 9827 32252
rect 9769 32243 9827 32249
rect 15102 32240 15108 32252
rect 15160 32240 15166 32292
rect 16850 32240 16856 32292
rect 16908 32280 16914 32292
rect 17494 32280 17500 32292
rect 16908 32252 17500 32280
rect 16908 32240 16914 32252
rect 17494 32240 17500 32252
rect 17552 32240 17558 32292
rect 18874 32240 18880 32292
rect 18932 32280 18938 32292
rect 19444 32280 19472 32311
rect 20530 32308 20536 32360
rect 20588 32308 20594 32360
rect 21542 32308 21548 32360
rect 21600 32348 21606 32360
rect 21910 32348 21916 32360
rect 21600 32320 21916 32348
rect 21600 32308 21606 32320
rect 21910 32308 21916 32320
rect 21968 32308 21974 32360
rect 18932 32252 19472 32280
rect 18932 32240 18938 32252
rect 19794 32240 19800 32292
rect 19852 32280 19858 32292
rect 19852 32252 20392 32280
rect 19852 32240 19858 32252
rect 6914 32172 6920 32224
rect 6972 32212 6978 32224
rect 7098 32212 7104 32224
rect 6972 32184 7104 32212
rect 6972 32172 6978 32184
rect 7098 32172 7104 32184
rect 7156 32172 7162 32224
rect 7282 32172 7288 32224
rect 7340 32212 7346 32224
rect 10962 32212 10968 32224
rect 7340 32184 10968 32212
rect 7340 32172 7346 32184
rect 10962 32172 10968 32184
rect 11020 32172 11026 32224
rect 14826 32172 14832 32224
rect 14884 32172 14890 32224
rect 14918 32172 14924 32224
rect 14976 32212 14982 32224
rect 15289 32215 15347 32221
rect 15289 32212 15301 32215
rect 14976 32184 15301 32212
rect 14976 32172 14982 32184
rect 15289 32181 15301 32184
rect 15335 32181 15347 32215
rect 15289 32175 15347 32181
rect 17586 32172 17592 32224
rect 17644 32172 17650 32224
rect 18785 32215 18843 32221
rect 18785 32181 18797 32215
rect 18831 32212 18843 32215
rect 19150 32212 19156 32224
rect 18831 32184 19156 32212
rect 18831 32181 18843 32184
rect 18785 32175 18843 32181
rect 19150 32172 19156 32184
rect 19208 32172 19214 32224
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 19981 32215 20039 32221
rect 19981 32212 19993 32215
rect 19392 32184 19993 32212
rect 19392 32172 19398 32184
rect 19981 32181 19993 32184
rect 20027 32181 20039 32215
rect 20364 32212 20392 32252
rect 22066 32212 22094 32388
rect 22186 32308 22192 32360
rect 22244 32308 22250 32360
rect 22370 32308 22376 32360
rect 22428 32308 22434 32360
rect 22480 32348 22508 32388
rect 23474 32376 23480 32428
rect 23532 32376 23538 32428
rect 24210 32376 24216 32428
rect 24268 32416 24274 32428
rect 24670 32416 24676 32428
rect 24268 32388 24676 32416
rect 24268 32376 24274 32388
rect 24670 32376 24676 32388
rect 24728 32376 24734 32428
rect 25130 32348 25136 32360
rect 22480 32320 25136 32348
rect 25130 32308 25136 32320
rect 25188 32308 25194 32360
rect 25222 32308 25228 32360
rect 25280 32348 25286 32360
rect 25590 32348 25596 32360
rect 25280 32320 25596 32348
rect 25280 32308 25286 32320
rect 25590 32308 25596 32320
rect 25648 32308 25654 32360
rect 22204 32280 22232 32308
rect 24026 32280 24032 32292
rect 22204 32252 24032 32280
rect 24026 32240 24032 32252
rect 24084 32240 24090 32292
rect 20364 32184 22094 32212
rect 19981 32175 20039 32181
rect 22830 32172 22836 32224
rect 22888 32172 22894 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 6641 32011 6699 32017
rect 6641 31977 6653 32011
rect 6687 32008 6699 32011
rect 6914 32008 6920 32020
rect 6687 31980 6920 32008
rect 6687 31977 6699 31980
rect 6641 31971 6699 31977
rect 6914 31968 6920 31980
rect 6972 31968 6978 32020
rect 8757 32011 8815 32017
rect 8757 32008 8769 32011
rect 7024 31980 8769 32008
rect 7024 31790 7052 31980
rect 8757 31977 8769 31980
rect 8803 32008 8815 32011
rect 9674 32008 9680 32020
rect 8803 31980 9680 32008
rect 8803 31977 8815 31980
rect 8757 31971 8815 31977
rect 9674 31968 9680 31980
rect 9732 31968 9738 32020
rect 11146 31968 11152 32020
rect 11204 32008 11210 32020
rect 11609 32011 11667 32017
rect 11609 32008 11621 32011
rect 11204 31980 11621 32008
rect 11204 31968 11210 31980
rect 11609 31977 11621 31980
rect 11655 31977 11667 32011
rect 11609 31971 11667 31977
rect 11698 31968 11704 32020
rect 11756 32008 11762 32020
rect 11756 31980 12434 32008
rect 11756 31968 11762 31980
rect 12406 31940 12434 31980
rect 12618 31968 12624 32020
rect 12676 32008 12682 32020
rect 14277 32011 14335 32017
rect 14277 32008 14289 32011
rect 12676 31980 14289 32008
rect 12676 31968 12682 31980
rect 14277 31977 14289 31980
rect 14323 31977 14335 32011
rect 14277 31971 14335 31977
rect 15473 32011 15531 32017
rect 15473 31977 15485 32011
rect 15519 32008 15531 32011
rect 15654 32008 15660 32020
rect 15519 31980 15660 32008
rect 15519 31977 15531 31980
rect 15473 31971 15531 31977
rect 15654 31968 15660 31980
rect 15712 31968 15718 32020
rect 18322 32008 18328 32020
rect 15764 31980 18328 32008
rect 13817 31943 13875 31949
rect 13817 31940 13829 31943
rect 11440 31912 12296 31940
rect 12406 31912 13829 31940
rect 11440 31884 11468 31912
rect 8018 31832 8024 31884
rect 8076 31872 8082 31884
rect 8389 31875 8447 31881
rect 8389 31872 8401 31875
rect 8076 31844 8401 31872
rect 8076 31832 8082 31844
rect 8389 31841 8401 31844
rect 8435 31841 8447 31875
rect 8846 31872 8852 31884
rect 8389 31835 8447 31841
rect 8496 31844 8852 31872
rect 8496 31804 8524 31844
rect 8846 31832 8852 31844
rect 8904 31832 8910 31884
rect 9861 31875 9919 31881
rect 9861 31841 9873 31875
rect 9907 31872 9919 31875
rect 10226 31872 10232 31884
rect 9907 31844 10232 31872
rect 9907 31841 9919 31844
rect 9861 31835 9919 31841
rect 10226 31832 10232 31844
rect 10284 31872 10290 31884
rect 11422 31872 11428 31884
rect 10284 31844 11428 31872
rect 10284 31832 10290 31844
rect 11422 31832 11428 31844
rect 11480 31832 11486 31884
rect 11698 31832 11704 31884
rect 11756 31872 11762 31884
rect 12066 31872 12072 31884
rect 11756 31844 12072 31872
rect 11756 31832 11762 31844
rect 12066 31832 12072 31844
rect 12124 31832 12130 31884
rect 12268 31872 12296 31912
rect 13817 31909 13829 31912
rect 13863 31940 13875 31943
rect 13863 31912 14872 31940
rect 13863 31909 13875 31912
rect 13817 31903 13875 31909
rect 12342 31872 12348 31884
rect 12268 31844 12348 31872
rect 12342 31832 12348 31844
rect 12400 31832 12406 31884
rect 12802 31832 12808 31884
rect 12860 31832 12866 31884
rect 14844 31881 14872 31912
rect 14829 31875 14887 31881
rect 14829 31841 14841 31875
rect 14875 31841 14887 31875
rect 14829 31835 14887 31841
rect 8404 31776 8524 31804
rect 8113 31739 8171 31745
rect 8113 31705 8125 31739
rect 8159 31736 8171 31739
rect 8404 31736 8432 31776
rect 9582 31764 9588 31816
rect 9640 31804 9646 31816
rect 11885 31807 11943 31813
rect 11885 31804 11897 31807
rect 9640 31776 9904 31804
rect 11270 31776 11897 31804
rect 9640 31764 9646 31776
rect 8159 31708 8432 31736
rect 9876 31736 9904 31776
rect 11885 31773 11897 31776
rect 11931 31773 11943 31807
rect 11885 31767 11943 31773
rect 13354 31764 13360 31816
rect 13412 31804 13418 31816
rect 13633 31807 13691 31813
rect 13633 31804 13645 31807
rect 13412 31776 13645 31804
rect 13412 31764 13418 31776
rect 13633 31773 13645 31776
rect 13679 31773 13691 31807
rect 13633 31767 13691 31773
rect 14737 31807 14795 31813
rect 14737 31773 14749 31807
rect 14783 31804 14795 31807
rect 15764 31804 15792 31980
rect 18322 31968 18328 31980
rect 18380 31968 18386 32020
rect 19429 32011 19487 32017
rect 19429 31977 19441 32011
rect 19475 32008 19487 32011
rect 19610 32008 19616 32020
rect 19475 31980 19616 32008
rect 19475 31977 19487 31980
rect 19429 31971 19487 31977
rect 19610 31968 19616 31980
rect 19668 31968 19674 32020
rect 19794 31968 19800 32020
rect 19852 31968 19858 32020
rect 20622 31968 20628 32020
rect 20680 31968 20686 32020
rect 21637 32011 21695 32017
rect 21637 31977 21649 32011
rect 21683 32008 21695 32011
rect 22370 32008 22376 32020
rect 21683 31980 22376 32008
rect 21683 31977 21695 31980
rect 21637 31971 21695 31977
rect 22370 31968 22376 31980
rect 22428 31968 22434 32020
rect 22544 32011 22602 32017
rect 22544 31977 22556 32011
rect 22590 32008 22602 32011
rect 22646 32008 22652 32020
rect 22590 31980 22652 32008
rect 22590 31977 22602 31980
rect 22544 31971 22602 31977
rect 22646 31968 22652 31980
rect 22704 31968 22710 32020
rect 24026 31968 24032 32020
rect 24084 31968 24090 32020
rect 17402 31900 17408 31952
rect 17460 31940 17466 31952
rect 18414 31940 18420 31952
rect 17460 31912 18420 31940
rect 17460 31900 17466 31912
rect 18414 31900 18420 31912
rect 18472 31900 18478 31952
rect 19518 31900 19524 31952
rect 19576 31940 19582 31952
rect 20530 31940 20536 31952
rect 19576 31912 20536 31940
rect 19576 31900 19582 31912
rect 20530 31900 20536 31912
rect 20588 31900 20594 31952
rect 21910 31940 21916 31952
rect 21192 31912 21916 31940
rect 21192 31884 21220 31912
rect 21910 31900 21916 31912
rect 21968 31900 21974 31952
rect 16945 31875 17003 31881
rect 16945 31841 16957 31875
rect 16991 31872 17003 31875
rect 18325 31875 18383 31881
rect 18325 31872 18337 31875
rect 16991 31844 18337 31872
rect 16991 31841 17003 31844
rect 16945 31835 17003 31841
rect 18325 31841 18337 31844
rect 18371 31841 18383 31875
rect 18325 31835 18383 31841
rect 19426 31832 19432 31884
rect 19484 31872 19490 31884
rect 19613 31875 19671 31881
rect 19613 31872 19625 31875
rect 19484 31844 19625 31872
rect 19484 31832 19490 31844
rect 19613 31841 19625 31844
rect 19659 31841 19671 31875
rect 19613 31835 19671 31841
rect 21082 31832 21088 31884
rect 21140 31832 21146 31884
rect 21174 31832 21180 31884
rect 21232 31832 21238 31884
rect 22281 31875 22339 31881
rect 22281 31841 22293 31875
rect 22327 31872 22339 31875
rect 23290 31872 23296 31884
rect 22327 31844 23296 31872
rect 22327 31841 22339 31844
rect 22281 31835 22339 31841
rect 23290 31832 23296 31844
rect 23348 31832 23354 31884
rect 14783 31776 15792 31804
rect 17221 31807 17279 31813
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 17221 31773 17233 31807
rect 17267 31773 17279 31807
rect 17221 31767 17279 31773
rect 10137 31739 10195 31745
rect 10137 31736 10149 31739
rect 9876 31708 10149 31736
rect 8159 31705 8171 31708
rect 8113 31699 8171 31705
rect 10137 31705 10149 31708
rect 10183 31705 10195 31739
rect 10137 31699 10195 31705
rect 10686 31696 10692 31748
rect 10744 31696 10750 31748
rect 9122 31628 9128 31680
rect 9180 31628 9186 31680
rect 13648 31668 13676 31767
rect 13722 31696 13728 31748
rect 13780 31736 13786 31748
rect 15654 31736 15660 31748
rect 13780 31708 15660 31736
rect 13780 31696 13786 31708
rect 15654 31696 15660 31708
rect 15712 31696 15718 31748
rect 16514 31708 16620 31736
rect 16592 31680 16620 31708
rect 16666 31696 16672 31748
rect 16724 31736 16730 31748
rect 17236 31736 17264 31767
rect 17678 31764 17684 31816
rect 17736 31764 17742 31816
rect 24044 31804 24072 31968
rect 24581 31807 24639 31813
rect 24581 31804 24593 31807
rect 24044 31776 24593 31804
rect 24581 31773 24593 31776
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 18874 31736 18880 31748
rect 16724 31708 18880 31736
rect 16724 31696 16730 31708
rect 18874 31696 18880 31708
rect 18932 31736 18938 31748
rect 19242 31736 19248 31748
rect 18932 31708 19248 31736
rect 18932 31696 18938 31708
rect 19242 31696 19248 31708
rect 19300 31696 19306 31748
rect 24486 31736 24492 31748
rect 23782 31708 24492 31736
rect 24486 31696 24492 31708
rect 24544 31696 24550 31748
rect 13998 31668 14004 31680
rect 13648 31640 14004 31668
rect 13998 31628 14004 31640
rect 14056 31668 14062 31680
rect 14642 31668 14648 31680
rect 14056 31640 14648 31668
rect 14056 31628 14062 31640
rect 14642 31628 14648 31640
rect 14700 31628 14706 31680
rect 15102 31628 15108 31680
rect 15160 31668 15166 31680
rect 15930 31668 15936 31680
rect 15160 31640 15936 31668
rect 15160 31628 15166 31640
rect 15930 31628 15936 31640
rect 15988 31628 15994 31680
rect 16574 31628 16580 31680
rect 16632 31668 16638 31680
rect 17494 31668 17500 31680
rect 16632 31640 17500 31668
rect 16632 31628 16638 31640
rect 17494 31628 17500 31640
rect 17552 31628 17558 31680
rect 17770 31628 17776 31680
rect 17828 31668 17834 31680
rect 20346 31668 20352 31680
rect 17828 31640 20352 31668
rect 17828 31628 17834 31640
rect 20346 31628 20352 31640
rect 20404 31628 20410 31680
rect 21269 31671 21327 31677
rect 21269 31637 21281 31671
rect 21315 31668 21327 31671
rect 21358 31668 21364 31680
rect 21315 31640 21364 31668
rect 21315 31637 21327 31640
rect 21269 31631 21327 31637
rect 21358 31628 21364 31640
rect 21416 31668 21422 31680
rect 21634 31668 21640 31680
rect 21416 31640 21640 31668
rect 21416 31628 21422 31640
rect 21634 31628 21640 31640
rect 21692 31628 21698 31680
rect 22094 31628 22100 31680
rect 22152 31668 22158 31680
rect 23842 31668 23848 31680
rect 22152 31640 23848 31668
rect 22152 31628 22158 31640
rect 23842 31628 23848 31640
rect 23900 31628 23906 31680
rect 24946 31628 24952 31680
rect 25004 31668 25010 31680
rect 25225 31671 25283 31677
rect 25225 31668 25237 31671
rect 25004 31640 25237 31668
rect 25004 31628 25010 31640
rect 25225 31637 25237 31640
rect 25271 31637 25283 31671
rect 25225 31631 25283 31637
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 7837 31467 7895 31473
rect 7837 31433 7849 31467
rect 7883 31464 7895 31467
rect 9122 31464 9128 31476
rect 7883 31436 9128 31464
rect 7883 31433 7895 31436
rect 7837 31427 7895 31433
rect 9122 31424 9128 31436
rect 9180 31424 9186 31476
rect 15654 31424 15660 31476
rect 15712 31464 15718 31476
rect 15712 31436 16252 31464
rect 15712 31424 15718 31436
rect 13906 31356 13912 31408
rect 13964 31356 13970 31408
rect 16022 31356 16028 31408
rect 16080 31356 16086 31408
rect 16224 31396 16252 31436
rect 16298 31424 16304 31476
rect 16356 31424 16362 31476
rect 16942 31424 16948 31476
rect 17000 31464 17006 31476
rect 18325 31467 18383 31473
rect 17000 31436 17540 31464
rect 17000 31424 17006 31436
rect 17512 31396 17540 31436
rect 18325 31433 18337 31467
rect 18371 31464 18383 31467
rect 18598 31464 18604 31476
rect 18371 31436 18604 31464
rect 18371 31433 18383 31436
rect 18325 31427 18383 31433
rect 18598 31424 18604 31436
rect 18656 31424 18662 31476
rect 18690 31424 18696 31476
rect 18748 31424 18754 31476
rect 19889 31467 19947 31473
rect 19889 31433 19901 31467
rect 19935 31464 19947 31467
rect 20714 31464 20720 31476
rect 19935 31436 20720 31464
rect 19935 31433 19947 31436
rect 19889 31427 19947 31433
rect 20714 31424 20720 31436
rect 20772 31424 20778 31476
rect 20990 31424 20996 31476
rect 21048 31464 21054 31476
rect 21085 31467 21143 31473
rect 21085 31464 21097 31467
rect 21048 31436 21097 31464
rect 21048 31424 21054 31436
rect 21085 31433 21097 31436
rect 21131 31433 21143 31467
rect 21085 31427 21143 31433
rect 21174 31424 21180 31476
rect 21232 31424 21238 31476
rect 23290 31424 23296 31476
rect 23348 31464 23354 31476
rect 23348 31436 25268 31464
rect 23348 31424 23354 31436
rect 18708 31396 18736 31424
rect 16224 31368 17448 31396
rect 17512 31368 18736 31396
rect 19981 31399 20039 31405
rect 3694 31288 3700 31340
rect 3752 31328 3758 31340
rect 3789 31331 3847 31337
rect 3789 31328 3801 31331
rect 3752 31300 3801 31328
rect 3752 31288 3758 31300
rect 3789 31297 3801 31300
rect 3835 31297 3847 31331
rect 3789 31291 3847 31297
rect 10505 31331 10563 31337
rect 10505 31297 10517 31331
rect 10551 31328 10563 31331
rect 11330 31328 11336 31340
rect 10551 31300 11336 31328
rect 10551 31297 10563 31300
rect 10505 31291 10563 31297
rect 11330 31288 11336 31300
rect 11388 31288 11394 31340
rect 12342 31288 12348 31340
rect 12400 31328 12406 31340
rect 12621 31331 12679 31337
rect 12621 31328 12633 31331
rect 12400 31300 12633 31328
rect 12400 31288 12406 31300
rect 12621 31297 12633 31300
rect 12667 31297 12679 31331
rect 12621 31291 12679 31297
rect 15197 31331 15255 31337
rect 15197 31297 15209 31331
rect 15243 31297 15255 31331
rect 15197 31291 15255 31297
rect 15289 31331 15347 31337
rect 15289 31297 15301 31331
rect 15335 31328 15347 31331
rect 16040 31328 16068 31356
rect 15335 31300 16068 31328
rect 15335 31297 15347 31300
rect 15289 31291 15347 31297
rect 3970 31220 3976 31272
rect 4028 31220 4034 31272
rect 4890 31220 4896 31272
rect 4948 31220 4954 31272
rect 7006 31220 7012 31272
rect 7064 31260 7070 31272
rect 7193 31263 7251 31269
rect 7193 31260 7205 31263
rect 7064 31232 7205 31260
rect 7064 31220 7070 31232
rect 7193 31229 7205 31232
rect 7239 31260 7251 31263
rect 7650 31260 7656 31272
rect 7239 31232 7656 31260
rect 7239 31229 7251 31232
rect 7193 31223 7251 31229
rect 7650 31220 7656 31232
rect 7708 31220 7714 31272
rect 7745 31263 7803 31269
rect 7745 31229 7757 31263
rect 7791 31260 7803 31263
rect 8294 31260 8300 31272
rect 7791 31232 8300 31260
rect 7791 31229 7803 31232
rect 7745 31223 7803 31229
rect 5258 31152 5264 31204
rect 5316 31192 5322 31204
rect 6917 31195 6975 31201
rect 6917 31192 6929 31195
rect 5316 31164 6929 31192
rect 5316 31152 5322 31164
rect 6917 31161 6929 31164
rect 6963 31192 6975 31195
rect 7760 31192 7788 31223
rect 8294 31220 8300 31232
rect 8352 31220 8358 31272
rect 12897 31263 12955 31269
rect 12897 31229 12909 31263
rect 12943 31260 12955 31263
rect 14918 31260 14924 31272
rect 12943 31232 14924 31260
rect 12943 31229 12955 31232
rect 12897 31223 12955 31229
rect 14918 31220 14924 31232
rect 14976 31220 14982 31272
rect 6963 31164 7788 31192
rect 6963 31161 6975 31164
rect 6917 31155 6975 31161
rect 7834 31152 7840 31204
rect 7892 31192 7898 31204
rect 8205 31195 8263 31201
rect 8205 31192 8217 31195
rect 7892 31164 8217 31192
rect 7892 31152 7898 31164
rect 8205 31161 8217 31164
rect 8251 31161 8263 31195
rect 14829 31195 14887 31201
rect 14829 31192 14841 31195
rect 8205 31155 8263 31161
rect 13924 31164 14841 31192
rect 11149 31127 11207 31133
rect 11149 31093 11161 31127
rect 11195 31124 11207 31127
rect 11238 31124 11244 31136
rect 11195 31096 11244 31124
rect 11195 31093 11207 31096
rect 11149 31087 11207 31093
rect 11238 31084 11244 31096
rect 11296 31084 11302 31136
rect 12066 31084 12072 31136
rect 12124 31124 12130 31136
rect 13924 31124 13952 31164
rect 14829 31161 14841 31164
rect 14875 31161 14887 31195
rect 15212 31192 15240 31291
rect 17218 31288 17224 31340
rect 17276 31288 17282 31340
rect 15470 31220 15476 31272
rect 15528 31220 15534 31272
rect 17420 31269 17448 31368
rect 19981 31365 19993 31399
rect 20027 31396 20039 31399
rect 20898 31396 20904 31408
rect 20027 31368 20904 31396
rect 20027 31365 20039 31368
rect 19981 31359 20039 31365
rect 20898 31356 20904 31368
rect 20956 31356 20962 31408
rect 22281 31399 22339 31405
rect 22281 31365 22293 31399
rect 22327 31396 22339 31399
rect 23109 31399 23167 31405
rect 23109 31396 23121 31399
rect 22327 31368 23121 31396
rect 22327 31365 22339 31368
rect 22281 31359 22339 31365
rect 23109 31365 23121 31368
rect 23155 31396 23167 31399
rect 23382 31396 23388 31408
rect 23155 31368 23388 31396
rect 23155 31365 23167 31368
rect 23109 31359 23167 31365
rect 23382 31356 23388 31368
rect 23440 31356 23446 31408
rect 24486 31356 24492 31408
rect 24544 31356 24550 31408
rect 24946 31356 24952 31408
rect 25004 31356 25010 31408
rect 18690 31288 18696 31340
rect 18748 31288 18754 31340
rect 25240 31337 25268 31436
rect 18785 31331 18843 31337
rect 18785 31297 18797 31331
rect 18831 31328 18843 31331
rect 22373 31331 22431 31337
rect 22373 31328 22385 31331
rect 18831 31300 22385 31328
rect 18831 31297 18843 31300
rect 18785 31291 18843 31297
rect 22373 31297 22385 31300
rect 22419 31328 22431 31331
rect 25225 31331 25283 31337
rect 22419 31300 23612 31328
rect 22419 31297 22431 31300
rect 22373 31291 22431 31297
rect 17313 31263 17371 31269
rect 17313 31229 17325 31263
rect 17359 31229 17371 31263
rect 17313 31223 17371 31229
rect 17405 31263 17463 31269
rect 17405 31229 17417 31263
rect 17451 31229 17463 31263
rect 17405 31223 17463 31229
rect 18877 31263 18935 31269
rect 18877 31229 18889 31263
rect 18923 31229 18935 31263
rect 18877 31223 18935 31229
rect 16298 31192 16304 31204
rect 15212 31164 16304 31192
rect 14829 31155 14887 31161
rect 16298 31152 16304 31164
rect 16356 31152 16362 31204
rect 16666 31152 16672 31204
rect 16724 31192 16730 31204
rect 16853 31195 16911 31201
rect 16853 31192 16865 31195
rect 16724 31164 16865 31192
rect 16724 31152 16730 31164
rect 16853 31161 16865 31164
rect 16899 31161 16911 31195
rect 17328 31192 17356 31223
rect 17770 31192 17776 31204
rect 17328 31164 17776 31192
rect 16853 31155 16911 31161
rect 17770 31152 17776 31164
rect 17828 31152 17834 31204
rect 12124 31096 13952 31124
rect 12124 31084 12130 31096
rect 14090 31084 14096 31136
rect 14148 31124 14154 31136
rect 14369 31127 14427 31133
rect 14369 31124 14381 31127
rect 14148 31096 14381 31124
rect 14148 31084 14154 31096
rect 14369 31093 14381 31096
rect 14415 31124 14427 31127
rect 14458 31124 14464 31136
rect 14415 31096 14464 31124
rect 14415 31093 14427 31096
rect 14369 31087 14427 31093
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 14642 31084 14648 31136
rect 14700 31124 14706 31136
rect 15841 31127 15899 31133
rect 15841 31124 15853 31127
rect 14700 31096 15853 31124
rect 14700 31084 14706 31096
rect 15841 31093 15853 31096
rect 15887 31093 15899 31127
rect 15841 31087 15899 31093
rect 15930 31084 15936 31136
rect 15988 31124 15994 31136
rect 18892 31124 18920 31223
rect 18966 31220 18972 31272
rect 19024 31260 19030 31272
rect 20073 31263 20131 31269
rect 20073 31260 20085 31263
rect 19024 31232 20085 31260
rect 19024 31220 19030 31232
rect 20073 31229 20085 31232
rect 20119 31229 20131 31263
rect 20073 31223 20131 31229
rect 21266 31220 21272 31272
rect 21324 31220 21330 31272
rect 22094 31220 22100 31272
rect 22152 31220 22158 31272
rect 23474 31220 23480 31272
rect 23532 31220 23538 31272
rect 23584 31260 23612 31300
rect 25225 31297 25237 31331
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 25498 31260 25504 31272
rect 23584 31232 25504 31260
rect 25498 31220 25504 31232
rect 25556 31220 25562 31272
rect 15988 31096 18920 31124
rect 19521 31127 19579 31133
rect 15988 31084 15994 31096
rect 19521 31093 19533 31127
rect 19567 31124 19579 31127
rect 19610 31124 19616 31136
rect 19567 31096 19616 31124
rect 19567 31093 19579 31096
rect 19521 31087 19579 31093
rect 19610 31084 19616 31096
rect 19668 31084 19674 31136
rect 20714 31084 20720 31136
rect 20772 31084 20778 31136
rect 22646 31084 22652 31136
rect 22704 31124 22710 31136
rect 22741 31127 22799 31133
rect 22741 31124 22753 31127
rect 22704 31096 22753 31124
rect 22704 31084 22710 31096
rect 22741 31093 22753 31096
rect 22787 31093 22799 31127
rect 22741 31087 22799 31093
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 7650 30880 7656 30932
rect 7708 30880 7714 30932
rect 8297 30923 8355 30929
rect 8297 30889 8309 30923
rect 8343 30920 8355 30923
rect 8478 30920 8484 30932
rect 8343 30892 8484 30920
rect 8343 30889 8355 30892
rect 8297 30883 8355 30889
rect 8478 30880 8484 30892
rect 8536 30880 8542 30932
rect 8588 30892 11376 30920
rect 7668 30852 7696 30880
rect 8588 30852 8616 30892
rect 7668 30824 8616 30852
rect 11348 30852 11376 30892
rect 12158 30880 12164 30932
rect 12216 30920 12222 30932
rect 12621 30923 12679 30929
rect 12621 30920 12633 30923
rect 12216 30892 12633 30920
rect 12216 30880 12222 30892
rect 12621 30889 12633 30892
rect 12667 30889 12679 30923
rect 12621 30883 12679 30889
rect 14274 30880 14280 30932
rect 14332 30920 14338 30932
rect 16666 30920 16672 30932
rect 14332 30892 16672 30920
rect 14332 30880 14338 30892
rect 16666 30880 16672 30892
rect 16724 30880 16730 30932
rect 17126 30880 17132 30932
rect 17184 30880 17190 30932
rect 17862 30880 17868 30932
rect 17920 30920 17926 30932
rect 17920 30892 19012 30920
rect 17920 30880 17926 30892
rect 11348 30824 13216 30852
rect 6914 30744 6920 30796
rect 6972 30784 6978 30796
rect 7653 30787 7711 30793
rect 7653 30784 7665 30787
rect 6972 30756 7665 30784
rect 6972 30744 6978 30756
rect 7653 30753 7665 30756
rect 7699 30753 7711 30787
rect 7653 30747 7711 30753
rect 11146 30744 11152 30796
rect 11204 30744 11210 30796
rect 11422 30744 11428 30796
rect 11480 30744 11486 30796
rect 13188 30793 13216 30824
rect 15838 30812 15844 30864
rect 15896 30812 15902 30864
rect 17494 30812 17500 30864
rect 17552 30812 17558 30864
rect 13173 30787 13231 30793
rect 13173 30753 13185 30787
rect 13219 30784 13231 30787
rect 13633 30787 13691 30793
rect 13633 30784 13645 30787
rect 13219 30756 13645 30784
rect 13219 30753 13231 30756
rect 13173 30747 13231 30753
rect 13633 30753 13645 30756
rect 13679 30753 13691 30787
rect 13633 30747 13691 30753
rect 13906 30744 13912 30796
rect 13964 30784 13970 30796
rect 14642 30784 14648 30796
rect 13964 30756 14648 30784
rect 13964 30744 13970 30756
rect 14642 30744 14648 30756
rect 14700 30744 14706 30796
rect 16022 30744 16028 30796
rect 16080 30784 16086 30796
rect 16485 30787 16543 30793
rect 16485 30784 16497 30787
rect 16080 30756 16497 30784
rect 16080 30744 16086 30756
rect 16485 30753 16497 30756
rect 16531 30784 16543 30787
rect 16942 30784 16948 30796
rect 16531 30756 16948 30784
rect 16531 30753 16543 30756
rect 16485 30747 16543 30753
rect 16942 30744 16948 30756
rect 17000 30744 17006 30796
rect 17512 30784 17540 30812
rect 17862 30784 17868 30796
rect 17512 30756 17868 30784
rect 17862 30744 17868 30756
rect 17920 30744 17926 30796
rect 7742 30676 7748 30728
rect 7800 30716 7806 30728
rect 7929 30719 7987 30725
rect 7929 30716 7941 30719
rect 7800 30688 7941 30716
rect 7800 30676 7806 30688
rect 7929 30685 7941 30688
rect 7975 30685 7987 30719
rect 7929 30679 7987 30685
rect 14369 30719 14427 30725
rect 14369 30685 14381 30719
rect 14415 30716 14427 30719
rect 15194 30716 15200 30728
rect 14415 30688 15200 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 15194 30676 15200 30688
rect 15252 30716 15258 30728
rect 15252 30688 15424 30716
rect 15252 30676 15258 30688
rect 10686 30608 10692 30660
rect 10744 30648 10750 30660
rect 10870 30648 10876 30660
rect 10744 30620 10876 30648
rect 10744 30608 10750 30620
rect 10870 30608 10876 30620
rect 10928 30608 10934 30660
rect 15396 30657 15424 30688
rect 18874 30676 18880 30728
rect 18932 30676 18938 30728
rect 18984 30716 19012 30892
rect 21174 30880 21180 30932
rect 21232 30920 21238 30932
rect 21545 30923 21603 30929
rect 21545 30920 21557 30923
rect 21232 30892 21557 30920
rect 21232 30880 21238 30892
rect 21545 30889 21557 30892
rect 21591 30889 21603 30923
rect 21545 30883 21603 30889
rect 20257 30855 20315 30861
rect 20257 30821 20269 30855
rect 20303 30852 20315 30855
rect 22922 30852 22928 30864
rect 20303 30824 22928 30852
rect 20303 30821 20315 30824
rect 20257 30815 20315 30821
rect 22922 30812 22928 30824
rect 22980 30812 22986 30864
rect 19705 30787 19763 30793
rect 19705 30753 19717 30787
rect 19751 30784 19763 30787
rect 20070 30784 20076 30796
rect 19751 30756 20076 30784
rect 19751 30753 19763 30756
rect 19705 30747 19763 30753
rect 20070 30744 20076 30756
rect 20128 30744 20134 30796
rect 23109 30787 23167 30793
rect 23109 30753 23121 30787
rect 23155 30784 23167 30787
rect 23474 30784 23480 30796
rect 23155 30756 23480 30784
rect 23155 30753 23167 30756
rect 23109 30747 23167 30753
rect 23474 30744 23480 30756
rect 23532 30744 23538 30796
rect 20717 30719 20775 30725
rect 20717 30716 20729 30719
rect 18984 30688 20729 30716
rect 20717 30685 20729 30688
rect 20763 30685 20775 30719
rect 20717 30679 20775 30685
rect 22830 30676 22836 30728
rect 22888 30716 22894 30728
rect 23201 30719 23259 30725
rect 23201 30716 23213 30719
rect 22888 30688 23213 30716
rect 22888 30676 22894 30688
rect 23201 30685 23213 30688
rect 23247 30685 23259 30719
rect 23201 30679 23259 30685
rect 24578 30676 24584 30728
rect 24636 30676 24642 30728
rect 15381 30651 15439 30657
rect 15381 30617 15393 30651
rect 15427 30648 15439 30651
rect 15427 30620 16804 30648
rect 15427 30617 15439 30620
rect 15381 30611 15439 30617
rect 7837 30583 7895 30589
rect 7837 30549 7849 30583
rect 7883 30580 7895 30583
rect 8386 30580 8392 30592
rect 7883 30552 8392 30580
rect 7883 30549 7895 30552
rect 7837 30543 7895 30549
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 9677 30583 9735 30589
rect 9677 30549 9689 30583
rect 9723 30580 9735 30583
rect 11330 30580 11336 30592
rect 9723 30552 11336 30580
rect 9723 30549 9735 30552
rect 9677 30543 9735 30549
rect 11330 30540 11336 30552
rect 11388 30540 11394 30592
rect 11882 30540 11888 30592
rect 11940 30540 11946 30592
rect 12434 30540 12440 30592
rect 12492 30580 12498 30592
rect 12989 30583 13047 30589
rect 12989 30580 13001 30583
rect 12492 30552 13001 30580
rect 12492 30540 12498 30552
rect 12989 30549 13001 30552
rect 13035 30549 13047 30583
rect 12989 30543 13047 30549
rect 13081 30583 13139 30589
rect 13081 30549 13093 30583
rect 13127 30580 13139 30583
rect 13722 30580 13728 30592
rect 13127 30552 13728 30580
rect 13127 30549 13139 30552
rect 13081 30543 13139 30549
rect 13722 30540 13728 30552
rect 13780 30540 13786 30592
rect 15102 30540 15108 30592
rect 15160 30580 15166 30592
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 15160 30552 15485 30580
rect 15160 30540 15166 30552
rect 15473 30549 15485 30552
rect 15519 30580 15531 30583
rect 16209 30583 16267 30589
rect 16209 30580 16221 30583
rect 15519 30552 16221 30580
rect 15519 30549 15531 30552
rect 15473 30543 15531 30549
rect 16209 30549 16221 30552
rect 16255 30549 16267 30583
rect 16209 30543 16267 30549
rect 16298 30540 16304 30592
rect 16356 30540 16362 30592
rect 16776 30580 16804 30620
rect 17862 30608 17868 30660
rect 17920 30608 17926 30660
rect 18601 30651 18659 30657
rect 18601 30617 18613 30651
rect 18647 30648 18659 30651
rect 19702 30648 19708 30660
rect 18647 30620 19708 30648
rect 18647 30617 18659 30620
rect 18601 30611 18659 30617
rect 19702 30608 19708 30620
rect 19760 30608 19766 30660
rect 19794 30608 19800 30660
rect 19852 30648 19858 30660
rect 21177 30651 21235 30657
rect 21177 30648 21189 30651
rect 19852 30620 21189 30648
rect 19852 30608 19858 30620
rect 21177 30617 21189 30620
rect 21223 30617 21235 30651
rect 21177 30611 21235 30617
rect 18322 30580 18328 30592
rect 16776 30552 18328 30580
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 19518 30540 19524 30592
rect 19576 30580 19582 30592
rect 19889 30583 19947 30589
rect 19889 30580 19901 30583
rect 19576 30552 19901 30580
rect 19576 30540 19582 30552
rect 19889 30549 19901 30552
rect 19935 30549 19947 30583
rect 19889 30543 19947 30549
rect 20901 30583 20959 30589
rect 20901 30549 20913 30583
rect 20947 30580 20959 30583
rect 21082 30580 21088 30592
rect 20947 30552 21088 30580
rect 20947 30549 20959 30552
rect 20901 30543 20959 30549
rect 21082 30540 21088 30552
rect 21140 30540 21146 30592
rect 21358 30540 21364 30592
rect 21416 30580 21422 30592
rect 21913 30583 21971 30589
rect 21913 30580 21925 30583
rect 21416 30552 21925 30580
rect 21416 30540 21422 30552
rect 21913 30549 21925 30552
rect 21959 30549 21971 30583
rect 21913 30543 21971 30549
rect 23290 30540 23296 30592
rect 23348 30540 23354 30592
rect 23661 30583 23719 30589
rect 23661 30549 23673 30583
rect 23707 30580 23719 30583
rect 23934 30580 23940 30592
rect 23707 30552 23940 30580
rect 23707 30549 23719 30552
rect 23661 30543 23719 30549
rect 23934 30540 23940 30552
rect 23992 30540 23998 30592
rect 24765 30583 24823 30589
rect 24765 30549 24777 30583
rect 24811 30580 24823 30583
rect 24854 30580 24860 30592
rect 24811 30552 24860 30580
rect 24811 30549 24823 30552
rect 24765 30543 24823 30549
rect 24854 30540 24860 30552
rect 24912 30540 24918 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 9766 30336 9772 30388
rect 9824 30376 9830 30388
rect 15470 30376 15476 30388
rect 9824 30348 15476 30376
rect 9824 30336 9830 30348
rect 15470 30336 15476 30348
rect 15528 30336 15534 30388
rect 16298 30336 16304 30388
rect 16356 30376 16362 30388
rect 16761 30379 16819 30385
rect 16761 30376 16773 30379
rect 16356 30348 16773 30376
rect 16356 30336 16362 30348
rect 16761 30345 16773 30348
rect 16807 30376 16819 30379
rect 17402 30376 17408 30388
rect 16807 30348 17408 30376
rect 16807 30345 16819 30348
rect 16761 30339 16819 30345
rect 17402 30336 17408 30348
rect 17460 30336 17466 30388
rect 17770 30336 17776 30388
rect 17828 30336 17834 30388
rect 18322 30336 18328 30388
rect 18380 30376 18386 30388
rect 25222 30376 25228 30388
rect 18380 30348 25228 30376
rect 18380 30336 18386 30348
rect 25222 30336 25228 30348
rect 25280 30376 25286 30388
rect 25280 30348 25360 30376
rect 25280 30336 25286 30348
rect 4338 30268 4344 30320
rect 4396 30308 4402 30320
rect 8662 30308 8668 30320
rect 4396 30280 8668 30308
rect 4396 30268 4402 30280
rect 8662 30268 8668 30280
rect 8720 30308 8726 30320
rect 9585 30311 9643 30317
rect 9585 30308 9597 30311
rect 8720 30280 9597 30308
rect 8720 30268 8726 30280
rect 9585 30277 9597 30280
rect 9631 30277 9643 30311
rect 9585 30271 9643 30277
rect 10781 30311 10839 30317
rect 10781 30277 10793 30311
rect 10827 30308 10839 30311
rect 11882 30308 11888 30320
rect 10827 30280 11888 30308
rect 10827 30277 10839 30280
rect 10781 30271 10839 30277
rect 11882 30268 11888 30280
rect 11940 30268 11946 30320
rect 12710 30268 12716 30320
rect 12768 30308 12774 30320
rect 12897 30311 12955 30317
rect 12897 30308 12909 30311
rect 12768 30280 12909 30308
rect 12768 30268 12774 30280
rect 12897 30277 12909 30280
rect 12943 30277 12955 30311
rect 12897 30271 12955 30277
rect 14734 30268 14740 30320
rect 14792 30308 14798 30320
rect 17037 30311 17095 30317
rect 17037 30308 17049 30311
rect 14792 30280 17049 30308
rect 14792 30268 14798 30280
rect 8570 30200 8576 30252
rect 8628 30240 8634 30252
rect 8846 30240 8852 30252
rect 8628 30212 8852 30240
rect 8628 30200 8634 30212
rect 8846 30200 8852 30212
rect 8904 30240 8910 30252
rect 9493 30243 9551 30249
rect 9493 30240 9505 30243
rect 8904 30212 9505 30240
rect 8904 30200 8910 30212
rect 9493 30209 9505 30212
rect 9539 30209 9551 30243
rect 11054 30240 11060 30252
rect 9493 30203 9551 30209
rect 10612 30212 11060 30240
rect 10612 30181 10640 30212
rect 11054 30200 11060 30212
rect 11112 30200 11118 30252
rect 12989 30243 13047 30249
rect 12989 30240 13001 30243
rect 11164 30212 13001 30240
rect 9401 30175 9459 30181
rect 9401 30141 9413 30175
rect 9447 30141 9459 30175
rect 9401 30135 9459 30141
rect 10597 30175 10655 30181
rect 10597 30141 10609 30175
rect 10643 30141 10655 30175
rect 10597 30135 10655 30141
rect 10689 30175 10747 30181
rect 10689 30141 10701 30175
rect 10735 30141 10747 30175
rect 10689 30135 10747 30141
rect 9416 30104 9444 30135
rect 9582 30104 9588 30116
rect 9416 30076 9588 30104
rect 9582 30064 9588 30076
rect 9640 30064 9646 30116
rect 9950 30064 9956 30116
rect 10008 30064 10014 30116
rect 8662 29996 8668 30048
rect 8720 29996 8726 30048
rect 8846 29996 8852 30048
rect 8904 29996 8910 30048
rect 9858 29996 9864 30048
rect 9916 30036 9922 30048
rect 10704 30036 10732 30135
rect 11164 30113 11192 30212
rect 12989 30209 13001 30212
rect 13035 30209 13047 30243
rect 12989 30203 13047 30209
rect 11330 30132 11336 30184
rect 11388 30172 11394 30184
rect 12713 30175 12771 30181
rect 12713 30172 12725 30175
rect 11388 30144 12725 30172
rect 11388 30132 11394 30144
rect 12713 30141 12725 30144
rect 12759 30141 12771 30175
rect 12713 30135 12771 30141
rect 11149 30107 11207 30113
rect 11149 30073 11161 30107
rect 11195 30073 11207 30107
rect 11149 30067 11207 30073
rect 11609 30107 11667 30113
rect 11609 30073 11621 30107
rect 11655 30104 11667 30107
rect 11882 30104 11888 30116
rect 11655 30076 11888 30104
rect 11655 30073 11667 30076
rect 11609 30067 11667 30073
rect 11882 30064 11888 30076
rect 11940 30064 11946 30116
rect 16868 30104 16896 30280
rect 17037 30277 17049 30280
rect 17083 30277 17095 30311
rect 17037 30271 17095 30277
rect 17126 30268 17132 30320
rect 17184 30308 17190 30320
rect 17788 30308 17816 30336
rect 17184 30280 18736 30308
rect 17184 30268 17190 30280
rect 16942 30200 16948 30252
rect 17000 30240 17006 30252
rect 18708 30249 18736 30280
rect 19702 30268 19708 30320
rect 19760 30308 19766 30320
rect 19797 30311 19855 30317
rect 19797 30308 19809 30311
rect 19760 30280 19809 30308
rect 19760 30268 19766 30280
rect 19797 30277 19809 30280
rect 19843 30277 19855 30311
rect 24946 30308 24952 30320
rect 19797 30271 19855 30277
rect 23216 30280 24952 30308
rect 17681 30243 17739 30249
rect 17681 30240 17693 30243
rect 17000 30212 17693 30240
rect 17000 30200 17006 30212
rect 17681 30209 17693 30212
rect 17727 30209 17739 30243
rect 17681 30203 17739 30209
rect 17773 30243 17831 30249
rect 17773 30209 17785 30243
rect 17819 30209 17831 30243
rect 17773 30203 17831 30209
rect 18693 30243 18751 30249
rect 18693 30209 18705 30243
rect 18739 30209 18751 30243
rect 18693 30203 18751 30209
rect 17494 30132 17500 30184
rect 17552 30132 17558 30184
rect 17788 30172 17816 30203
rect 19886 30200 19892 30252
rect 19944 30240 19950 30252
rect 20438 30240 20444 30252
rect 19944 30212 20444 30240
rect 19944 30200 19950 30212
rect 20438 30200 20444 30212
rect 20496 30200 20502 30252
rect 23216 30249 23244 30280
rect 24946 30268 24952 30280
rect 25004 30268 25010 30320
rect 25332 30317 25360 30348
rect 25317 30311 25375 30317
rect 25317 30277 25329 30311
rect 25363 30308 25375 30311
rect 25406 30308 25412 30320
rect 25363 30280 25412 30308
rect 25363 30277 25375 30280
rect 25317 30271 25375 30277
rect 25406 30268 25412 30280
rect 25464 30268 25470 30320
rect 22741 30243 22799 30249
rect 22741 30209 22753 30243
rect 22787 30240 22799 30243
rect 23201 30243 23259 30249
rect 23201 30240 23213 30243
rect 22787 30212 23213 30240
rect 22787 30209 22799 30212
rect 22741 30203 22799 30209
rect 23201 30209 23213 30212
rect 23247 30209 23259 30243
rect 23201 30203 23259 30209
rect 23658 30200 23664 30252
rect 23716 30200 23722 30252
rect 24486 30200 24492 30252
rect 24544 30200 24550 30252
rect 17696 30144 17816 30172
rect 17126 30104 17132 30116
rect 16868 30076 17132 30104
rect 17126 30064 17132 30076
rect 17184 30104 17190 30116
rect 17696 30104 17724 30144
rect 19242 30132 19248 30184
rect 19300 30172 19306 30184
rect 19426 30172 19432 30184
rect 19300 30144 19432 30172
rect 19300 30132 19306 30144
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 20898 30132 20904 30184
rect 20956 30132 20962 30184
rect 17184 30076 17724 30104
rect 18141 30107 18199 30113
rect 17184 30064 17190 30076
rect 18141 30073 18153 30107
rect 18187 30104 18199 30107
rect 19794 30104 19800 30116
rect 18187 30076 19800 30104
rect 18187 30073 18199 30076
rect 18141 30067 18199 30073
rect 19794 30064 19800 30076
rect 19852 30064 19858 30116
rect 20254 30064 20260 30116
rect 20312 30104 20318 30116
rect 20530 30104 20536 30116
rect 20312 30076 20536 30104
rect 20312 30064 20318 30076
rect 20530 30064 20536 30076
rect 20588 30104 20594 30116
rect 23017 30107 23075 30113
rect 23017 30104 23029 30107
rect 20588 30076 23029 30104
rect 20588 30064 20594 30076
rect 23017 30073 23029 30076
rect 23063 30073 23075 30107
rect 23017 30067 23075 30073
rect 11790 30036 11796 30048
rect 9916 30008 11796 30036
rect 9916 29996 9922 30008
rect 11790 29996 11796 30008
rect 11848 29996 11854 30048
rect 12342 29996 12348 30048
rect 12400 29996 12406 30048
rect 13357 30039 13415 30045
rect 13357 30005 13369 30039
rect 13403 30036 13415 30039
rect 14366 30036 14372 30048
rect 13403 30008 14372 30036
rect 13403 30005 13415 30008
rect 13357 29999 13415 30005
rect 14366 29996 14372 30008
rect 14424 29996 14430 30048
rect 18414 29996 18420 30048
rect 18472 30036 18478 30048
rect 19337 30039 19395 30045
rect 19337 30036 19349 30039
rect 18472 30008 19349 30036
rect 18472 29996 18478 30008
rect 19337 30005 19349 30008
rect 19383 30005 19395 30039
rect 19337 29999 19395 30005
rect 19978 29996 19984 30048
rect 20036 30036 20042 30048
rect 20438 30036 20444 30048
rect 20036 30008 20444 30036
rect 20036 29996 20042 30008
rect 20438 29996 20444 30008
rect 20496 30036 20502 30048
rect 21910 30036 21916 30048
rect 20496 30008 21916 30036
rect 20496 29996 20502 30008
rect 21910 29996 21916 30008
rect 21968 29996 21974 30048
rect 23845 30039 23903 30045
rect 23845 30005 23857 30039
rect 23891 30036 23903 30039
rect 24026 30036 24032 30048
rect 23891 30008 24032 30036
rect 23891 30005 23903 30008
rect 23845 29999 23903 30005
rect 24026 29996 24032 30008
rect 24084 29996 24090 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 5074 29792 5080 29844
rect 5132 29832 5138 29844
rect 8021 29835 8079 29841
rect 8021 29832 8033 29835
rect 5132 29804 8033 29832
rect 5132 29792 5138 29804
rect 8021 29801 8033 29804
rect 8067 29832 8079 29835
rect 8570 29832 8576 29844
rect 8067 29804 8576 29832
rect 8067 29801 8079 29804
rect 8021 29795 8079 29801
rect 8570 29792 8576 29804
rect 8628 29792 8634 29844
rect 11882 29792 11888 29844
rect 11940 29832 11946 29844
rect 13906 29832 13912 29844
rect 11940 29804 13912 29832
rect 11940 29792 11946 29804
rect 13906 29792 13912 29804
rect 13964 29792 13970 29844
rect 15197 29835 15255 29841
rect 15197 29801 15209 29835
rect 15243 29832 15255 29835
rect 15286 29832 15292 29844
rect 15243 29804 15292 29832
rect 15243 29801 15255 29804
rect 15197 29795 15255 29801
rect 15286 29792 15292 29804
rect 15344 29792 15350 29844
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 16945 29835 17003 29841
rect 16945 29832 16957 29835
rect 16632 29804 16957 29832
rect 16632 29792 16638 29804
rect 16945 29801 16957 29804
rect 16991 29832 17003 29835
rect 17678 29832 17684 29844
rect 16991 29804 17684 29832
rect 16991 29801 17003 29804
rect 16945 29795 17003 29801
rect 17678 29792 17684 29804
rect 17736 29792 17742 29844
rect 18046 29792 18052 29844
rect 18104 29832 18110 29844
rect 21818 29832 21824 29844
rect 18104 29804 21824 29832
rect 18104 29792 18110 29804
rect 21818 29792 21824 29804
rect 21876 29792 21882 29844
rect 22005 29835 22063 29841
rect 22005 29801 22017 29835
rect 22051 29832 22063 29835
rect 23290 29832 23296 29844
rect 22051 29804 23296 29832
rect 22051 29801 22063 29804
rect 22005 29795 22063 29801
rect 23290 29792 23296 29804
rect 23348 29792 23354 29844
rect 25406 29792 25412 29844
rect 25464 29792 25470 29844
rect 4062 29656 4068 29708
rect 4120 29656 4126 29708
rect 11238 29656 11244 29708
rect 11296 29656 11302 29708
rect 11514 29656 11520 29708
rect 11572 29656 11578 29708
rect 3510 29520 3516 29572
rect 3568 29560 3574 29572
rect 4249 29563 4307 29569
rect 4249 29560 4261 29563
rect 3568 29532 4261 29560
rect 3568 29520 3574 29532
rect 4249 29529 4261 29532
rect 4295 29529 4307 29563
rect 4249 29523 4307 29529
rect 5905 29563 5963 29569
rect 5905 29529 5917 29563
rect 5951 29560 5963 29563
rect 6178 29560 6184 29572
rect 5951 29532 6184 29560
rect 5951 29529 5963 29532
rect 5905 29523 5963 29529
rect 6178 29520 6184 29532
rect 6236 29520 6242 29572
rect 11900 29560 11928 29792
rect 20901 29767 20959 29773
rect 20901 29764 20913 29767
rect 18984 29736 20913 29764
rect 17218 29656 17224 29708
rect 17276 29696 17282 29708
rect 18046 29696 18052 29708
rect 17276 29668 18052 29696
rect 17276 29656 17282 29668
rect 18046 29656 18052 29668
rect 18104 29656 18110 29708
rect 18414 29656 18420 29708
rect 18472 29656 18478 29708
rect 18693 29699 18751 29705
rect 18693 29665 18705 29699
rect 18739 29696 18751 29699
rect 18874 29696 18880 29708
rect 18739 29668 18880 29696
rect 18739 29665 18751 29668
rect 18693 29659 18751 29665
rect 18874 29656 18880 29668
rect 18932 29656 18938 29708
rect 18984 29628 19012 29736
rect 20901 29733 20913 29736
rect 20947 29733 20959 29767
rect 20901 29727 20959 29733
rect 19426 29656 19432 29708
rect 19484 29696 19490 29708
rect 19613 29699 19671 29705
rect 19613 29696 19625 29699
rect 19484 29668 19625 29696
rect 19484 29656 19490 29668
rect 19613 29665 19625 29668
rect 19659 29665 19671 29699
rect 19613 29659 19671 29665
rect 19794 29656 19800 29708
rect 19852 29656 19858 29708
rect 18708 29600 19012 29628
rect 19889 29631 19947 29637
rect 10810 29532 11928 29560
rect 16485 29563 16543 29569
rect 10888 29504 10916 29532
rect 16485 29529 16497 29563
rect 16531 29560 16543 29563
rect 16758 29560 16764 29572
rect 16531 29532 16764 29560
rect 16531 29529 16543 29532
rect 16485 29523 16543 29529
rect 16758 29520 16764 29532
rect 16816 29520 16822 29572
rect 17862 29520 17868 29572
rect 17920 29520 17926 29572
rect 18414 29520 18420 29572
rect 18472 29560 18478 29572
rect 18708 29560 18736 29600
rect 19889 29597 19901 29631
rect 19935 29628 19947 29631
rect 20806 29628 20812 29640
rect 19935 29600 20812 29628
rect 19935 29597 19947 29600
rect 19889 29591 19947 29597
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 20916 29628 20944 29727
rect 20990 29724 20996 29776
rect 21048 29764 21054 29776
rect 22465 29767 22523 29773
rect 22465 29764 22477 29767
rect 21048 29736 22477 29764
rect 21048 29724 21054 29736
rect 22465 29733 22477 29736
rect 22511 29733 22523 29767
rect 24581 29767 24639 29773
rect 24581 29764 24593 29767
rect 22465 29727 22523 29733
rect 22664 29736 24593 29764
rect 21453 29699 21511 29705
rect 21453 29665 21465 29699
rect 21499 29696 21511 29699
rect 22186 29696 22192 29708
rect 21499 29668 22192 29696
rect 21499 29665 21511 29668
rect 21453 29659 21511 29665
rect 22186 29656 22192 29668
rect 22244 29656 22250 29708
rect 21545 29631 21603 29637
rect 21545 29628 21557 29631
rect 20916 29600 21557 29628
rect 21545 29597 21557 29600
rect 21591 29597 21603 29631
rect 21545 29591 21603 29597
rect 18472 29532 18736 29560
rect 18472 29520 18478 29532
rect 19794 29520 19800 29572
rect 19852 29560 19858 29572
rect 19852 29532 21036 29560
rect 19852 29520 19858 29532
rect 9769 29495 9827 29501
rect 9769 29461 9781 29495
rect 9815 29492 9827 29495
rect 10318 29492 10324 29504
rect 9815 29464 10324 29492
rect 9815 29461 9827 29464
rect 9769 29455 9827 29461
rect 10318 29452 10324 29464
rect 10376 29452 10382 29504
rect 10870 29452 10876 29504
rect 10928 29452 10934 29504
rect 16942 29452 16948 29504
rect 17000 29492 17006 29504
rect 18969 29495 19027 29501
rect 18969 29492 18981 29495
rect 17000 29464 18981 29492
rect 17000 29452 17006 29464
rect 18969 29461 18981 29464
rect 19015 29492 19027 29495
rect 19058 29492 19064 29504
rect 19015 29464 19064 29492
rect 19015 29461 19027 29464
rect 18969 29455 19027 29461
rect 19058 29452 19064 29464
rect 19116 29452 19122 29504
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20257 29495 20315 29501
rect 20257 29492 20269 29495
rect 20036 29464 20269 29492
rect 20036 29452 20042 29464
rect 20257 29461 20269 29464
rect 20303 29461 20315 29495
rect 21008 29492 21036 29532
rect 21818 29520 21824 29572
rect 21876 29560 21882 29572
rect 22664 29560 22692 29736
rect 24581 29733 24593 29736
rect 24627 29733 24639 29767
rect 24581 29727 24639 29733
rect 22922 29656 22928 29708
rect 22980 29656 22986 29708
rect 23109 29699 23167 29705
rect 23109 29665 23121 29699
rect 23155 29696 23167 29699
rect 23474 29696 23480 29708
rect 23155 29668 23480 29696
rect 23155 29665 23167 29668
rect 23109 29659 23167 29665
rect 23474 29656 23480 29668
rect 23532 29656 23538 29708
rect 22738 29588 22744 29640
rect 22796 29628 22802 29640
rect 22833 29631 22891 29637
rect 22833 29628 22845 29631
rect 22796 29600 22845 29628
rect 22796 29588 22802 29600
rect 22833 29597 22845 29600
rect 22879 29597 22891 29631
rect 22833 29591 22891 29597
rect 23569 29631 23627 29637
rect 23569 29597 23581 29631
rect 23615 29628 23627 29631
rect 24029 29631 24087 29637
rect 24029 29628 24041 29631
rect 23615 29600 24041 29628
rect 23615 29597 23627 29600
rect 23569 29591 23627 29597
rect 24029 29597 24041 29600
rect 24075 29597 24087 29631
rect 24029 29591 24087 29597
rect 24044 29560 24072 29591
rect 24670 29588 24676 29640
rect 24728 29628 24734 29640
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 24728 29600 24777 29628
rect 24728 29588 24734 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 24765 29591 24823 29597
rect 24946 29560 24952 29572
rect 21876 29532 22692 29560
rect 22848 29532 23888 29560
rect 24044 29532 24952 29560
rect 21876 29520 21882 29532
rect 21450 29492 21456 29504
rect 21008 29464 21456 29492
rect 20257 29455 20315 29461
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 21634 29452 21640 29504
rect 21692 29452 21698 29504
rect 21910 29452 21916 29504
rect 21968 29492 21974 29504
rect 22848 29492 22876 29532
rect 23860 29501 23888 29532
rect 24946 29520 24952 29532
rect 25004 29520 25010 29572
rect 21968 29464 22876 29492
rect 23845 29495 23903 29501
rect 21968 29452 21974 29464
rect 23845 29461 23857 29495
rect 23891 29461 23903 29495
rect 23845 29455 23903 29461
rect 24670 29452 24676 29504
rect 24728 29492 24734 29504
rect 25041 29495 25099 29501
rect 25041 29492 25053 29495
rect 24728 29464 25053 29492
rect 24728 29452 24734 29464
rect 25041 29461 25053 29464
rect 25087 29461 25099 29495
rect 25041 29455 25099 29461
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 3559 29291 3617 29297
rect 3559 29257 3571 29291
rect 3605 29288 3617 29291
rect 3970 29288 3976 29300
rect 3605 29260 3976 29288
rect 3605 29257 3617 29260
rect 3559 29251 3617 29257
rect 3970 29248 3976 29260
rect 4028 29248 4034 29300
rect 8386 29248 8392 29300
rect 8444 29248 8450 29300
rect 8570 29248 8576 29300
rect 8628 29288 8634 29300
rect 8757 29291 8815 29297
rect 8757 29288 8769 29291
rect 8628 29260 8769 29288
rect 8628 29248 8634 29260
rect 8757 29257 8769 29260
rect 8803 29288 8815 29291
rect 9122 29288 9128 29300
rect 8803 29260 9128 29288
rect 8803 29257 8815 29260
rect 8757 29251 8815 29257
rect 9122 29248 9128 29260
rect 9180 29248 9186 29300
rect 12713 29291 12771 29297
rect 12713 29257 12725 29291
rect 12759 29288 12771 29291
rect 13817 29291 13875 29297
rect 13817 29288 13829 29291
rect 12759 29260 13829 29288
rect 12759 29257 12771 29260
rect 12713 29251 12771 29257
rect 13817 29257 13829 29260
rect 13863 29257 13875 29291
rect 13817 29251 13875 29257
rect 13909 29291 13967 29297
rect 13909 29257 13921 29291
rect 13955 29288 13967 29291
rect 15562 29288 15568 29300
rect 13955 29260 15568 29288
rect 13955 29257 13967 29260
rect 13909 29251 13967 29257
rect 15562 29248 15568 29260
rect 15620 29248 15626 29300
rect 15838 29248 15844 29300
rect 15896 29248 15902 29300
rect 17957 29291 18015 29297
rect 17957 29257 17969 29291
rect 18003 29288 18015 29291
rect 18693 29291 18751 29297
rect 18693 29288 18705 29291
rect 18003 29260 18705 29288
rect 18003 29257 18015 29260
rect 17957 29251 18015 29257
rect 18693 29257 18705 29260
rect 18739 29257 18751 29291
rect 18693 29251 18751 29257
rect 19153 29291 19211 29297
rect 19153 29257 19165 29291
rect 19199 29288 19211 29291
rect 20530 29288 20536 29300
rect 19199 29260 20536 29288
rect 19199 29257 19211 29260
rect 19153 29251 19211 29257
rect 20530 29248 20536 29260
rect 20588 29248 20594 29300
rect 21453 29291 21511 29297
rect 21453 29257 21465 29291
rect 21499 29288 21511 29291
rect 21634 29288 21640 29300
rect 21499 29260 21640 29288
rect 21499 29257 21511 29260
rect 21453 29251 21511 29257
rect 21634 29248 21640 29260
rect 21692 29248 21698 29300
rect 14182 29220 14188 29232
rect 12176 29192 14188 29220
rect 3488 29155 3546 29161
rect 3488 29121 3500 29155
rect 3534 29152 3546 29155
rect 3602 29152 3608 29164
rect 3534 29124 3608 29152
rect 3534 29121 3546 29124
rect 3488 29115 3546 29121
rect 3602 29112 3608 29124
rect 3660 29112 3666 29164
rect 7650 29112 7656 29164
rect 7708 29112 7714 29164
rect 10318 29112 10324 29164
rect 10376 29152 10382 29164
rect 11054 29152 11060 29164
rect 10376 29124 11060 29152
rect 10376 29112 10382 29124
rect 11054 29112 11060 29124
rect 11112 29112 11118 29164
rect 8849 29087 8907 29093
rect 8849 29053 8861 29087
rect 8895 29053 8907 29087
rect 8849 29047 8907 29053
rect 7374 28976 7380 29028
rect 7432 29016 7438 29028
rect 8021 29019 8079 29025
rect 8021 29016 8033 29019
rect 7432 28988 8033 29016
rect 7432 28976 7438 28988
rect 8021 28985 8033 28988
rect 8067 29016 8079 29019
rect 8864 29016 8892 29047
rect 8938 29044 8944 29096
rect 8996 29044 9002 29096
rect 12176 29093 12204 29192
rect 14182 29180 14188 29192
rect 14240 29180 14246 29232
rect 15378 29180 15384 29232
rect 15436 29220 15442 29232
rect 15654 29220 15660 29232
rect 15436 29192 15660 29220
rect 15436 29180 15442 29192
rect 15654 29180 15660 29192
rect 15712 29180 15718 29232
rect 15749 29223 15807 29229
rect 15749 29189 15761 29223
rect 15795 29220 15807 29223
rect 17034 29220 17040 29232
rect 15795 29192 17040 29220
rect 15795 29189 15807 29192
rect 15749 29183 15807 29189
rect 17034 29180 17040 29192
rect 17092 29180 17098 29232
rect 17865 29223 17923 29229
rect 17865 29189 17877 29223
rect 17911 29220 17923 29223
rect 20898 29220 20904 29232
rect 17911 29192 20904 29220
rect 17911 29189 17923 29192
rect 17865 29183 17923 29189
rect 20898 29180 20904 29192
rect 20956 29180 20962 29232
rect 23750 29180 23756 29232
rect 23808 29220 23814 29232
rect 24581 29223 24639 29229
rect 24581 29220 24593 29223
rect 23808 29192 24593 29220
rect 23808 29180 23814 29192
rect 24581 29189 24593 29192
rect 24627 29189 24639 29223
rect 24581 29183 24639 29189
rect 24762 29180 24768 29232
rect 24820 29180 24826 29232
rect 12342 29112 12348 29164
rect 12400 29112 12406 29164
rect 15562 29112 15568 29164
rect 15620 29152 15626 29164
rect 16850 29152 16856 29164
rect 15620 29124 16856 29152
rect 15620 29112 15626 29124
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 17494 29112 17500 29164
rect 17552 29152 17558 29164
rect 17552 29124 18184 29152
rect 17552 29112 17558 29124
rect 12161 29087 12219 29093
rect 12161 29053 12173 29087
rect 12207 29053 12219 29087
rect 12161 29047 12219 29053
rect 12253 29087 12311 29093
rect 12253 29053 12265 29087
rect 12299 29053 12311 29087
rect 12253 29047 12311 29053
rect 9398 29016 9404 29028
rect 8067 28988 9404 29016
rect 8067 28985 8079 28988
rect 8021 28979 8079 28985
rect 9398 28976 9404 28988
rect 9456 28976 9462 29028
rect 11422 28976 11428 29028
rect 11480 29016 11486 29028
rect 11609 29019 11667 29025
rect 11609 29016 11621 29019
rect 11480 28988 11621 29016
rect 11480 28976 11486 28988
rect 11609 28985 11621 28988
rect 11655 29016 11667 29019
rect 12268 29016 12296 29047
rect 14090 29044 14096 29096
rect 14148 29044 14154 29096
rect 15930 29044 15936 29096
rect 15988 29044 15994 29096
rect 16684 29056 17724 29084
rect 11655 28988 12296 29016
rect 11655 28985 11667 28988
rect 11609 28979 11667 28985
rect 12618 28976 12624 29028
rect 12676 29016 12682 29028
rect 13449 29019 13507 29025
rect 13449 29016 13461 29019
rect 12676 28988 13461 29016
rect 12676 28976 12682 28988
rect 13449 28985 13461 28988
rect 13495 28985 13507 29019
rect 13449 28979 13507 28985
rect 15378 28976 15384 29028
rect 15436 28976 15442 29028
rect 15654 28976 15660 29028
rect 15712 29016 15718 29028
rect 16684 29016 16712 29056
rect 15712 28988 16712 29016
rect 15712 28976 15718 28988
rect 16758 28976 16764 29028
rect 16816 28976 16822 29028
rect 17696 29016 17724 29056
rect 17770 29044 17776 29096
rect 17828 29084 17834 29096
rect 18049 29087 18107 29093
rect 18049 29084 18061 29087
rect 17828 29056 18061 29084
rect 17828 29044 17834 29056
rect 18049 29053 18061 29056
rect 18095 29053 18107 29087
rect 18156 29084 18184 29124
rect 19058 29112 19064 29164
rect 19116 29112 19122 29164
rect 19794 29152 19800 29164
rect 19168 29124 19800 29152
rect 19168 29084 19196 29124
rect 19794 29112 19800 29124
rect 19852 29152 19858 29164
rect 19889 29155 19947 29161
rect 19889 29152 19901 29155
rect 19852 29124 19901 29152
rect 19852 29112 19858 29124
rect 19889 29121 19901 29124
rect 19935 29121 19947 29155
rect 22005 29155 22063 29161
rect 22005 29152 22017 29155
rect 19889 29115 19947 29121
rect 20088 29124 22017 29152
rect 18156 29056 19196 29084
rect 19337 29087 19395 29093
rect 18049 29047 18107 29053
rect 19337 29053 19349 29087
rect 19383 29053 19395 29087
rect 19337 29047 19395 29053
rect 17696 28988 18276 29016
rect 7006 28908 7012 28960
rect 7064 28908 7070 28960
rect 9674 28908 9680 28960
rect 9732 28908 9738 28960
rect 17494 28908 17500 28960
rect 17552 28908 17558 28960
rect 18248 28948 18276 28988
rect 18322 28976 18328 29028
rect 18380 29016 18386 29028
rect 19352 29016 19380 29047
rect 19426 29044 19432 29096
rect 19484 29084 19490 29096
rect 20088 29084 20116 29124
rect 22005 29121 22017 29124
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 23293 29155 23351 29161
rect 23293 29121 23305 29155
rect 23339 29121 23351 29155
rect 23293 29115 23351 29121
rect 19484 29056 20116 29084
rect 20180 29056 22094 29084
rect 19484 29044 19490 29056
rect 19886 29016 19892 29028
rect 18380 28988 19288 29016
rect 19352 28988 19892 29016
rect 18380 28976 18386 28988
rect 18414 28948 18420 28960
rect 18248 28920 18420 28948
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 19260 28948 19288 28988
rect 19886 28976 19892 28988
rect 19944 28976 19950 29028
rect 20180 29016 20208 29056
rect 19996 28988 20208 29016
rect 22066 29016 22094 29056
rect 22370 29044 22376 29096
rect 22428 29084 22434 29096
rect 22649 29087 22707 29093
rect 22649 29084 22661 29087
rect 22428 29056 22661 29084
rect 22428 29044 22434 29056
rect 22649 29053 22661 29056
rect 22695 29053 22707 29087
rect 23308 29084 23336 29115
rect 23934 29112 23940 29164
rect 23992 29112 23998 29164
rect 23308 29056 24348 29084
rect 22649 29047 22707 29053
rect 24320 29028 24348 29056
rect 23109 29019 23167 29025
rect 23109 29016 23121 29019
rect 22066 28988 23121 29016
rect 19996 28948 20024 28988
rect 23109 28985 23121 28988
rect 23155 28985 23167 29019
rect 23109 28979 23167 28985
rect 23290 28976 23296 29028
rect 23348 29016 23354 29028
rect 23753 29019 23811 29025
rect 23753 29016 23765 29019
rect 23348 28988 23765 29016
rect 23348 28976 23354 28988
rect 23753 28985 23765 28988
rect 23799 28985 23811 29019
rect 23753 28979 23811 28985
rect 24302 28976 24308 29028
rect 24360 28976 24366 29028
rect 19260 28920 20024 28948
rect 20530 28908 20536 28960
rect 20588 28908 20594 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 18414 28744 18420 28756
rect 5736 28716 18420 28744
rect 5736 28620 5764 28716
rect 18414 28704 18420 28716
rect 18472 28704 18478 28756
rect 18877 28747 18935 28753
rect 18877 28713 18889 28747
rect 18923 28744 18935 28747
rect 18966 28744 18972 28756
rect 18923 28716 18972 28744
rect 18923 28713 18935 28716
rect 18877 28707 18935 28713
rect 11054 28636 11060 28688
rect 11112 28676 11118 28688
rect 18782 28676 18788 28688
rect 11112 28648 14872 28676
rect 11112 28636 11118 28648
rect 4154 28568 4160 28620
rect 4212 28608 4218 28620
rect 4249 28611 4307 28617
rect 4249 28608 4261 28611
rect 4212 28580 4261 28608
rect 4212 28568 4218 28580
rect 4249 28577 4261 28580
rect 4295 28577 4307 28611
rect 4249 28571 4307 28577
rect 5718 28568 5724 28620
rect 5776 28568 5782 28620
rect 11793 28611 11851 28617
rect 11793 28577 11805 28611
rect 11839 28608 11851 28611
rect 12342 28608 12348 28620
rect 11839 28580 12348 28608
rect 11839 28577 11851 28580
rect 11793 28571 11851 28577
rect 12342 28568 12348 28580
rect 12400 28568 12406 28620
rect 12802 28568 12808 28620
rect 12860 28568 12866 28620
rect 14090 28568 14096 28620
rect 14148 28608 14154 28620
rect 14734 28608 14740 28620
rect 14148 28580 14740 28608
rect 14148 28568 14154 28580
rect 14734 28568 14740 28580
rect 14792 28568 14798 28620
rect 14844 28617 14872 28648
rect 18064 28648 18788 28676
rect 14829 28611 14887 28617
rect 14829 28577 14841 28611
rect 14875 28577 14887 28611
rect 14829 28571 14887 28577
rect 16574 28568 16580 28620
rect 16632 28568 16638 28620
rect 16669 28611 16727 28617
rect 16669 28577 16681 28611
rect 16715 28608 16727 28611
rect 17586 28608 17592 28620
rect 16715 28580 17592 28608
rect 16715 28577 16727 28580
rect 16669 28571 16727 28577
rect 17586 28568 17592 28580
rect 17644 28568 17650 28620
rect 18064 28617 18092 28648
rect 18782 28636 18788 28648
rect 18840 28676 18846 28688
rect 18892 28676 18920 28707
rect 18966 28704 18972 28716
rect 19024 28704 19030 28756
rect 22554 28704 22560 28756
rect 22612 28744 22618 28756
rect 22738 28744 22744 28756
rect 22612 28716 22744 28744
rect 22612 28704 22618 28716
rect 22738 28704 22744 28716
rect 22796 28704 22802 28756
rect 18840 28648 18920 28676
rect 18840 28636 18846 28648
rect 18049 28611 18107 28617
rect 18049 28577 18061 28611
rect 18095 28577 18107 28611
rect 18049 28571 18107 28577
rect 18230 28568 18236 28620
rect 18288 28568 18294 28620
rect 18414 28568 18420 28620
rect 18472 28608 18478 28620
rect 18969 28611 19027 28617
rect 18969 28608 18981 28611
rect 18472 28580 18981 28608
rect 18472 28568 18478 28580
rect 18969 28577 18981 28580
rect 19015 28608 19027 28611
rect 19058 28608 19064 28620
rect 19015 28580 19064 28608
rect 19015 28577 19027 28580
rect 18969 28571 19027 28577
rect 19058 28568 19064 28580
rect 19116 28568 19122 28620
rect 20530 28568 20536 28620
rect 20588 28608 20594 28620
rect 20901 28611 20959 28617
rect 20901 28608 20913 28611
rect 20588 28580 20913 28608
rect 20588 28568 20594 28580
rect 20901 28577 20913 28580
rect 20947 28577 20959 28611
rect 20901 28571 20959 28577
rect 8570 28500 8576 28552
rect 8628 28500 8634 28552
rect 9766 28500 9772 28552
rect 9824 28500 9830 28552
rect 11514 28500 11520 28552
rect 11572 28540 11578 28552
rect 12713 28543 12771 28549
rect 12713 28540 12725 28543
rect 11572 28512 12725 28540
rect 11572 28500 11578 28512
rect 12713 28509 12725 28512
rect 12759 28540 12771 28543
rect 13541 28543 13599 28549
rect 13541 28540 13553 28543
rect 12759 28512 13553 28540
rect 12759 28509 12771 28512
rect 12713 28503 12771 28509
rect 13541 28509 13553 28512
rect 13587 28540 13599 28543
rect 16761 28543 16819 28549
rect 13587 28512 15700 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 3418 28432 3424 28484
rect 3476 28472 3482 28484
rect 4433 28475 4491 28481
rect 4433 28472 4445 28475
rect 3476 28444 4445 28472
rect 3476 28432 3482 28444
rect 4433 28441 4445 28444
rect 4479 28441 4491 28475
rect 4433 28435 4491 28441
rect 7742 28432 7748 28484
rect 7800 28432 7806 28484
rect 8297 28475 8355 28481
rect 8297 28441 8309 28475
rect 8343 28472 8355 28475
rect 9125 28475 9183 28481
rect 9125 28472 9137 28475
rect 8343 28444 9137 28472
rect 8343 28441 8355 28444
rect 8297 28435 8355 28441
rect 9125 28441 9137 28444
rect 9171 28441 9183 28475
rect 9125 28435 9183 28441
rect 14645 28475 14703 28481
rect 14645 28441 14657 28475
rect 14691 28472 14703 28475
rect 15672 28472 15700 28512
rect 16761 28509 16773 28543
rect 16807 28540 16819 28543
rect 17494 28540 17500 28552
rect 16807 28512 17500 28540
rect 16807 28509 16819 28512
rect 16761 28503 16819 28509
rect 17494 28500 17500 28512
rect 17552 28500 17558 28552
rect 17957 28543 18015 28549
rect 17957 28509 17969 28543
rect 18003 28540 18015 28543
rect 18601 28543 18659 28549
rect 18601 28540 18613 28543
rect 18003 28512 18613 28540
rect 18003 28509 18015 28512
rect 17957 28503 18015 28509
rect 18601 28509 18613 28512
rect 18647 28509 18659 28543
rect 18601 28503 18659 28509
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28540 21235 28543
rect 22186 28540 22192 28552
rect 21223 28512 22192 28540
rect 21223 28509 21235 28512
rect 21177 28503 21235 28509
rect 15746 28472 15752 28484
rect 14691 28444 15608 28472
rect 15672 28444 15752 28472
rect 14691 28441 14703 28444
rect 14645 28435 14703 28441
rect 15580 28416 15608 28444
rect 15746 28432 15752 28444
rect 15804 28472 15810 28484
rect 17972 28472 18000 28503
rect 22186 28500 22192 28512
rect 22244 28540 22250 28552
rect 22281 28543 22339 28549
rect 22281 28540 22293 28543
rect 22244 28512 22293 28540
rect 22244 28500 22250 28512
rect 22281 28509 22293 28512
rect 22327 28509 22339 28543
rect 22281 28503 22339 28509
rect 24394 28500 24400 28552
rect 24452 28540 24458 28552
rect 24673 28543 24731 28549
rect 24673 28540 24685 28543
rect 24452 28512 24685 28540
rect 24452 28500 24458 28512
rect 24673 28509 24685 28512
rect 24719 28509 24731 28543
rect 24673 28503 24731 28509
rect 21453 28475 21511 28481
rect 21453 28472 21465 28475
rect 15804 28444 18000 28472
rect 18064 28444 19564 28472
rect 20470 28444 21465 28472
rect 15804 28432 15810 28444
rect 6825 28407 6883 28413
rect 6825 28373 6837 28407
rect 6871 28404 6883 28407
rect 7650 28404 7656 28416
rect 6871 28376 7656 28404
rect 6871 28373 6883 28376
rect 6825 28367 6883 28373
rect 7650 28364 7656 28376
rect 7708 28364 7714 28416
rect 10870 28364 10876 28416
rect 10928 28404 10934 28416
rect 12253 28407 12311 28413
rect 12253 28404 12265 28407
rect 10928 28376 12265 28404
rect 10928 28364 10934 28376
rect 12253 28373 12265 28376
rect 12299 28373 12311 28407
rect 12253 28367 12311 28373
rect 12621 28407 12679 28413
rect 12621 28373 12633 28407
rect 12667 28404 12679 28407
rect 13357 28407 13415 28413
rect 13357 28404 13369 28407
rect 12667 28376 13369 28404
rect 12667 28373 12679 28376
rect 12621 28367 12679 28373
rect 13357 28373 13369 28376
rect 13403 28404 13415 28407
rect 13446 28404 13452 28416
rect 13403 28376 13452 28404
rect 13403 28373 13415 28376
rect 13357 28367 13415 28373
rect 13446 28364 13452 28376
rect 13504 28364 13510 28416
rect 13538 28364 13544 28416
rect 13596 28404 13602 28416
rect 14277 28407 14335 28413
rect 14277 28404 14289 28407
rect 13596 28376 14289 28404
rect 13596 28364 13602 28376
rect 14277 28373 14289 28376
rect 14323 28373 14335 28407
rect 14277 28367 14335 28373
rect 14734 28364 14740 28416
rect 14792 28404 14798 28416
rect 15289 28407 15347 28413
rect 15289 28404 15301 28407
rect 14792 28376 15301 28404
rect 14792 28364 14798 28376
rect 15289 28373 15301 28376
rect 15335 28373 15347 28407
rect 15289 28367 15347 28373
rect 15562 28364 15568 28416
rect 15620 28364 15626 28416
rect 17034 28364 17040 28416
rect 17092 28404 17098 28416
rect 17129 28407 17187 28413
rect 17129 28404 17141 28407
rect 17092 28376 17141 28404
rect 17092 28364 17098 28376
rect 17129 28373 17141 28376
rect 17175 28373 17187 28407
rect 17129 28367 17187 28373
rect 17586 28364 17592 28416
rect 17644 28364 17650 28416
rect 17678 28364 17684 28416
rect 17736 28404 17742 28416
rect 18064 28404 18092 28444
rect 17736 28376 18092 28404
rect 17736 28364 17742 28376
rect 18230 28364 18236 28416
rect 18288 28404 18294 28416
rect 18414 28404 18420 28416
rect 18288 28376 18420 28404
rect 18288 28364 18294 28376
rect 18414 28364 18420 28376
rect 18472 28404 18478 28416
rect 19242 28404 19248 28416
rect 18472 28376 19248 28404
rect 18472 28364 18478 28376
rect 19242 28364 19248 28376
rect 19300 28364 19306 28416
rect 19426 28364 19432 28416
rect 19484 28364 19490 28416
rect 19536 28404 19564 28444
rect 20548 28404 20576 28444
rect 21453 28441 21465 28444
rect 21499 28472 21511 28475
rect 21542 28472 21548 28484
rect 21499 28444 21548 28472
rect 21499 28441 21511 28444
rect 21453 28435 21511 28441
rect 21542 28432 21548 28444
rect 21600 28432 21606 28484
rect 22462 28432 22468 28484
rect 22520 28472 22526 28484
rect 22557 28475 22615 28481
rect 22557 28472 22569 28475
rect 22520 28444 22569 28472
rect 22520 28432 22526 28444
rect 22557 28441 22569 28444
rect 22603 28441 22615 28475
rect 22557 28435 22615 28441
rect 23014 28432 23020 28484
rect 23072 28432 23078 28484
rect 24857 28475 24915 28481
rect 24857 28441 24869 28475
rect 24903 28472 24915 28475
rect 25130 28472 25136 28484
rect 24903 28444 25136 28472
rect 24903 28441 24915 28444
rect 24857 28435 24915 28441
rect 25130 28432 25136 28444
rect 25188 28432 25194 28484
rect 19536 28376 20576 28404
rect 23474 28364 23480 28416
rect 23532 28404 23538 28416
rect 24029 28407 24087 28413
rect 24029 28404 24041 28407
rect 23532 28376 24041 28404
rect 23532 28364 23538 28376
rect 24029 28373 24041 28376
rect 24075 28404 24087 28407
rect 24302 28404 24308 28416
rect 24075 28376 24308 28404
rect 24075 28373 24087 28376
rect 24029 28367 24087 28373
rect 24302 28364 24308 28376
rect 24360 28364 24366 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 7834 28160 7840 28212
rect 7892 28200 7898 28212
rect 8573 28203 8631 28209
rect 8573 28200 8585 28203
rect 7892 28172 8585 28200
rect 7892 28160 7898 28172
rect 8573 28169 8585 28172
rect 8619 28200 8631 28203
rect 12802 28200 12808 28212
rect 8619 28172 12808 28200
rect 8619 28169 8631 28172
rect 8573 28163 8631 28169
rect 12802 28160 12808 28172
rect 12860 28160 12866 28212
rect 13446 28160 13452 28212
rect 13504 28200 13510 28212
rect 15654 28200 15660 28212
rect 13504 28172 15660 28200
rect 13504 28160 13510 28172
rect 15654 28160 15660 28172
rect 15712 28160 15718 28212
rect 16574 28160 16580 28212
rect 16632 28200 16638 28212
rect 17037 28203 17095 28209
rect 17037 28200 17049 28203
rect 16632 28172 17049 28200
rect 16632 28160 16638 28172
rect 17037 28169 17049 28172
rect 17083 28200 17095 28203
rect 17678 28200 17684 28212
rect 17083 28172 17684 28200
rect 17083 28169 17095 28172
rect 17037 28163 17095 28169
rect 17678 28160 17684 28172
rect 17736 28160 17742 28212
rect 18230 28160 18236 28212
rect 18288 28200 18294 28212
rect 18414 28200 18420 28212
rect 18288 28172 18420 28200
rect 18288 28160 18294 28172
rect 18414 28160 18420 28172
rect 18472 28160 18478 28212
rect 18966 28160 18972 28212
rect 19024 28200 19030 28212
rect 19702 28200 19708 28212
rect 19024 28172 19708 28200
rect 19024 28160 19030 28172
rect 19702 28160 19708 28172
rect 19760 28160 19766 28212
rect 19886 28160 19892 28212
rect 19944 28200 19950 28212
rect 22097 28203 22155 28209
rect 22097 28200 22109 28203
rect 19944 28172 22109 28200
rect 19944 28160 19950 28172
rect 22097 28169 22109 28172
rect 22143 28169 22155 28203
rect 23290 28200 23296 28212
rect 22097 28163 22155 28169
rect 22296 28172 23296 28200
rect 7006 28092 7012 28144
rect 7064 28132 7070 28144
rect 7101 28135 7159 28141
rect 7101 28132 7113 28135
rect 7064 28104 7113 28132
rect 7064 28092 7070 28104
rect 7101 28101 7113 28104
rect 7147 28101 7159 28135
rect 7101 28095 7159 28101
rect 7742 28092 7748 28144
rect 7800 28092 7806 28144
rect 10505 28135 10563 28141
rect 10505 28101 10517 28135
rect 10551 28132 10563 28135
rect 11701 28135 11759 28141
rect 11701 28132 11713 28135
rect 10551 28104 11713 28132
rect 10551 28101 10563 28104
rect 10505 28095 10563 28101
rect 11701 28101 11713 28104
rect 11747 28101 11759 28135
rect 11701 28095 11759 28101
rect 13081 28135 13139 28141
rect 13081 28101 13093 28135
rect 13127 28132 13139 28135
rect 13354 28132 13360 28144
rect 13127 28104 13360 28132
rect 13127 28101 13139 28104
rect 13081 28095 13139 28101
rect 13354 28092 13360 28104
rect 13412 28092 13418 28144
rect 14458 28132 14464 28144
rect 14306 28104 14464 28132
rect 14458 28092 14464 28104
rect 14516 28092 14522 28144
rect 17494 28092 17500 28144
rect 17552 28132 17558 28144
rect 17773 28135 17831 28141
rect 17773 28132 17785 28135
rect 17552 28104 17785 28132
rect 17552 28092 17558 28104
rect 17773 28101 17785 28104
rect 17819 28132 17831 28135
rect 18601 28135 18659 28141
rect 18601 28132 18613 28135
rect 17819 28104 18613 28132
rect 17819 28101 17831 28104
rect 17773 28095 17831 28101
rect 18601 28101 18613 28104
rect 18647 28132 18659 28135
rect 21174 28132 21180 28144
rect 18647 28104 21180 28132
rect 18647 28101 18659 28104
rect 18601 28095 18659 28101
rect 21174 28092 21180 28104
rect 21232 28092 21238 28144
rect 8956 28036 9430 28064
rect 6822 27956 6828 28008
rect 6880 27956 6886 28008
rect 7742 27956 7748 28008
rect 7800 27996 7806 28008
rect 8956 27996 8984 28036
rect 12342 28024 12348 28076
rect 12400 28024 12406 28076
rect 15657 28067 15715 28073
rect 15657 28064 15669 28067
rect 14568 28036 15669 28064
rect 7800 27968 8984 27996
rect 9033 27999 9091 28005
rect 7800 27956 7806 27968
rect 9033 27965 9045 27999
rect 9079 27996 9091 27999
rect 9766 27996 9772 28008
rect 9079 27968 9772 27996
rect 9079 27965 9091 27968
rect 9033 27959 9091 27965
rect 9766 27956 9772 27968
rect 9824 27956 9830 28008
rect 10781 27999 10839 28005
rect 10781 27965 10793 27999
rect 10827 27996 10839 27999
rect 12434 27996 12440 28008
rect 10827 27968 12440 27996
rect 10827 27965 10839 27968
rect 10781 27959 10839 27965
rect 12434 27956 12440 27968
rect 12492 27996 12498 28008
rect 12805 27999 12863 28005
rect 12805 27996 12817 27999
rect 12492 27968 12817 27996
rect 12492 27956 12498 27968
rect 12805 27965 12817 27968
rect 12851 27965 12863 27999
rect 12805 27959 12863 27965
rect 14274 27820 14280 27872
rect 14332 27860 14338 27872
rect 14568 27869 14596 28036
rect 15657 28033 15669 28036
rect 15703 28064 15715 28067
rect 15930 28064 15936 28076
rect 15703 28036 15936 28064
rect 15703 28033 15715 28036
rect 15657 28027 15715 28033
rect 15930 28024 15936 28036
rect 15988 28024 15994 28076
rect 17862 28064 17868 28076
rect 17144 28036 17868 28064
rect 16298 27888 16304 27940
rect 16356 27928 16362 27940
rect 17144 27937 17172 28036
rect 17862 28024 17868 28036
rect 17920 28024 17926 28076
rect 19242 28024 19248 28076
rect 19300 28064 19306 28076
rect 19797 28067 19855 28073
rect 19797 28064 19809 28067
rect 19300 28036 19809 28064
rect 19300 28024 19306 28036
rect 19797 28033 19809 28036
rect 19843 28033 19855 28067
rect 21358 28064 21364 28076
rect 19797 28027 19855 28033
rect 19904 28036 21364 28064
rect 17681 27999 17739 28005
rect 17681 27965 17693 27999
rect 17727 27996 17739 27999
rect 18598 27996 18604 28008
rect 17727 27968 18604 27996
rect 17727 27965 17739 27968
rect 17681 27959 17739 27965
rect 18598 27956 18604 27968
rect 18656 27996 18662 28008
rect 18874 27996 18880 28008
rect 18656 27968 18880 27996
rect 18656 27956 18662 27968
rect 18874 27956 18880 27968
rect 18932 27956 18938 28008
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27996 19671 27999
rect 19702 27996 19708 28008
rect 19659 27968 19708 27996
rect 19659 27965 19671 27968
rect 19613 27959 19671 27965
rect 19702 27956 19708 27968
rect 19760 27956 19766 28008
rect 17129 27931 17187 27937
rect 17129 27928 17141 27931
rect 16356 27900 17141 27928
rect 16356 27888 16362 27900
rect 17129 27897 17141 27900
rect 17175 27897 17187 27931
rect 19904 27928 19932 28036
rect 21358 28024 21364 28036
rect 21416 28024 21422 28076
rect 21453 28067 21511 28073
rect 21453 28033 21465 28067
rect 21499 28064 21511 28067
rect 22296 28064 22324 28172
rect 23290 28160 23296 28172
rect 23348 28160 23354 28212
rect 24118 28092 24124 28144
rect 24176 28132 24182 28144
rect 24765 28135 24823 28141
rect 24765 28132 24777 28135
rect 24176 28104 24777 28132
rect 24176 28092 24182 28104
rect 24765 28101 24777 28104
rect 24811 28101 24823 28135
rect 24765 28095 24823 28101
rect 21499 28036 22324 28064
rect 21499 28033 21511 28036
rect 21453 28027 21511 28033
rect 22462 28024 22468 28076
rect 22520 28024 22526 28076
rect 21174 27956 21180 28008
rect 21232 27956 21238 28008
rect 22480 27996 22508 28024
rect 23014 27996 23020 28008
rect 22480 27968 23020 27996
rect 23014 27956 23020 27968
rect 23072 27956 23078 28008
rect 23566 27956 23572 28008
rect 23624 27956 23630 28008
rect 23845 27999 23903 28005
rect 23845 27965 23857 27999
rect 23891 27965 23903 27999
rect 23845 27959 23903 27965
rect 22002 27928 22008 27940
rect 17129 27891 17187 27897
rect 18156 27900 19932 27928
rect 20088 27900 22008 27928
rect 14553 27863 14611 27869
rect 14553 27860 14565 27863
rect 14332 27832 14565 27860
rect 14332 27820 14338 27832
rect 14553 27829 14565 27832
rect 14599 27829 14611 27863
rect 14553 27823 14611 27829
rect 15010 27820 15016 27872
rect 15068 27820 15074 27872
rect 16390 27820 16396 27872
rect 16448 27860 16454 27872
rect 18156 27860 18184 27900
rect 16448 27832 18184 27860
rect 18233 27863 18291 27869
rect 16448 27820 16454 27832
rect 18233 27829 18245 27863
rect 18279 27860 18291 27863
rect 18322 27860 18328 27872
rect 18279 27832 18328 27860
rect 18279 27829 18291 27832
rect 18233 27823 18291 27829
rect 18322 27820 18328 27832
rect 18380 27820 18386 27872
rect 18874 27820 18880 27872
rect 18932 27860 18938 27872
rect 19061 27863 19119 27869
rect 19061 27860 19073 27863
rect 18932 27832 19073 27860
rect 18932 27820 18938 27832
rect 19061 27829 19073 27832
rect 19107 27860 19119 27863
rect 19242 27860 19248 27872
rect 19107 27832 19248 27860
rect 19107 27829 19119 27832
rect 19061 27823 19119 27829
rect 19242 27820 19248 27832
rect 19300 27820 19306 27872
rect 19702 27820 19708 27872
rect 19760 27860 19766 27872
rect 20088 27860 20116 27900
rect 22002 27888 22008 27900
rect 22060 27888 22066 27940
rect 19760 27832 20116 27860
rect 20165 27863 20223 27869
rect 19760 27820 19766 27832
rect 20165 27829 20177 27863
rect 20211 27860 20223 27863
rect 20622 27860 20628 27872
rect 20211 27832 20628 27860
rect 20211 27829 20223 27832
rect 20165 27823 20223 27829
rect 20622 27820 20628 27832
rect 20680 27820 20686 27872
rect 23382 27820 23388 27872
rect 23440 27860 23446 27872
rect 23860 27860 23888 27959
rect 24578 27888 24584 27940
rect 24636 27888 24642 27940
rect 23440 27832 23888 27860
rect 23440 27820 23446 27832
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 9572 27659 9630 27665
rect 9572 27625 9584 27659
rect 9618 27656 9630 27659
rect 9674 27656 9680 27668
rect 9618 27628 9680 27656
rect 9618 27625 9630 27628
rect 9572 27619 9630 27625
rect 9674 27616 9680 27628
rect 9732 27616 9738 27668
rect 11057 27659 11115 27665
rect 11057 27625 11069 27659
rect 11103 27656 11115 27659
rect 12342 27656 12348 27668
rect 11103 27628 12348 27656
rect 11103 27625 11115 27628
rect 11057 27619 11115 27625
rect 12342 27616 12348 27628
rect 12400 27616 12406 27668
rect 14090 27616 14096 27668
rect 14148 27656 14154 27668
rect 16850 27656 16856 27668
rect 14148 27628 16856 27656
rect 14148 27616 14154 27628
rect 16850 27616 16856 27628
rect 16908 27656 16914 27668
rect 19794 27656 19800 27668
rect 16908 27628 19800 27656
rect 16908 27616 16914 27628
rect 19794 27616 19800 27628
rect 19852 27656 19858 27668
rect 19852 27628 20484 27656
rect 19852 27616 19858 27628
rect 12250 27548 12256 27600
rect 12308 27588 12314 27600
rect 12989 27591 13047 27597
rect 12989 27588 13001 27591
rect 12308 27560 13001 27588
rect 12308 27548 12314 27560
rect 12989 27557 13001 27560
rect 13035 27557 13047 27591
rect 12989 27551 13047 27557
rect 16945 27591 17003 27597
rect 16945 27557 16957 27591
rect 16991 27588 17003 27591
rect 17402 27588 17408 27600
rect 16991 27560 17408 27588
rect 16991 27557 17003 27560
rect 16945 27551 17003 27557
rect 17402 27548 17408 27560
rect 17460 27588 17466 27600
rect 17678 27588 17684 27600
rect 17460 27560 17684 27588
rect 17460 27548 17466 27560
rect 17678 27548 17684 27560
rect 17736 27548 17742 27600
rect 18877 27591 18935 27597
rect 18877 27557 18889 27591
rect 18923 27588 18935 27591
rect 20254 27588 20260 27600
rect 18923 27560 20260 27588
rect 18923 27557 18935 27560
rect 18877 27551 18935 27557
rect 20254 27548 20260 27560
rect 20312 27548 20318 27600
rect 20456 27597 20484 27628
rect 20441 27591 20499 27597
rect 20441 27557 20453 27591
rect 20487 27557 20499 27591
rect 20441 27551 20499 27557
rect 2774 27480 2780 27532
rect 2832 27480 2838 27532
rect 3237 27523 3295 27529
rect 3237 27489 3249 27523
rect 3283 27520 3295 27523
rect 3602 27520 3608 27532
rect 3283 27492 3608 27520
rect 3283 27489 3295 27492
rect 3237 27483 3295 27489
rect 3602 27480 3608 27492
rect 3660 27480 3666 27532
rect 3878 27480 3884 27532
rect 3936 27520 3942 27532
rect 3973 27523 4031 27529
rect 3973 27520 3985 27523
rect 3936 27492 3985 27520
rect 3936 27480 3942 27492
rect 3973 27489 3985 27492
rect 4019 27489 4031 27523
rect 3973 27483 4031 27489
rect 7650 27480 7656 27532
rect 7708 27520 7714 27532
rect 11701 27523 11759 27529
rect 11701 27520 11713 27523
rect 7708 27492 11713 27520
rect 7708 27480 7714 27492
rect 11701 27489 11713 27492
rect 11747 27489 11759 27523
rect 11701 27483 11759 27489
rect 11885 27523 11943 27529
rect 11885 27489 11897 27523
rect 11931 27520 11943 27523
rect 12066 27520 12072 27532
rect 11931 27492 12072 27520
rect 11931 27489 11943 27492
rect 11885 27483 11943 27489
rect 12066 27480 12072 27492
rect 12124 27480 12130 27532
rect 13541 27523 13599 27529
rect 13541 27520 13553 27523
rect 12406 27492 13553 27520
rect 3421 27455 3479 27461
rect 3421 27421 3433 27455
rect 3467 27421 3479 27455
rect 3421 27415 3479 27421
rect 7469 27455 7527 27461
rect 7469 27421 7481 27455
rect 7515 27421 7527 27455
rect 7469 27415 7527 27421
rect 3436 27316 3464 27415
rect 4157 27387 4215 27393
rect 4157 27353 4169 27387
rect 4203 27384 4215 27387
rect 4246 27384 4252 27396
rect 4203 27356 4252 27384
rect 4203 27353 4215 27356
rect 4157 27347 4215 27353
rect 4246 27344 4252 27356
rect 4304 27344 4310 27396
rect 5813 27387 5871 27393
rect 5813 27353 5825 27387
rect 5859 27384 5871 27387
rect 5902 27384 5908 27396
rect 5859 27356 5908 27384
rect 5859 27353 5871 27356
rect 5813 27347 5871 27353
rect 5902 27344 5908 27356
rect 5960 27344 5966 27396
rect 6546 27344 6552 27396
rect 6604 27384 6610 27396
rect 7484 27384 7512 27415
rect 9306 27412 9312 27464
rect 9364 27412 9370 27464
rect 9490 27384 9496 27396
rect 6604 27356 9496 27384
rect 6604 27344 6610 27356
rect 9490 27344 9496 27356
rect 9548 27344 9554 27396
rect 11146 27384 11152 27396
rect 10810 27356 11152 27384
rect 11146 27344 11152 27356
rect 11204 27344 11210 27396
rect 12406 27384 12434 27492
rect 13541 27489 13553 27492
rect 13587 27489 13599 27523
rect 13541 27483 13599 27489
rect 13630 27480 13636 27532
rect 13688 27520 13694 27532
rect 14918 27520 14924 27532
rect 13688 27492 14924 27520
rect 13688 27480 13694 27492
rect 14918 27480 14924 27492
rect 14976 27480 14982 27532
rect 15197 27523 15255 27529
rect 15197 27489 15209 27523
rect 15243 27520 15255 27523
rect 16114 27520 16120 27532
rect 15243 27492 16120 27520
rect 15243 27489 15255 27492
rect 15197 27483 15255 27489
rect 16114 27480 16120 27492
rect 16172 27480 16178 27532
rect 17586 27480 17592 27532
rect 17644 27520 17650 27532
rect 17957 27523 18015 27529
rect 17957 27520 17969 27523
rect 17644 27492 17969 27520
rect 17644 27480 17650 27492
rect 17957 27489 17969 27492
rect 18003 27489 18015 27523
rect 17957 27483 18015 27489
rect 18049 27523 18107 27529
rect 18049 27489 18061 27523
rect 18095 27489 18107 27523
rect 18049 27483 18107 27489
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 14182 27452 14188 27464
rect 13403 27424 14188 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 14182 27412 14188 27424
rect 14240 27412 14246 27464
rect 16574 27412 16580 27464
rect 16632 27412 16638 27464
rect 17862 27412 17868 27464
rect 17920 27452 17926 27464
rect 18064 27452 18092 27483
rect 18230 27480 18236 27532
rect 18288 27520 18294 27532
rect 19613 27523 19671 27529
rect 18288 27492 18920 27520
rect 18288 27480 18294 27492
rect 18892 27464 18920 27492
rect 19613 27489 19625 27523
rect 19659 27520 19671 27523
rect 19659 27492 20024 27520
rect 19659 27489 19671 27492
rect 19613 27483 19671 27489
rect 17920 27424 18092 27452
rect 18693 27455 18751 27461
rect 17920 27412 17926 27424
rect 18693 27421 18705 27455
rect 18739 27421 18751 27455
rect 18693 27415 18751 27421
rect 14277 27387 14335 27393
rect 14277 27384 14289 27387
rect 11256 27356 12434 27384
rect 13464 27356 14289 27384
rect 4522 27316 4528 27328
rect 3436 27288 4528 27316
rect 4522 27276 4528 27288
rect 4580 27276 4586 27328
rect 6825 27319 6883 27325
rect 6825 27285 6837 27319
rect 6871 27316 6883 27319
rect 7098 27316 7104 27328
rect 6871 27288 7104 27316
rect 6871 27285 6883 27288
rect 6825 27279 6883 27285
rect 7098 27276 7104 27288
rect 7156 27276 7162 27328
rect 8846 27276 8852 27328
rect 8904 27316 8910 27328
rect 11256 27316 11284 27356
rect 13464 27328 13492 27356
rect 14277 27353 14289 27356
rect 14323 27384 14335 27387
rect 15102 27384 15108 27396
rect 14323 27356 15108 27384
rect 14323 27353 14335 27356
rect 14277 27347 14335 27353
rect 15102 27344 15108 27356
rect 15160 27344 15166 27396
rect 15470 27344 15476 27396
rect 15528 27344 15534 27396
rect 18708 27384 18736 27415
rect 18874 27412 18880 27464
rect 18932 27412 18938 27464
rect 19794 27412 19800 27464
rect 19852 27412 19858 27464
rect 16776 27356 18736 27384
rect 19996 27384 20024 27492
rect 20070 27480 20076 27532
rect 20128 27520 20134 27532
rect 21637 27523 21695 27529
rect 21637 27520 21649 27523
rect 20128 27492 21649 27520
rect 20128 27480 20134 27492
rect 21637 27489 21649 27492
rect 21683 27520 21695 27523
rect 22554 27520 22560 27532
rect 21683 27492 22560 27520
rect 21683 27489 21695 27492
rect 21637 27483 21695 27489
rect 22554 27480 22560 27492
rect 22612 27480 22618 27532
rect 23109 27523 23167 27529
rect 23109 27489 23121 27523
rect 23155 27520 23167 27523
rect 23842 27520 23848 27532
rect 23155 27492 23848 27520
rect 23155 27489 23167 27492
rect 23109 27483 23167 27489
rect 23842 27480 23848 27492
rect 23900 27480 23906 27532
rect 21085 27455 21143 27461
rect 21085 27421 21097 27455
rect 21131 27452 21143 27455
rect 21358 27452 21364 27464
rect 21131 27424 21364 27452
rect 21131 27421 21143 27424
rect 21085 27415 21143 27421
rect 21358 27412 21364 27424
rect 21416 27412 21422 27464
rect 23382 27412 23388 27464
rect 23440 27412 23446 27464
rect 24302 27412 24308 27464
rect 24360 27452 24366 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24360 27424 24593 27452
rect 24360 27412 24366 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 20530 27384 20536 27396
rect 19996 27356 20536 27384
rect 8904 27288 11284 27316
rect 8904 27276 8910 27288
rect 11974 27276 11980 27328
rect 12032 27276 12038 27328
rect 12345 27319 12403 27325
rect 12345 27285 12357 27319
rect 12391 27316 12403 27319
rect 12710 27316 12716 27328
rect 12391 27288 12716 27316
rect 12391 27285 12403 27288
rect 12345 27279 12403 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 13446 27276 13452 27328
rect 13504 27276 13510 27328
rect 14182 27276 14188 27328
rect 14240 27276 14246 27328
rect 14458 27276 14464 27328
rect 14516 27316 14522 27328
rect 14645 27319 14703 27325
rect 14645 27316 14657 27319
rect 14516 27288 14657 27316
rect 14516 27276 14522 27288
rect 14645 27285 14657 27288
rect 14691 27285 14703 27319
rect 14645 27279 14703 27285
rect 14826 27276 14832 27328
rect 14884 27316 14890 27328
rect 16776 27316 16804 27356
rect 20530 27344 20536 27356
rect 20588 27384 20594 27396
rect 21266 27384 21272 27396
rect 20588 27356 21272 27384
rect 20588 27344 20594 27356
rect 21266 27344 21272 27356
rect 21324 27344 21330 27396
rect 22554 27344 22560 27396
rect 22612 27344 22618 27396
rect 23400 27384 23428 27412
rect 23308 27356 23428 27384
rect 14884 27288 16804 27316
rect 14884 27276 14890 27288
rect 17494 27276 17500 27328
rect 17552 27276 17558 27328
rect 17865 27319 17923 27325
rect 17865 27285 17877 27319
rect 17911 27316 17923 27319
rect 19334 27316 19340 27328
rect 17911 27288 19340 27316
rect 17911 27285 17923 27288
rect 17865 27279 17923 27285
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 19702 27276 19708 27328
rect 19760 27276 19766 27328
rect 20162 27276 20168 27328
rect 20220 27276 20226 27328
rect 20898 27276 20904 27328
rect 20956 27276 20962 27328
rect 22186 27276 22192 27328
rect 22244 27316 22250 27328
rect 23308 27316 23336 27356
rect 22244 27288 23336 27316
rect 22244 27276 22250 27288
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 23845 27319 23903 27325
rect 23845 27316 23857 27319
rect 23532 27288 23857 27316
rect 23532 27276 23538 27288
rect 23845 27285 23857 27288
rect 23891 27285 23903 27319
rect 23845 27279 23903 27285
rect 24486 27276 24492 27328
rect 24544 27316 24550 27328
rect 25225 27319 25283 27325
rect 25225 27316 25237 27319
rect 24544 27288 25237 27316
rect 24544 27276 24550 27288
rect 25225 27285 25237 27288
rect 25271 27285 25283 27319
rect 25225 27279 25283 27285
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 3510 27121 3516 27124
rect 3467 27115 3516 27121
rect 3467 27081 3479 27115
rect 3513 27081 3516 27115
rect 3467 27075 3516 27081
rect 3510 27072 3516 27075
rect 3568 27072 3574 27124
rect 6546 27072 6552 27124
rect 6604 27072 6610 27124
rect 7834 27072 7840 27124
rect 7892 27112 7898 27124
rect 10045 27115 10103 27121
rect 7892 27084 8064 27112
rect 7892 27072 7898 27084
rect 7742 27044 7748 27056
rect 7590 27016 7748 27044
rect 7742 27004 7748 27016
rect 7800 27004 7806 27056
rect 8036 27053 8064 27084
rect 10045 27081 10057 27115
rect 10091 27112 10103 27115
rect 11974 27112 11980 27124
rect 10091 27084 11980 27112
rect 10091 27081 10103 27084
rect 10045 27075 10103 27081
rect 11974 27072 11980 27084
rect 12032 27072 12038 27124
rect 13722 27072 13728 27124
rect 13780 27112 13786 27124
rect 15749 27115 15807 27121
rect 15749 27112 15761 27115
rect 13780 27084 15761 27112
rect 13780 27072 13786 27084
rect 15749 27081 15761 27084
rect 15795 27081 15807 27115
rect 15749 27075 15807 27081
rect 18325 27115 18383 27121
rect 18325 27081 18337 27115
rect 18371 27112 18383 27115
rect 18414 27112 18420 27124
rect 18371 27084 18420 27112
rect 18371 27081 18383 27084
rect 18325 27075 18383 27081
rect 8021 27047 8079 27053
rect 8021 27013 8033 27047
rect 8067 27013 8079 27047
rect 8021 27007 8079 27013
rect 11057 27047 11115 27053
rect 11057 27013 11069 27047
rect 11103 27044 11115 27047
rect 11698 27044 11704 27056
rect 11103 27016 11704 27044
rect 11103 27013 11115 27016
rect 11057 27007 11115 27013
rect 11698 27004 11704 27016
rect 11756 27004 11762 27056
rect 13630 27044 13636 27056
rect 11992 27016 13636 27044
rect 3326 26936 3332 26988
rect 3384 26985 3390 26988
rect 3384 26979 3422 26985
rect 3410 26945 3422 26979
rect 3384 26939 3422 26945
rect 3384 26936 3390 26939
rect 3786 26936 3792 26988
rect 3844 26976 3850 26988
rect 4525 26979 4583 26985
rect 4525 26976 4537 26979
rect 3844 26948 4537 26976
rect 3844 26936 3850 26948
rect 4525 26945 4537 26948
rect 4571 26945 4583 26979
rect 4525 26939 4583 26945
rect 8297 26979 8355 26985
rect 8297 26945 8309 26979
rect 8343 26976 8355 26979
rect 8570 26976 8576 26988
rect 8343 26948 8576 26976
rect 8343 26945 8355 26948
rect 8297 26939 8355 26945
rect 8570 26936 8576 26948
rect 8628 26936 8634 26988
rect 9030 26936 9036 26988
rect 9088 26976 9094 26988
rect 9585 26979 9643 26985
rect 9585 26976 9597 26979
rect 9088 26948 9597 26976
rect 9088 26936 9094 26948
rect 9585 26945 9597 26948
rect 9631 26945 9643 26979
rect 9585 26939 9643 26945
rect 9677 26979 9735 26985
rect 9677 26945 9689 26979
rect 9723 26976 9735 26979
rect 10505 26979 10563 26985
rect 10505 26976 10517 26979
rect 9723 26948 10517 26976
rect 9723 26945 9735 26948
rect 9677 26939 9735 26945
rect 10505 26945 10517 26948
rect 10551 26945 10563 26979
rect 11882 26976 11888 26988
rect 10505 26939 10563 26945
rect 11072 26948 11888 26976
rect 3602 26868 3608 26920
rect 3660 26908 3666 26920
rect 4065 26911 4123 26917
rect 4065 26908 4077 26911
rect 3660 26880 4077 26908
rect 3660 26868 3666 26880
rect 4065 26877 4077 26880
rect 4111 26877 4123 26911
rect 4065 26871 4123 26877
rect 6178 26868 6184 26920
rect 6236 26908 6242 26920
rect 9493 26911 9551 26917
rect 6236 26880 9444 26908
rect 6236 26868 6242 26880
rect 4430 26732 4436 26784
rect 4488 26732 4494 26784
rect 9030 26732 9036 26784
rect 9088 26732 9094 26784
rect 9416 26772 9444 26880
rect 9493 26877 9505 26911
rect 9539 26877 9551 26911
rect 9600 26908 9628 26939
rect 11072 26908 11100 26948
rect 11882 26936 11888 26948
rect 11940 26936 11946 26988
rect 9600 26880 11100 26908
rect 9493 26871 9551 26877
rect 9508 26840 9536 26871
rect 11146 26868 11152 26920
rect 11204 26868 11210 26920
rect 11238 26868 11244 26920
rect 11296 26908 11302 26920
rect 11701 26911 11759 26917
rect 11701 26908 11713 26911
rect 11296 26880 11713 26908
rect 11296 26868 11302 26880
rect 11701 26877 11713 26880
rect 11747 26877 11759 26911
rect 11701 26871 11759 26877
rect 9766 26840 9772 26852
rect 9508 26812 9772 26840
rect 9766 26800 9772 26812
rect 9824 26800 9830 26852
rect 11992 26840 12020 27016
rect 13630 27004 13636 27016
rect 13688 27004 13694 27056
rect 14918 27004 14924 27056
rect 14976 27044 14982 27056
rect 15654 27044 15660 27056
rect 14976 27016 15660 27044
rect 14976 27004 14982 27016
rect 15654 27004 15660 27016
rect 15712 27004 15718 27056
rect 15764 27044 15792 27075
rect 18414 27072 18420 27084
rect 18472 27072 18478 27124
rect 20898 27112 20904 27124
rect 19306 27084 20904 27112
rect 19306 27044 19334 27084
rect 20898 27072 20904 27084
rect 20956 27072 20962 27124
rect 21358 27072 21364 27124
rect 21416 27112 21422 27124
rect 23290 27112 23296 27124
rect 21416 27084 23296 27112
rect 21416 27072 21422 27084
rect 23290 27072 23296 27084
rect 23348 27072 23354 27124
rect 23842 27072 23848 27124
rect 23900 27072 23906 27124
rect 15764 27016 19334 27044
rect 20346 27004 20352 27056
rect 20404 27044 20410 27056
rect 20404 27016 23244 27044
rect 20404 27004 20410 27016
rect 14458 26936 14464 26988
rect 14516 26976 14522 26988
rect 16301 26979 16359 26985
rect 16301 26976 16313 26979
rect 14516 26948 15148 26976
rect 14516 26936 14522 26948
rect 12434 26868 12440 26920
rect 12492 26908 12498 26920
rect 13081 26911 13139 26917
rect 13081 26908 13093 26911
rect 12492 26880 13093 26908
rect 12492 26868 12498 26880
rect 13081 26877 13093 26880
rect 13127 26877 13139 26911
rect 13081 26871 13139 26877
rect 13357 26911 13415 26917
rect 13357 26877 13369 26911
rect 13403 26908 13415 26911
rect 15010 26908 15016 26920
rect 13403 26880 15016 26908
rect 13403 26877 13415 26880
rect 13357 26871 13415 26877
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 15120 26908 15148 26948
rect 15764 26948 16313 26976
rect 15764 26908 15792 26948
rect 16301 26945 16313 26948
rect 16347 26945 16359 26979
rect 16301 26939 16359 26945
rect 17221 26979 17279 26985
rect 17221 26945 17233 26979
rect 17267 26976 17279 26979
rect 17586 26976 17592 26988
rect 17267 26948 17592 26976
rect 17267 26945 17279 26948
rect 17221 26939 17279 26945
rect 17586 26936 17592 26948
rect 17644 26936 17650 26988
rect 17770 26936 17776 26988
rect 17828 26976 17834 26988
rect 18417 26979 18475 26985
rect 18417 26976 18429 26979
rect 17828 26948 18429 26976
rect 17828 26936 17834 26948
rect 18417 26945 18429 26948
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 20438 26936 20444 26988
rect 20496 26936 20502 26988
rect 20533 26979 20591 26985
rect 20533 26945 20545 26979
rect 20579 26945 20591 26979
rect 20533 26939 20591 26945
rect 21637 26979 21695 26985
rect 21637 26945 21649 26979
rect 21683 26976 21695 26979
rect 21726 26976 21732 26988
rect 21683 26948 21732 26976
rect 21683 26945 21695 26948
rect 21637 26939 21695 26945
rect 15120 26880 15792 26908
rect 15933 26911 15991 26917
rect 15933 26877 15945 26911
rect 15979 26908 15991 26911
rect 16022 26908 16028 26920
rect 15979 26880 16028 26908
rect 15979 26877 15991 26880
rect 15933 26871 15991 26877
rect 16022 26868 16028 26880
rect 16080 26868 16086 26920
rect 16758 26868 16764 26920
rect 16816 26908 16822 26920
rect 17310 26908 17316 26920
rect 16816 26880 17316 26908
rect 16816 26868 16822 26880
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 17405 26911 17463 26917
rect 17405 26877 17417 26911
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 11072 26812 12020 26840
rect 11072 26772 11100 26812
rect 15102 26800 15108 26852
rect 15160 26840 15166 26852
rect 17420 26840 17448 26871
rect 17678 26868 17684 26920
rect 17736 26908 17742 26920
rect 18141 26911 18199 26917
rect 18141 26908 18153 26911
rect 17736 26880 18153 26908
rect 17736 26868 17742 26880
rect 18141 26877 18153 26880
rect 18187 26877 18199 26911
rect 19426 26908 19432 26920
rect 18141 26871 18199 26877
rect 18708 26880 19432 26908
rect 15160 26812 17448 26840
rect 15160 26800 15166 26812
rect 9416 26744 11100 26772
rect 11146 26732 11152 26784
rect 11204 26772 11210 26784
rect 14458 26772 14464 26784
rect 11204 26744 14464 26772
rect 11204 26732 11210 26744
rect 14458 26732 14464 26744
rect 14516 26732 14522 26784
rect 14734 26732 14740 26784
rect 14792 26772 14798 26784
rect 14829 26775 14887 26781
rect 14829 26772 14841 26775
rect 14792 26744 14841 26772
rect 14792 26732 14798 26744
rect 14829 26741 14841 26744
rect 14875 26741 14887 26775
rect 14829 26735 14887 26741
rect 15010 26732 15016 26784
rect 15068 26772 15074 26784
rect 15289 26775 15347 26781
rect 15289 26772 15301 26775
rect 15068 26744 15301 26772
rect 15068 26732 15074 26744
rect 15289 26741 15301 26744
rect 15335 26741 15347 26775
rect 15289 26735 15347 26741
rect 16850 26732 16856 26784
rect 16908 26732 16914 26784
rect 17310 26732 17316 26784
rect 17368 26772 17374 26784
rect 18708 26772 18736 26880
rect 19426 26868 19432 26880
rect 19484 26868 19490 26920
rect 19518 26868 19524 26920
rect 19576 26868 19582 26920
rect 20070 26868 20076 26920
rect 20128 26908 20134 26920
rect 20257 26911 20315 26917
rect 20257 26908 20269 26911
rect 20128 26880 20269 26908
rect 20128 26868 20134 26880
rect 20257 26877 20269 26880
rect 20303 26877 20315 26911
rect 20257 26871 20315 26877
rect 19242 26800 19248 26852
rect 19300 26840 19306 26852
rect 20548 26840 20576 26939
rect 21726 26936 21732 26948
rect 21784 26976 21790 26988
rect 22281 26979 22339 26985
rect 22281 26976 22293 26979
rect 21784 26948 22293 26976
rect 21784 26936 21790 26948
rect 22281 26945 22293 26948
rect 22327 26945 22339 26979
rect 22281 26939 22339 26945
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26976 22431 26979
rect 22738 26976 22744 26988
rect 22419 26948 22744 26976
rect 22419 26945 22431 26948
rect 22373 26939 22431 26945
rect 22738 26936 22744 26948
rect 22796 26936 22802 26988
rect 23216 26985 23244 27016
rect 23566 27004 23572 27056
rect 23624 27044 23630 27056
rect 24305 27047 24363 27053
rect 24305 27044 24317 27047
rect 23624 27016 24317 27044
rect 23624 27004 23630 27016
rect 24305 27013 24317 27016
rect 24351 27013 24363 27047
rect 24305 27007 24363 27013
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26945 23259 26979
rect 23201 26939 23259 26945
rect 23290 26936 23296 26988
rect 23348 26976 23354 26988
rect 24949 26979 25007 26985
rect 24949 26976 24961 26979
rect 23348 26948 24961 26976
rect 23348 26936 23354 26948
rect 24949 26945 24961 26948
rect 24995 26945 25007 26979
rect 24949 26939 25007 26945
rect 20806 26868 20812 26920
rect 20864 26908 20870 26920
rect 21450 26908 21456 26920
rect 20864 26880 21456 26908
rect 20864 26868 20870 26880
rect 21450 26868 21456 26880
rect 21508 26868 21514 26920
rect 22094 26868 22100 26920
rect 22152 26868 22158 26920
rect 22756 26908 22784 26936
rect 25225 26911 25283 26917
rect 25225 26908 25237 26911
rect 22756 26880 25237 26908
rect 25225 26877 25237 26880
rect 25271 26877 25283 26911
rect 25225 26871 25283 26877
rect 19300 26812 20576 26840
rect 20901 26843 20959 26849
rect 19300 26800 19306 26812
rect 20901 26809 20913 26843
rect 20947 26840 20959 26843
rect 22462 26840 22468 26852
rect 20947 26812 22468 26840
rect 20947 26809 20959 26812
rect 20901 26803 20959 26809
rect 22462 26800 22468 26812
rect 22520 26800 22526 26852
rect 23382 26840 23388 26852
rect 22572 26812 23388 26840
rect 17368 26744 18736 26772
rect 18785 26775 18843 26781
rect 17368 26732 17374 26744
rect 18785 26741 18797 26775
rect 18831 26772 18843 26775
rect 19426 26772 19432 26784
rect 18831 26744 19432 26772
rect 18831 26741 18843 26744
rect 18785 26735 18843 26741
rect 19426 26732 19432 26744
rect 19484 26732 19490 26784
rect 19702 26732 19708 26784
rect 19760 26772 19766 26784
rect 21177 26775 21235 26781
rect 21177 26772 21189 26775
rect 19760 26744 21189 26772
rect 19760 26732 19766 26744
rect 21177 26741 21189 26744
rect 21223 26772 21235 26775
rect 22572 26772 22600 26812
rect 23382 26800 23388 26812
rect 23440 26800 23446 26852
rect 21223 26744 22600 26772
rect 21223 26741 21235 26744
rect 21177 26735 21235 26741
rect 22646 26732 22652 26784
rect 22704 26772 22710 26784
rect 22741 26775 22799 26781
rect 22741 26772 22753 26775
rect 22704 26744 22753 26772
rect 22704 26732 22710 26744
rect 22741 26741 22753 26744
rect 22787 26741 22799 26775
rect 22741 26735 22799 26741
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 3786 26528 3792 26580
rect 3844 26528 3850 26580
rect 5902 26528 5908 26580
rect 5960 26568 5966 26580
rect 8573 26571 8631 26577
rect 5960 26540 8524 26568
rect 5960 26528 5966 26540
rect 8496 26500 8524 26540
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 8846 26568 8852 26580
rect 8619 26540 8852 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 8846 26528 8852 26540
rect 8904 26528 8910 26580
rect 14182 26528 14188 26580
rect 14240 26568 14246 26580
rect 14240 26540 15148 26568
rect 14240 26528 14246 26540
rect 11422 26500 11428 26512
rect 8496 26472 11428 26500
rect 11422 26460 11428 26472
rect 11480 26460 11486 26512
rect 11609 26503 11667 26509
rect 11609 26469 11621 26503
rect 11655 26500 11667 26503
rect 12986 26500 12992 26512
rect 11655 26472 12992 26500
rect 11655 26469 11667 26472
rect 11609 26463 11667 26469
rect 12986 26460 12992 26472
rect 13044 26460 13050 26512
rect 14274 26500 14280 26512
rect 13188 26472 14280 26500
rect 7098 26392 7104 26444
rect 7156 26392 7162 26444
rect 7742 26392 7748 26444
rect 7800 26432 7806 26444
rect 7800 26404 8340 26432
rect 7800 26392 7806 26404
rect 4430 26324 4436 26376
rect 4488 26364 4494 26376
rect 4893 26367 4951 26373
rect 4893 26364 4905 26367
rect 4488 26336 4905 26364
rect 4488 26324 4494 26336
rect 4893 26333 4905 26336
rect 4939 26333 4951 26367
rect 4893 26327 4951 26333
rect 6822 26324 6828 26376
rect 6880 26324 6886 26376
rect 8312 26296 8340 26404
rect 11054 26392 11060 26444
rect 11112 26392 11118 26444
rect 11146 26392 11152 26444
rect 11204 26432 11210 26444
rect 11698 26432 11704 26444
rect 11204 26404 11704 26432
rect 11204 26392 11210 26404
rect 11698 26392 11704 26404
rect 11756 26392 11762 26444
rect 13188 26441 13216 26472
rect 14274 26460 14280 26472
rect 14332 26460 14338 26512
rect 14369 26503 14427 26509
rect 14369 26469 14381 26503
rect 14415 26500 14427 26503
rect 14550 26500 14556 26512
rect 14415 26472 14556 26500
rect 14415 26469 14427 26472
rect 14369 26463 14427 26469
rect 14550 26460 14556 26472
rect 14608 26460 14614 26512
rect 15010 26500 15016 26512
rect 14660 26472 15016 26500
rect 13173 26435 13231 26441
rect 13173 26401 13185 26435
rect 13219 26401 13231 26435
rect 13173 26395 13231 26401
rect 13265 26435 13323 26441
rect 13265 26401 13277 26435
rect 13311 26432 13323 26435
rect 14660 26432 14688 26472
rect 15010 26460 15016 26472
rect 15068 26460 15074 26512
rect 15120 26500 15148 26540
rect 15470 26528 15476 26580
rect 15528 26568 15534 26580
rect 16209 26571 16267 26577
rect 16209 26568 16221 26571
rect 15528 26540 16221 26568
rect 15528 26528 15534 26540
rect 16209 26537 16221 26540
rect 16255 26537 16267 26571
rect 16209 26531 16267 26537
rect 16390 26528 16396 26580
rect 16448 26568 16454 26580
rect 16761 26571 16819 26577
rect 16761 26568 16773 26571
rect 16448 26540 16773 26568
rect 16448 26528 16454 26540
rect 16761 26537 16773 26540
rect 16807 26568 16819 26571
rect 16807 26540 19334 26568
rect 16807 26537 16819 26540
rect 16761 26531 16819 26537
rect 16666 26500 16672 26512
rect 15120 26472 16672 26500
rect 16666 26460 16672 26472
rect 16724 26500 16730 26512
rect 17310 26500 17316 26512
rect 16724 26472 17316 26500
rect 16724 26460 16730 26472
rect 17310 26460 17316 26472
rect 17368 26460 17374 26512
rect 19306 26500 19334 26540
rect 20346 26528 20352 26580
rect 20404 26528 20410 26580
rect 20622 26528 20628 26580
rect 20680 26568 20686 26580
rect 20680 26540 23060 26568
rect 20680 26528 20686 26540
rect 19702 26500 19708 26512
rect 19306 26472 19708 26500
rect 19702 26460 19708 26472
rect 19760 26500 19766 26512
rect 20806 26500 20812 26512
rect 19760 26472 20812 26500
rect 19760 26460 19766 26472
rect 20806 26460 20812 26472
rect 20864 26460 20870 26512
rect 13311 26404 14688 26432
rect 13311 26401 13323 26404
rect 13265 26395 13323 26401
rect 14826 26392 14832 26444
rect 14884 26432 14890 26444
rect 14921 26435 14979 26441
rect 14921 26432 14933 26435
rect 14884 26404 14933 26432
rect 14884 26392 14890 26404
rect 14921 26401 14933 26404
rect 14967 26401 14979 26435
rect 14921 26395 14979 26401
rect 15654 26392 15660 26444
rect 15712 26432 15718 26444
rect 16853 26435 16911 26441
rect 16853 26432 16865 26435
rect 15712 26404 16865 26432
rect 15712 26392 15718 26404
rect 16853 26401 16865 26404
rect 16899 26401 16911 26435
rect 16853 26395 16911 26401
rect 11238 26324 11244 26376
rect 11296 26324 11302 26376
rect 14734 26324 14740 26376
rect 14792 26364 14798 26376
rect 15565 26367 15623 26373
rect 15565 26364 15577 26367
rect 14792 26336 15577 26364
rect 14792 26324 14798 26336
rect 15565 26333 15577 26336
rect 15611 26333 15623 26367
rect 16868 26364 16896 26395
rect 17586 26392 17592 26444
rect 17644 26432 17650 26444
rect 17773 26435 17831 26441
rect 17773 26432 17785 26435
rect 17644 26404 17785 26432
rect 17644 26392 17650 26404
rect 17773 26401 17785 26404
rect 17819 26432 17831 26435
rect 21726 26432 21732 26444
rect 17819 26404 21732 26432
rect 17819 26401 17831 26404
rect 17773 26395 17831 26401
rect 21726 26392 21732 26404
rect 21784 26392 21790 26444
rect 23032 26441 23060 26540
rect 23017 26435 23075 26441
rect 23017 26401 23029 26435
rect 23063 26401 23075 26435
rect 23017 26395 23075 26401
rect 23106 26392 23112 26444
rect 23164 26392 23170 26444
rect 19242 26364 19248 26376
rect 16868 26336 19248 26364
rect 15565 26327 15623 26333
rect 19242 26324 19248 26336
rect 19300 26364 19306 26376
rect 19981 26367 20039 26373
rect 19981 26364 19993 26367
rect 19300 26336 19993 26364
rect 19300 26324 19306 26336
rect 19981 26333 19993 26336
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26364 22155 26367
rect 22186 26364 22192 26376
rect 22143 26336 22192 26364
rect 22143 26333 22155 26336
rect 22097 26327 22155 26333
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 22554 26324 22560 26376
rect 22612 26324 22618 26376
rect 22738 26324 22744 26376
rect 22796 26364 22802 26376
rect 22925 26367 22983 26373
rect 22925 26364 22937 26367
rect 22796 26336 22937 26364
rect 22796 26324 22802 26336
rect 22925 26333 22937 26336
rect 22971 26333 22983 26367
rect 22925 26327 22983 26333
rect 23658 26324 23664 26376
rect 23716 26364 23722 26376
rect 23937 26367 23995 26373
rect 23937 26364 23949 26367
rect 23716 26336 23949 26364
rect 23716 26324 23722 26336
rect 23937 26333 23949 26336
rect 23983 26333 23995 26367
rect 23937 26327 23995 26333
rect 24026 26324 24032 26376
rect 24084 26364 24090 26376
rect 24765 26367 24823 26373
rect 24765 26364 24777 26367
rect 24084 26336 24777 26364
rect 24084 26324 24090 26336
rect 24765 26333 24777 26336
rect 24811 26333 24823 26367
rect 24765 26327 24823 26333
rect 9214 26296 9220 26308
rect 8312 26282 9220 26296
rect 8326 26268 9220 26282
rect 9214 26256 9220 26268
rect 9272 26256 9278 26308
rect 10042 26256 10048 26308
rect 10100 26296 10106 26308
rect 10137 26299 10195 26305
rect 10137 26296 10149 26299
rect 10100 26268 10149 26296
rect 10100 26256 10106 26268
rect 10137 26265 10149 26268
rect 10183 26265 10195 26299
rect 10137 26259 10195 26265
rect 10321 26299 10379 26305
rect 10321 26265 10333 26299
rect 10367 26296 10379 26299
rect 11606 26296 11612 26308
rect 10367 26268 11612 26296
rect 10367 26265 10379 26268
rect 10321 26259 10379 26265
rect 11606 26256 11612 26268
rect 11664 26256 11670 26308
rect 14829 26299 14887 26305
rect 14829 26265 14841 26299
rect 14875 26296 14887 26299
rect 14918 26296 14924 26308
rect 14875 26268 14924 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 14918 26256 14924 26268
rect 14976 26256 14982 26308
rect 16758 26256 16764 26308
rect 16816 26296 16822 26308
rect 17037 26299 17095 26305
rect 17037 26296 17049 26299
rect 16816 26268 17049 26296
rect 16816 26256 16822 26268
rect 17037 26265 17049 26268
rect 17083 26265 17095 26299
rect 21821 26299 21879 26305
rect 21390 26268 21772 26296
rect 17037 26259 17095 26265
rect 5534 26188 5540 26240
rect 5592 26188 5598 26240
rect 13354 26188 13360 26240
rect 13412 26188 13418 26240
rect 13725 26231 13783 26237
rect 13725 26197 13737 26231
rect 13771 26228 13783 26231
rect 14642 26228 14648 26240
rect 13771 26200 14648 26228
rect 13771 26197 13783 26200
rect 13725 26191 13783 26197
rect 14642 26188 14648 26200
rect 14700 26188 14706 26240
rect 14737 26231 14795 26237
rect 14737 26197 14749 26231
rect 14783 26228 14795 26231
rect 15194 26228 15200 26240
rect 14783 26200 15200 26228
rect 14783 26197 14795 26200
rect 14737 26191 14795 26197
rect 15194 26188 15200 26200
rect 15252 26188 15258 26240
rect 16577 26231 16635 26237
rect 16577 26197 16589 26231
rect 16623 26228 16635 26231
rect 17126 26228 17132 26240
rect 16623 26200 17132 26228
rect 16623 26197 16635 26200
rect 16577 26191 16635 26197
rect 17126 26188 17132 26200
rect 17184 26188 17190 26240
rect 17770 26188 17776 26240
rect 17828 26228 17834 26240
rect 17865 26231 17923 26237
rect 17865 26228 17877 26231
rect 17828 26200 17877 26228
rect 17828 26188 17834 26200
rect 17865 26197 17877 26200
rect 17911 26197 17923 26231
rect 21744 26228 21772 26268
rect 21821 26265 21833 26299
rect 21867 26296 21879 26299
rect 22370 26296 22376 26308
rect 21867 26268 22376 26296
rect 21867 26265 21879 26268
rect 21821 26259 21879 26265
rect 22370 26256 22376 26268
rect 22428 26256 22434 26308
rect 22572 26296 22600 26324
rect 23382 26296 23388 26308
rect 22480 26268 23388 26296
rect 22480 26228 22508 26268
rect 23382 26256 23388 26268
rect 23440 26256 23446 26308
rect 23750 26256 23756 26308
rect 23808 26256 23814 26308
rect 24118 26256 24124 26308
rect 24176 26296 24182 26308
rect 24581 26299 24639 26305
rect 24581 26296 24593 26299
rect 24176 26268 24593 26296
rect 24176 26256 24182 26268
rect 24581 26265 24593 26268
rect 24627 26265 24639 26299
rect 24581 26259 24639 26265
rect 21744 26200 22508 26228
rect 17865 26191 17923 26197
rect 22554 26188 22560 26240
rect 22612 26188 22618 26240
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 3283 26027 3341 26033
rect 3283 25993 3295 26027
rect 3329 26024 3341 26027
rect 3418 26024 3424 26036
rect 3329 25996 3424 26024
rect 3329 25993 3341 25996
rect 3283 25987 3341 25993
rect 3418 25984 3424 25996
rect 3476 25984 3482 26036
rect 5534 26024 5540 26036
rect 5276 25996 5540 26024
rect 5276 25965 5304 25996
rect 5534 25984 5540 25996
rect 5592 25984 5598 26036
rect 12986 25984 12992 26036
rect 13044 25984 13050 26036
rect 13262 25984 13268 26036
rect 13320 26024 13326 26036
rect 14553 26027 14611 26033
rect 14553 26024 14565 26027
rect 13320 25996 14565 26024
rect 13320 25984 13326 25996
rect 14553 25993 14565 25996
rect 14599 26024 14611 26027
rect 15930 26024 15936 26036
rect 14599 25996 15936 26024
rect 14599 25993 14611 25996
rect 14553 25987 14611 25993
rect 15930 25984 15936 25996
rect 15988 25984 15994 26036
rect 16574 26024 16580 26036
rect 16040 25996 16580 26024
rect 5261 25959 5319 25965
rect 5261 25925 5273 25959
rect 5307 25925 5319 25959
rect 6822 25956 6828 25968
rect 5261 25919 5319 25925
rect 5552 25928 6828 25956
rect 3212 25891 3270 25897
rect 3212 25857 3224 25891
rect 3258 25888 3270 25891
rect 3418 25888 3424 25900
rect 3258 25860 3424 25888
rect 3258 25857 3270 25860
rect 3212 25851 3270 25857
rect 3418 25848 3424 25860
rect 3476 25848 3482 25900
rect 5552 25897 5580 25928
rect 6822 25916 6828 25928
rect 6880 25956 6886 25968
rect 8570 25956 8576 25968
rect 6880 25928 8576 25956
rect 6880 25916 6886 25928
rect 8220 25897 8248 25928
rect 8570 25916 8576 25928
rect 8628 25916 8634 25968
rect 9214 25916 9220 25968
rect 9272 25916 9278 25968
rect 12897 25959 12955 25965
rect 12897 25925 12909 25959
rect 12943 25956 12955 25959
rect 13538 25956 13544 25968
rect 12943 25928 13544 25956
rect 12943 25925 12955 25928
rect 12897 25919 12955 25925
rect 13538 25916 13544 25928
rect 13596 25916 13602 25968
rect 16040 25956 16068 25996
rect 16574 25984 16580 25996
rect 16632 26024 16638 26036
rect 16669 26027 16727 26033
rect 16669 26024 16681 26027
rect 16632 25996 16681 26024
rect 16632 25984 16638 25996
rect 16669 25993 16681 25996
rect 16715 25993 16727 26027
rect 16669 25987 16727 25993
rect 18322 25984 18328 26036
rect 18380 25984 18386 26036
rect 19058 25984 19064 26036
rect 19116 26024 19122 26036
rect 19116 25996 19288 26024
rect 19116 25984 19122 25996
rect 15594 25928 16068 25956
rect 16114 25916 16120 25968
rect 16172 25956 16178 25968
rect 18233 25959 18291 25965
rect 16172 25928 16344 25956
rect 16172 25916 16178 25928
rect 5537 25891 5595 25897
rect 4172 25820 4200 25874
rect 5537 25857 5549 25891
rect 5583 25857 5595 25891
rect 5537 25851 5595 25857
rect 8205 25891 8263 25897
rect 8205 25857 8217 25891
rect 8251 25857 8263 25891
rect 11057 25891 11115 25897
rect 11057 25888 11069 25891
rect 8205 25851 8263 25857
rect 9968 25860 11069 25888
rect 4172 25792 5856 25820
rect 5828 25696 5856 25792
rect 7742 25780 7748 25832
rect 7800 25780 7806 25832
rect 8481 25823 8539 25829
rect 8481 25789 8493 25823
rect 8527 25820 8539 25823
rect 8846 25820 8852 25832
rect 8527 25792 8852 25820
rect 8527 25789 8539 25792
rect 8481 25783 8539 25789
rect 8846 25780 8852 25792
rect 8904 25780 8910 25832
rect 9968 25829 9996 25860
rect 11057 25857 11069 25860
rect 11103 25888 11115 25891
rect 11882 25888 11888 25900
rect 11103 25860 11888 25888
rect 11103 25857 11115 25860
rect 11057 25851 11115 25857
rect 11882 25848 11888 25860
rect 11940 25848 11946 25900
rect 12342 25848 12348 25900
rect 12400 25888 12406 25900
rect 16316 25897 16344 25928
rect 18233 25925 18245 25959
rect 18279 25956 18291 25959
rect 19150 25956 19156 25968
rect 18279 25928 19156 25956
rect 18279 25925 18291 25928
rect 18233 25919 18291 25925
rect 19150 25916 19156 25928
rect 19208 25916 19214 25968
rect 19260 25956 19288 25996
rect 19518 25984 19524 26036
rect 19576 26024 19582 26036
rect 19613 26027 19671 26033
rect 19613 26024 19625 26027
rect 19576 25996 19625 26024
rect 19576 25984 19582 25996
rect 19613 25993 19625 25996
rect 19659 25993 19671 26027
rect 19613 25987 19671 25993
rect 21913 26027 21971 26033
rect 21913 25993 21925 26027
rect 21959 26024 21971 26027
rect 23198 26024 23204 26036
rect 21959 25996 23204 26024
rect 21959 25993 21971 25996
rect 21913 25987 21971 25993
rect 20438 25956 20444 25968
rect 19260 25928 20444 25956
rect 20438 25916 20444 25928
rect 20496 25916 20502 25968
rect 16301 25891 16359 25897
rect 12400 25860 12756 25888
rect 12400 25848 12406 25860
rect 9953 25823 10011 25829
rect 9953 25789 9965 25823
rect 9999 25789 10011 25823
rect 9953 25783 10011 25789
rect 12161 25823 12219 25829
rect 12161 25789 12173 25823
rect 12207 25820 12219 25823
rect 12526 25820 12532 25832
rect 12207 25792 12532 25820
rect 12207 25789 12219 25792
rect 12161 25783 12219 25789
rect 12526 25780 12532 25792
rect 12584 25780 12590 25832
rect 12728 25829 12756 25860
rect 16301 25857 16313 25891
rect 16347 25888 16359 25891
rect 17126 25888 17132 25900
rect 16347 25860 17132 25888
rect 16347 25857 16359 25860
rect 16301 25851 16359 25857
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19521 25891 19579 25897
rect 19521 25888 19533 25891
rect 19484 25860 19533 25888
rect 19484 25848 19490 25860
rect 19521 25857 19533 25860
rect 19567 25857 19579 25891
rect 19521 25851 19579 25857
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25888 21511 25891
rect 21928 25888 21956 25987
rect 23198 25984 23204 25996
rect 23256 25984 23262 26036
rect 22278 25916 22284 25968
rect 22336 25956 22342 25968
rect 22465 25959 22523 25965
rect 22465 25956 22477 25959
rect 22336 25928 22477 25956
rect 22336 25916 22342 25928
rect 22465 25925 22477 25928
rect 22511 25925 22523 25959
rect 22465 25919 22523 25925
rect 24486 25916 24492 25968
rect 24544 25916 24550 25968
rect 23198 25888 23204 25900
rect 21499 25860 21956 25888
rect 23032 25860 23204 25888
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 12713 25823 12771 25829
rect 12713 25789 12725 25823
rect 12759 25789 12771 25823
rect 12713 25783 12771 25789
rect 16022 25780 16028 25832
rect 16080 25780 16086 25832
rect 18509 25823 18567 25829
rect 18509 25789 18521 25823
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 9674 25712 9680 25764
rect 9732 25752 9738 25764
rect 10413 25755 10471 25761
rect 10413 25752 10425 25755
rect 9732 25724 10425 25752
rect 9732 25712 9738 25724
rect 10413 25721 10425 25724
rect 10459 25721 10471 25755
rect 10413 25715 10471 25721
rect 3789 25687 3847 25693
rect 3789 25653 3801 25687
rect 3835 25684 3847 25687
rect 4154 25684 4160 25696
rect 3835 25656 4160 25684
rect 3835 25653 3847 25656
rect 3789 25647 3847 25653
rect 4154 25644 4160 25656
rect 4212 25644 4218 25696
rect 5810 25644 5816 25696
rect 5868 25644 5874 25696
rect 12802 25644 12808 25696
rect 12860 25684 12866 25696
rect 13262 25684 13268 25696
rect 12860 25656 13268 25684
rect 12860 25644 12866 25656
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 13357 25687 13415 25693
rect 13357 25653 13369 25687
rect 13403 25684 13415 25687
rect 13630 25684 13636 25696
rect 13403 25656 13636 25684
rect 13403 25653 13415 25656
rect 13357 25647 13415 25653
rect 13630 25644 13636 25656
rect 13688 25644 13694 25696
rect 17865 25687 17923 25693
rect 17865 25653 17877 25687
rect 17911 25684 17923 25687
rect 18322 25684 18328 25696
rect 17911 25656 18328 25684
rect 17911 25653 17923 25656
rect 17865 25647 17923 25653
rect 18322 25644 18328 25656
rect 18380 25644 18386 25696
rect 18524 25684 18552 25783
rect 19334 25780 19340 25832
rect 19392 25780 19398 25832
rect 22830 25780 22836 25832
rect 22888 25820 22894 25832
rect 23032 25829 23060 25860
rect 23198 25848 23204 25860
rect 23256 25848 23262 25900
rect 23382 25848 23388 25900
rect 23440 25848 23446 25900
rect 23017 25823 23075 25829
rect 23017 25820 23029 25823
rect 22888 25792 23029 25820
rect 22888 25780 22894 25792
rect 23017 25789 23029 25792
rect 23063 25789 23075 25823
rect 23017 25783 23075 25789
rect 24762 25780 24768 25832
rect 24820 25780 24826 25832
rect 18690 25712 18696 25764
rect 18748 25752 18754 25764
rect 20898 25752 20904 25764
rect 18748 25724 20904 25752
rect 18748 25712 18754 25724
rect 20898 25712 20904 25724
rect 20956 25752 20962 25764
rect 21269 25755 21327 25761
rect 21269 25752 21281 25755
rect 20956 25724 21281 25752
rect 20956 25712 20962 25724
rect 21269 25721 21281 25724
rect 21315 25721 21327 25755
rect 21269 25715 21327 25721
rect 19426 25684 19432 25696
rect 18524 25656 19432 25684
rect 19426 25644 19432 25656
rect 19484 25644 19490 25696
rect 19518 25644 19524 25696
rect 19576 25684 19582 25696
rect 19702 25684 19708 25696
rect 19576 25656 19708 25684
rect 19576 25644 19582 25656
rect 19702 25644 19708 25656
rect 19760 25644 19766 25696
rect 19886 25644 19892 25696
rect 19944 25684 19950 25696
rect 19981 25687 20039 25693
rect 19981 25684 19993 25687
rect 19944 25656 19993 25684
rect 19944 25644 19950 25656
rect 19981 25653 19993 25656
rect 20027 25653 20039 25687
rect 19981 25647 20039 25653
rect 22370 25644 22376 25696
rect 22428 25644 22434 25696
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 3329 25483 3387 25489
rect 3329 25449 3341 25483
rect 3375 25480 3387 25483
rect 4154 25480 4160 25492
rect 3375 25452 4160 25480
rect 3375 25449 3387 25452
rect 3329 25443 3387 25449
rect 4154 25440 4160 25452
rect 4212 25440 4218 25492
rect 4430 25440 4436 25492
rect 4488 25440 4494 25492
rect 11422 25440 11428 25492
rect 11480 25480 11486 25492
rect 11793 25483 11851 25489
rect 11793 25480 11805 25483
rect 11480 25452 11805 25480
rect 11480 25440 11486 25452
rect 11793 25449 11805 25452
rect 11839 25449 11851 25483
rect 11793 25443 11851 25449
rect 12897 25483 12955 25489
rect 12897 25449 12909 25483
rect 12943 25480 12955 25483
rect 13354 25480 13360 25492
rect 12943 25452 13360 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 13354 25440 13360 25452
rect 13412 25440 13418 25492
rect 15749 25483 15807 25489
rect 15749 25449 15761 25483
rect 15795 25480 15807 25483
rect 16022 25480 16028 25492
rect 15795 25452 16028 25480
rect 15795 25449 15807 25452
rect 15749 25443 15807 25449
rect 16022 25440 16028 25452
rect 16080 25440 16086 25492
rect 9861 25415 9919 25421
rect 9861 25381 9873 25415
rect 9907 25412 9919 25415
rect 12066 25412 12072 25424
rect 9907 25384 12072 25412
rect 9907 25381 9919 25384
rect 9861 25375 9919 25381
rect 12066 25372 12072 25384
rect 12124 25372 12130 25424
rect 14366 25372 14372 25424
rect 14424 25412 14430 25424
rect 18233 25415 18291 25421
rect 14424 25384 16528 25412
rect 14424 25372 14430 25384
rect 6181 25347 6239 25353
rect 6181 25313 6193 25347
rect 6227 25344 6239 25347
rect 6822 25344 6828 25356
rect 6227 25316 6828 25344
rect 6227 25313 6239 25316
rect 6181 25307 6239 25313
rect 6822 25304 6828 25316
rect 6880 25344 6886 25356
rect 7098 25344 7104 25356
rect 6880 25316 7104 25344
rect 6880 25304 6886 25316
rect 7098 25304 7104 25316
rect 7156 25304 7162 25356
rect 7834 25304 7840 25356
rect 7892 25344 7898 25356
rect 7929 25347 7987 25353
rect 7929 25344 7941 25347
rect 7892 25316 7941 25344
rect 7892 25304 7898 25316
rect 7929 25313 7941 25316
rect 7975 25313 7987 25347
rect 7929 25307 7987 25313
rect 8846 25304 8852 25356
rect 8904 25344 8910 25356
rect 9217 25347 9275 25353
rect 9217 25344 9229 25347
rect 8904 25316 9229 25344
rect 8904 25304 8910 25316
rect 9217 25313 9229 25316
rect 9263 25313 9275 25347
rect 9217 25307 9275 25313
rect 9490 25304 9496 25356
rect 9548 25344 9554 25356
rect 10689 25347 10747 25353
rect 10689 25344 10701 25347
rect 9548 25316 10701 25344
rect 9548 25304 9554 25316
rect 10689 25313 10701 25316
rect 10735 25313 10747 25347
rect 10689 25307 10747 25313
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 12345 25347 12403 25353
rect 12345 25313 12357 25347
rect 12391 25344 12403 25347
rect 12802 25344 12808 25356
rect 12391 25316 12808 25344
rect 12391 25313 12403 25316
rect 12345 25307 12403 25313
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 14553 25347 14611 25353
rect 14553 25313 14565 25347
rect 14599 25344 14611 25347
rect 14734 25344 14740 25356
rect 14599 25316 14740 25344
rect 14599 25313 14611 25316
rect 14553 25307 14611 25313
rect 14734 25304 14740 25316
rect 14792 25304 14798 25356
rect 2593 25279 2651 25285
rect 2593 25245 2605 25279
rect 2639 25276 2651 25279
rect 3421 25279 3479 25285
rect 3421 25276 3433 25279
rect 2639 25248 3433 25276
rect 2639 25245 2651 25248
rect 2593 25239 2651 25245
rect 3421 25245 3433 25248
rect 3467 25276 3479 25279
rect 3786 25276 3792 25288
rect 3467 25248 3792 25276
rect 3467 25245 3479 25248
rect 3421 25239 3479 25245
rect 3786 25236 3792 25248
rect 3844 25276 3850 25288
rect 4430 25276 4436 25288
rect 3844 25248 4436 25276
rect 3844 25236 3850 25248
rect 4430 25236 4436 25248
rect 4488 25236 4494 25288
rect 6270 25236 6276 25288
rect 6328 25276 6334 25288
rect 7285 25279 7343 25285
rect 7285 25276 7297 25279
rect 6328 25248 7297 25276
rect 6328 25236 6334 25248
rect 7285 25245 7297 25248
rect 7331 25245 7343 25279
rect 7285 25239 7343 25245
rect 7742 25236 7748 25288
rect 7800 25276 7806 25288
rect 8205 25279 8263 25285
rect 8205 25276 8217 25279
rect 7800 25248 8217 25276
rect 7800 25236 7806 25248
rect 8205 25245 8217 25248
rect 8251 25245 8263 25279
rect 8205 25239 8263 25245
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 9401 25279 9459 25285
rect 9401 25276 9413 25279
rect 8352 25248 9413 25276
rect 8352 25236 8358 25248
rect 9401 25245 9413 25248
rect 9447 25276 9459 25279
rect 10226 25276 10232 25288
rect 9447 25248 10232 25276
rect 9447 25245 9459 25248
rect 9401 25239 9459 25245
rect 10226 25236 10232 25248
rect 10284 25236 10290 25288
rect 12526 25236 12532 25288
rect 12584 25236 12590 25288
rect 14642 25236 14648 25288
rect 14700 25276 14706 25288
rect 14829 25279 14887 25285
rect 14829 25276 14841 25279
rect 14700 25248 14841 25276
rect 14700 25236 14706 25248
rect 14829 25245 14841 25248
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 16022 25236 16028 25288
rect 16080 25276 16086 25288
rect 16393 25279 16451 25285
rect 16393 25276 16405 25279
rect 16080 25248 16405 25276
rect 16080 25236 16086 25248
rect 16393 25245 16405 25248
rect 16439 25245 16451 25279
rect 16500 25276 16528 25384
rect 18233 25381 18245 25415
rect 18279 25412 18291 25415
rect 21910 25412 21916 25424
rect 18279 25384 21916 25412
rect 18279 25381 18291 25384
rect 18233 25375 18291 25381
rect 21910 25372 21916 25384
rect 21968 25372 21974 25424
rect 17218 25304 17224 25356
rect 17276 25344 17282 25356
rect 17313 25347 17371 25353
rect 17313 25344 17325 25347
rect 17276 25316 17325 25344
rect 17276 25304 17282 25316
rect 17313 25313 17325 25316
rect 17359 25313 17371 25347
rect 17313 25307 17371 25313
rect 17497 25347 17555 25353
rect 17497 25313 17509 25347
rect 17543 25344 17555 25347
rect 18690 25344 18696 25356
rect 17543 25316 18696 25344
rect 17543 25313 17555 25316
rect 17497 25307 17555 25313
rect 18690 25304 18696 25316
rect 18748 25344 18754 25356
rect 18874 25344 18880 25356
rect 18748 25316 18880 25344
rect 18748 25304 18754 25316
rect 18874 25304 18880 25316
rect 18932 25304 18938 25356
rect 20073 25347 20131 25353
rect 20073 25313 20085 25347
rect 20119 25344 20131 25347
rect 20809 25347 20867 25353
rect 20119 25316 20668 25344
rect 20119 25313 20131 25316
rect 20073 25307 20131 25313
rect 18049 25279 18107 25285
rect 18049 25276 18061 25279
rect 16500 25248 18061 25276
rect 16393 25239 16451 25245
rect 18049 25245 18061 25248
rect 18095 25245 18107 25279
rect 18049 25239 18107 25245
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 20162 25276 20168 25288
rect 19935 25248 20168 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 20162 25236 20168 25248
rect 20220 25236 20226 25288
rect 20640 25276 20668 25316
rect 20809 25313 20821 25347
rect 20855 25344 20867 25347
rect 21266 25344 21272 25356
rect 20855 25316 21272 25344
rect 20855 25313 20867 25316
rect 20809 25307 20867 25313
rect 21266 25304 21272 25316
rect 21324 25344 21330 25356
rect 22002 25344 22008 25356
rect 21324 25316 22008 25344
rect 21324 25304 21330 25316
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 22462 25304 22468 25356
rect 22520 25344 22526 25356
rect 22649 25347 22707 25353
rect 22649 25344 22661 25347
rect 22520 25316 22661 25344
rect 22520 25304 22526 25316
rect 22649 25313 22661 25316
rect 22695 25313 22707 25347
rect 22649 25307 22707 25313
rect 22833 25347 22891 25353
rect 22833 25313 22845 25347
rect 22879 25344 22891 25347
rect 24302 25344 24308 25356
rect 22879 25316 24308 25344
rect 22879 25313 22891 25316
rect 22833 25307 22891 25313
rect 24302 25304 24308 25316
rect 24360 25304 24366 25356
rect 21634 25276 21640 25288
rect 20640 25248 21640 25276
rect 21634 25236 21640 25248
rect 21692 25236 21698 25288
rect 22557 25279 22615 25285
rect 22557 25245 22569 25279
rect 22603 25276 22615 25279
rect 23474 25276 23480 25288
rect 22603 25248 23480 25276
rect 22603 25245 22615 25248
rect 22557 25239 22615 25245
rect 23474 25236 23480 25248
rect 23532 25236 23538 25288
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25276 23903 25279
rect 23934 25276 23940 25288
rect 23891 25248 23940 25276
rect 23891 25245 23903 25248
rect 23845 25239 23903 25245
rect 23934 25236 23940 25248
rect 23992 25236 23998 25288
rect 24854 25236 24860 25288
rect 24912 25236 24918 25288
rect 5810 25208 5816 25220
rect 5474 25180 5816 25208
rect 5810 25168 5816 25180
rect 5868 25168 5874 25220
rect 5905 25211 5963 25217
rect 5905 25177 5917 25211
rect 5951 25208 5963 25211
rect 6641 25211 6699 25217
rect 6641 25208 6653 25211
rect 5951 25180 6653 25208
rect 5951 25177 5963 25180
rect 5905 25171 5963 25177
rect 6641 25177 6653 25180
rect 6687 25177 6699 25211
rect 6641 25171 6699 25177
rect 7650 25168 7656 25220
rect 7708 25208 7714 25220
rect 8113 25211 8171 25217
rect 8113 25208 8125 25211
rect 7708 25180 8125 25208
rect 7708 25168 7714 25180
rect 8113 25177 8125 25180
rect 8159 25177 8171 25211
rect 10965 25211 11023 25217
rect 10965 25208 10977 25211
rect 8113 25171 8171 25177
rect 8588 25180 10977 25208
rect 2961 25143 3019 25149
rect 2961 25109 2973 25143
rect 3007 25140 3019 25143
rect 3326 25140 3332 25152
rect 3007 25112 3332 25140
rect 3007 25109 3019 25112
rect 2961 25103 3019 25109
rect 3326 25100 3332 25112
rect 3384 25100 3390 25152
rect 5828 25140 5856 25168
rect 6362 25140 6368 25152
rect 5828 25112 6368 25140
rect 6362 25100 6368 25112
rect 6420 25100 6426 25152
rect 8588 25149 8616 25180
rect 10965 25177 10977 25180
rect 11011 25177 11023 25211
rect 14090 25208 14096 25220
rect 10965 25171 11023 25177
rect 11348 25180 14096 25208
rect 8573 25143 8631 25149
rect 8573 25109 8585 25143
rect 8619 25109 8631 25143
rect 8573 25103 8631 25109
rect 9490 25100 9496 25152
rect 9548 25100 9554 25152
rect 10226 25100 10232 25152
rect 10284 25100 10290 25152
rect 11348 25149 11376 25180
rect 14090 25168 14096 25180
rect 14148 25168 14154 25220
rect 14737 25211 14795 25217
rect 14737 25177 14749 25211
rect 14783 25208 14795 25211
rect 15378 25208 15384 25220
rect 14783 25180 15384 25208
rect 14783 25177 14795 25180
rect 14737 25171 14795 25177
rect 15378 25168 15384 25180
rect 15436 25168 15442 25220
rect 16758 25168 16764 25220
rect 16816 25208 16822 25220
rect 17221 25211 17279 25217
rect 17221 25208 17233 25211
rect 16816 25180 17233 25208
rect 16816 25168 16822 25180
rect 17221 25177 17233 25180
rect 17267 25208 17279 25211
rect 17770 25208 17776 25220
rect 17267 25180 17776 25208
rect 17267 25177 17279 25180
rect 17221 25171 17279 25177
rect 17770 25168 17776 25180
rect 17828 25168 17834 25220
rect 19797 25211 19855 25217
rect 19797 25177 19809 25211
rect 19843 25208 19855 25211
rect 20714 25208 20720 25220
rect 19843 25180 20720 25208
rect 19843 25177 19855 25180
rect 19797 25171 19855 25177
rect 20714 25168 20720 25180
rect 20772 25168 20778 25220
rect 20898 25168 20904 25220
rect 20956 25168 20962 25220
rect 22094 25168 22100 25220
rect 22152 25208 22158 25220
rect 22462 25208 22468 25220
rect 22152 25180 22468 25208
rect 22152 25168 22158 25180
rect 22462 25168 22468 25180
rect 22520 25168 22526 25220
rect 11333 25143 11391 25149
rect 11333 25109 11345 25143
rect 11379 25109 11391 25143
rect 11333 25103 11391 25109
rect 11422 25100 11428 25152
rect 11480 25140 11486 25152
rect 12437 25143 12495 25149
rect 12437 25140 12449 25143
rect 11480 25112 12449 25140
rect 11480 25100 11486 25112
rect 12437 25109 12449 25112
rect 12483 25140 12495 25143
rect 13722 25140 13728 25152
rect 12483 25112 13728 25140
rect 12483 25109 12495 25112
rect 12437 25103 12495 25109
rect 13722 25100 13728 25112
rect 13780 25100 13786 25152
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 15470 25140 15476 25152
rect 15243 25112 15476 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 15470 25100 15476 25112
rect 15528 25100 15534 25152
rect 15838 25100 15844 25152
rect 15896 25140 15902 25152
rect 16853 25143 16911 25149
rect 16853 25140 16865 25143
rect 15896 25112 16865 25140
rect 15896 25100 15902 25112
rect 16853 25109 16865 25112
rect 16899 25109 16911 25143
rect 16853 25103 16911 25109
rect 19429 25143 19487 25149
rect 19429 25109 19441 25143
rect 19475 25140 19487 25143
rect 19702 25140 19708 25152
rect 19475 25112 19708 25140
rect 19475 25109 19487 25112
rect 19429 25103 19487 25109
rect 19702 25100 19708 25112
rect 19760 25100 19766 25152
rect 20438 25100 20444 25152
rect 20496 25140 20502 25152
rect 20993 25143 21051 25149
rect 20993 25140 21005 25143
rect 20496 25112 21005 25140
rect 20496 25100 20502 25112
rect 20993 25109 21005 25112
rect 21039 25109 21051 25143
rect 20993 25103 21051 25109
rect 21361 25143 21419 25149
rect 21361 25109 21373 25143
rect 21407 25140 21419 25143
rect 21726 25140 21732 25152
rect 21407 25112 21732 25140
rect 21407 25109 21419 25112
rect 21361 25103 21419 25109
rect 21726 25100 21732 25112
rect 21784 25100 21790 25152
rect 22189 25143 22247 25149
rect 22189 25109 22201 25143
rect 22235 25140 22247 25143
rect 22278 25140 22284 25152
rect 22235 25112 22284 25140
rect 22235 25109 22247 25112
rect 22189 25103 22247 25109
rect 22278 25100 22284 25112
rect 22336 25100 22342 25152
rect 23934 25100 23940 25152
rect 23992 25100 23998 25152
rect 24026 25100 24032 25152
rect 24084 25140 24090 25152
rect 24673 25143 24731 25149
rect 24673 25140 24685 25143
rect 24084 25112 24685 25140
rect 24084 25100 24090 25112
rect 24673 25109 24685 25112
rect 24719 25109 24731 25143
rect 24673 25103 24731 25109
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 7190 24896 7196 24948
rect 7248 24936 7254 24948
rect 7650 24936 7656 24948
rect 7248 24908 7656 24936
rect 7248 24896 7254 24908
rect 7650 24896 7656 24908
rect 7708 24896 7714 24948
rect 8941 24939 8999 24945
rect 8941 24905 8953 24939
rect 8987 24936 8999 24939
rect 9490 24936 9496 24948
rect 8987 24908 9496 24936
rect 8987 24905 8999 24908
rect 8941 24899 8999 24905
rect 9490 24896 9496 24908
rect 9548 24896 9554 24948
rect 16758 24896 16764 24948
rect 16816 24896 16822 24948
rect 19886 24896 19892 24948
rect 19944 24896 19950 24948
rect 21085 24939 21143 24945
rect 21085 24905 21097 24939
rect 21131 24936 21143 24939
rect 22278 24936 22284 24948
rect 21131 24908 22284 24936
rect 21131 24905 21143 24908
rect 21085 24899 21143 24905
rect 22278 24896 22284 24908
rect 22336 24896 22342 24948
rect 9674 24828 9680 24880
rect 9732 24828 9738 24880
rect 13096 24840 13768 24868
rect 4341 24803 4399 24809
rect 4341 24769 4353 24803
rect 4387 24800 4399 24803
rect 6546 24800 6552 24812
rect 4387 24772 6552 24800
rect 4387 24769 4399 24772
rect 4341 24763 4399 24769
rect 6546 24760 6552 24772
rect 6604 24760 6610 24812
rect 9306 24760 9312 24812
rect 9364 24800 9370 24812
rect 9401 24803 9459 24809
rect 9401 24800 9413 24803
rect 9364 24772 9413 24800
rect 9364 24760 9370 24772
rect 9401 24769 9413 24772
rect 9447 24769 9459 24803
rect 11974 24800 11980 24812
rect 10810 24786 11980 24800
rect 9401 24763 9459 24769
rect 10796 24772 11980 24786
rect 2866 24692 2872 24744
rect 2924 24692 2930 24744
rect 3326 24692 3332 24744
rect 3384 24732 3390 24744
rect 3513 24735 3571 24741
rect 3513 24732 3525 24735
rect 3384 24704 3525 24732
rect 3384 24692 3390 24704
rect 3513 24701 3525 24704
rect 3559 24701 3571 24735
rect 3513 24695 3571 24701
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24732 3755 24735
rect 3743 24704 4384 24732
rect 3743 24701 3755 24704
rect 3697 24695 3755 24701
rect 4356 24676 4384 24704
rect 9214 24692 9220 24744
rect 9272 24732 9278 24744
rect 10796 24732 10824 24772
rect 11974 24760 11980 24772
rect 12032 24760 12038 24812
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24800 12403 24803
rect 12391 24772 12425 24800
rect 12391 24769 12403 24772
rect 12345 24763 12403 24769
rect 12360 24732 12388 24763
rect 13096 24732 13124 24840
rect 13173 24803 13231 24809
rect 13173 24769 13185 24803
rect 13219 24769 13231 24803
rect 13740 24800 13768 24840
rect 14826 24800 14832 24812
rect 13740 24772 14832 24800
rect 13173 24763 13231 24769
rect 9272 24704 10824 24732
rect 11164 24704 13124 24732
rect 9272 24692 9278 24704
rect 4338 24624 4344 24676
rect 4396 24624 4402 24676
rect 11164 24608 11192 24704
rect 4157 24599 4215 24605
rect 4157 24565 4169 24599
rect 4203 24596 4215 24599
rect 4522 24596 4528 24608
rect 4203 24568 4528 24596
rect 4203 24565 4215 24568
rect 4157 24559 4215 24565
rect 4522 24556 4528 24568
rect 4580 24556 4586 24608
rect 6362 24556 6368 24608
rect 6420 24556 6426 24608
rect 11146 24556 11152 24608
rect 11204 24556 11210 24608
rect 11698 24556 11704 24608
rect 11756 24556 11762 24608
rect 11974 24556 11980 24608
rect 12032 24596 12038 24608
rect 12342 24596 12348 24608
rect 12032 24568 12348 24596
rect 12032 24556 12038 24568
rect 12342 24556 12348 24568
rect 12400 24596 12406 24608
rect 12897 24599 12955 24605
rect 12897 24596 12909 24599
rect 12400 24568 12909 24596
rect 12400 24556 12406 24568
rect 12897 24565 12909 24568
rect 12943 24565 12955 24599
rect 13188 24596 13216 24763
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 15838 24760 15844 24812
rect 15896 24760 15902 24812
rect 15933 24803 15991 24809
rect 15933 24769 15945 24803
rect 15979 24800 15991 24803
rect 16114 24800 16120 24812
rect 15979 24772 16120 24800
rect 15979 24769 15991 24772
rect 15933 24763 15991 24769
rect 16114 24760 16120 24772
rect 16172 24760 16178 24812
rect 16390 24760 16396 24812
rect 16448 24800 16454 24812
rect 16448 24772 17618 24800
rect 16448 24760 16454 24772
rect 19978 24760 19984 24812
rect 20036 24760 20042 24812
rect 20990 24760 20996 24812
rect 21048 24760 21054 24812
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 23385 24803 23443 24809
rect 21232 24772 23060 24800
rect 21232 24760 21238 24772
rect 15749 24735 15807 24741
rect 15749 24701 15761 24735
rect 15795 24732 15807 24735
rect 17221 24735 17279 24741
rect 17221 24732 17233 24735
rect 15795 24704 17233 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 17221 24701 17233 24704
rect 17267 24732 17279 24735
rect 17678 24732 17684 24744
rect 17267 24704 17684 24732
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 17678 24692 17684 24704
rect 17736 24692 17742 24744
rect 18690 24692 18696 24744
rect 18748 24692 18754 24744
rect 18969 24735 19027 24741
rect 18969 24701 18981 24735
rect 19015 24701 19027 24735
rect 18969 24695 19027 24701
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24732 20223 24735
rect 20346 24732 20352 24744
rect 20211 24704 20352 24732
rect 20211 24701 20223 24704
rect 20165 24695 20223 24701
rect 17126 24624 17132 24676
rect 17184 24664 17190 24676
rect 17184 24636 17724 24664
rect 17184 24624 17190 24636
rect 13633 24599 13691 24605
rect 13633 24596 13645 24599
rect 13188 24568 13645 24596
rect 12897 24559 12955 24565
rect 13633 24565 13645 24568
rect 13679 24596 13691 24599
rect 14826 24596 14832 24608
rect 13679 24568 14832 24596
rect 13679 24565 13691 24568
rect 13633 24559 13691 24565
rect 14826 24556 14832 24568
rect 14884 24556 14890 24608
rect 16301 24599 16359 24605
rect 16301 24565 16313 24599
rect 16347 24596 16359 24599
rect 16574 24596 16580 24608
rect 16347 24568 16580 24596
rect 16347 24565 16359 24568
rect 16301 24559 16359 24565
rect 16574 24556 16580 24568
rect 16632 24556 16638 24608
rect 17696 24596 17724 24636
rect 18984 24596 19012 24695
rect 20346 24692 20352 24704
rect 20404 24692 20410 24744
rect 20901 24735 20959 24741
rect 20901 24701 20913 24735
rect 20947 24701 20959 24735
rect 20901 24695 20959 24701
rect 22925 24735 22983 24741
rect 22925 24701 22937 24735
rect 22971 24701 22983 24735
rect 23032 24732 23060 24772
rect 23385 24769 23397 24803
rect 23431 24800 23443 24803
rect 23842 24800 23848 24812
rect 23431 24772 23848 24800
rect 23431 24769 23443 24772
rect 23385 24763 23443 24769
rect 23842 24760 23848 24772
rect 23900 24760 23906 24812
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24769 23995 24803
rect 23937 24763 23995 24769
rect 23952 24732 23980 24763
rect 23032 24704 23980 24732
rect 22925 24695 22983 24701
rect 19150 24624 19156 24676
rect 19208 24664 19214 24676
rect 19521 24667 19579 24673
rect 19521 24664 19533 24667
rect 19208 24636 19533 24664
rect 19208 24624 19214 24636
rect 19521 24633 19533 24636
rect 19567 24633 19579 24667
rect 20916 24664 20944 24695
rect 22830 24664 22836 24676
rect 20916 24636 22836 24664
rect 19521 24627 19579 24633
rect 22830 24624 22836 24636
rect 22888 24624 22894 24676
rect 22940 24664 22968 24695
rect 24670 24692 24676 24744
rect 24728 24692 24734 24744
rect 24854 24664 24860 24676
rect 22940 24636 24860 24664
rect 24854 24624 24860 24636
rect 24912 24624 24918 24676
rect 19334 24596 19340 24608
rect 17696 24568 19340 24596
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 21450 24556 21456 24608
rect 21508 24556 21514 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 5353 24395 5411 24401
rect 5353 24361 5365 24395
rect 5399 24392 5411 24395
rect 6086 24392 6092 24404
rect 5399 24364 6092 24392
rect 5399 24361 5411 24364
rect 5353 24355 5411 24361
rect 6086 24352 6092 24364
rect 6144 24392 6150 24404
rect 6270 24392 6276 24404
rect 6144 24364 6276 24392
rect 6144 24352 6150 24364
rect 6270 24352 6276 24364
rect 6328 24352 6334 24404
rect 10873 24395 10931 24401
rect 10873 24392 10885 24395
rect 10244 24364 10885 24392
rect 7098 24216 7104 24268
rect 7156 24256 7162 24268
rect 8386 24256 8392 24268
rect 7156 24228 8392 24256
rect 7156 24216 7162 24228
rect 8386 24216 8392 24228
rect 8444 24216 8450 24268
rect 10244 24265 10272 24364
rect 10873 24361 10885 24364
rect 10919 24392 10931 24395
rect 14918 24392 14924 24404
rect 10919 24364 14924 24392
rect 10919 24361 10931 24364
rect 10873 24355 10931 24361
rect 14918 24352 14924 24364
rect 14976 24352 14982 24404
rect 15746 24352 15752 24404
rect 15804 24392 15810 24404
rect 18690 24392 18696 24404
rect 15804 24364 18696 24392
rect 15804 24352 15810 24364
rect 18690 24352 18696 24364
rect 18748 24352 18754 24404
rect 23382 24392 23388 24404
rect 21284 24364 23388 24392
rect 10229 24259 10287 24265
rect 10229 24225 10241 24259
rect 10275 24225 10287 24259
rect 10229 24219 10287 24225
rect 10318 24216 10324 24268
rect 10376 24216 10382 24268
rect 12434 24256 12440 24268
rect 11440 24228 12440 24256
rect 11440 24200 11468 24228
rect 12434 24216 12440 24228
rect 12492 24216 12498 24268
rect 17126 24216 17132 24268
rect 17184 24216 17190 24268
rect 20165 24259 20223 24265
rect 20165 24225 20177 24259
rect 20211 24256 20223 24259
rect 20530 24256 20536 24268
rect 20211 24228 20536 24256
rect 20211 24225 20223 24228
rect 20165 24219 20223 24225
rect 20530 24216 20536 24228
rect 20588 24216 20594 24268
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 3602 24188 3608 24200
rect 2271 24160 3608 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 3602 24148 3608 24160
rect 3660 24148 3666 24200
rect 4154 24148 4160 24200
rect 4212 24188 4218 24200
rect 4249 24191 4307 24197
rect 4249 24188 4261 24191
rect 4212 24160 4261 24188
rect 4212 24148 4218 24160
rect 4249 24157 4261 24160
rect 4295 24157 4307 24191
rect 4249 24151 4307 24157
rect 7650 24148 7656 24200
rect 7708 24188 7714 24200
rect 8205 24191 8263 24197
rect 8205 24188 8217 24191
rect 7708 24160 8217 24188
rect 7708 24148 7714 24160
rect 8205 24157 8217 24160
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 9306 24148 9312 24200
rect 9364 24188 9370 24200
rect 11422 24188 11428 24200
rect 9364 24160 11428 24188
rect 9364 24148 9370 24160
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 17862 24148 17868 24200
rect 17920 24188 17926 24200
rect 18233 24191 18291 24197
rect 18233 24188 18245 24191
rect 17920 24160 18245 24188
rect 17920 24148 17926 24160
rect 18233 24157 18245 24160
rect 18279 24157 18291 24191
rect 18233 24151 18291 24157
rect 19334 24148 19340 24200
rect 19392 24188 19398 24200
rect 19889 24191 19947 24197
rect 19889 24188 19901 24191
rect 19392 24160 19901 24188
rect 19392 24148 19398 24160
rect 19889 24157 19901 24160
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 6362 24080 6368 24132
rect 6420 24120 6426 24132
rect 6825 24123 6883 24129
rect 6420 24092 6500 24120
rect 6420 24080 6426 24092
rect 1762 24012 1768 24064
rect 1820 24052 1826 24064
rect 2041 24055 2099 24061
rect 2041 24052 2053 24055
rect 1820 24024 2053 24052
rect 1820 24012 1826 24024
rect 2041 24021 2053 24024
rect 2087 24021 2099 24055
rect 2041 24015 2099 24021
rect 4614 24012 4620 24064
rect 4672 24052 4678 24064
rect 4893 24055 4951 24061
rect 4893 24052 4905 24055
rect 4672 24024 4905 24052
rect 4672 24012 4678 24024
rect 4893 24021 4905 24024
rect 4939 24021 4951 24055
rect 6472 24052 6500 24092
rect 6825 24089 6837 24123
rect 6871 24120 6883 24123
rect 7561 24123 7619 24129
rect 7561 24120 7573 24123
rect 6871 24092 7573 24120
rect 6871 24089 6883 24092
rect 6825 24083 6883 24089
rect 7561 24089 7573 24092
rect 7607 24089 7619 24123
rect 7561 24083 7619 24089
rect 11698 24080 11704 24132
rect 11756 24080 11762 24132
rect 12342 24080 12348 24132
rect 12400 24080 12406 24132
rect 16390 24080 16396 24132
rect 16448 24120 16454 24132
rect 16853 24123 16911 24129
rect 16448 24092 16804 24120
rect 16448 24080 16454 24092
rect 7466 24052 7472 24064
rect 6472 24024 7472 24052
rect 4893 24015 4951 24021
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 8846 24012 8852 24064
rect 8904 24052 8910 24064
rect 9769 24055 9827 24061
rect 9769 24052 9781 24055
rect 8904 24024 9781 24052
rect 8904 24012 8910 24024
rect 9769 24021 9781 24024
rect 9815 24021 9827 24055
rect 9769 24015 9827 24021
rect 9950 24012 9956 24064
rect 10008 24052 10014 24064
rect 10137 24055 10195 24061
rect 10137 24052 10149 24055
rect 10008 24024 10149 24052
rect 10008 24012 10014 24024
rect 10137 24021 10149 24024
rect 10183 24021 10195 24055
rect 10137 24015 10195 24021
rect 13173 24055 13231 24061
rect 13173 24021 13185 24055
rect 13219 24052 13231 24055
rect 13814 24052 13820 24064
rect 13219 24024 13820 24052
rect 13219 24021 13231 24024
rect 13173 24015 13231 24021
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 15381 24055 15439 24061
rect 15381 24021 15393 24055
rect 15427 24052 15439 24055
rect 16022 24052 16028 24064
rect 15427 24024 16028 24052
rect 15427 24021 15439 24024
rect 15381 24015 15439 24021
rect 16022 24012 16028 24024
rect 16080 24012 16086 24064
rect 16776 24052 16804 24092
rect 16853 24089 16865 24123
rect 16899 24120 16911 24123
rect 17589 24123 17647 24129
rect 17589 24120 17601 24123
rect 16899 24092 17601 24120
rect 16899 24089 16911 24092
rect 16853 24083 16911 24089
rect 17589 24089 17601 24092
rect 17635 24089 17647 24123
rect 17589 24083 17647 24089
rect 20272 24092 20654 24120
rect 20272 24052 20300 24092
rect 16776 24024 20300 24052
rect 20548 24052 20576 24092
rect 21284 24052 21312 24364
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 21634 24284 21640 24336
rect 21692 24284 21698 24336
rect 24026 24148 24032 24200
rect 24084 24148 24090 24200
rect 22830 24080 22836 24132
rect 22888 24080 22894 24132
rect 24394 24080 24400 24132
rect 24452 24120 24458 24132
rect 24949 24123 25007 24129
rect 24949 24120 24961 24123
rect 24452 24092 24961 24120
rect 24452 24080 24458 24092
rect 24949 24089 24961 24092
rect 24995 24120 25007 24123
rect 25317 24123 25375 24129
rect 25317 24120 25329 24123
rect 24995 24092 25329 24120
rect 24995 24089 25007 24092
rect 24949 24083 25007 24089
rect 25317 24089 25329 24092
rect 25363 24089 25375 24123
rect 25317 24083 25375 24089
rect 20548 24024 21312 24052
rect 22738 24012 22744 24064
rect 22796 24052 22802 24064
rect 23290 24052 23296 24064
rect 22796 24024 23296 24052
rect 22796 24012 22802 24024
rect 23290 24012 23296 24024
rect 23348 24012 23354 24064
rect 23382 24012 23388 24064
rect 23440 24052 23446 24064
rect 24670 24052 24676 24064
rect 23440 24024 24676 24052
rect 23440 24012 23446 24024
rect 24670 24012 24676 24024
rect 24728 24012 24734 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 4246 23857 4252 23860
rect 4203 23851 4252 23857
rect 4203 23817 4215 23851
rect 4249 23817 4252 23851
rect 4203 23811 4252 23817
rect 4246 23808 4252 23811
rect 4304 23808 4310 23860
rect 9122 23808 9128 23860
rect 9180 23848 9186 23860
rect 9401 23851 9459 23857
rect 9401 23848 9413 23851
rect 9180 23820 9413 23848
rect 9180 23808 9186 23820
rect 9401 23817 9413 23820
rect 9447 23817 9459 23851
rect 9401 23811 9459 23817
rect 9416 23780 9444 23811
rect 9950 23808 9956 23860
rect 10008 23808 10014 23860
rect 10686 23848 10692 23860
rect 10060 23820 10692 23848
rect 10060 23780 10088 23820
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 12066 23808 12072 23860
rect 12124 23848 12130 23860
rect 12161 23851 12219 23857
rect 12161 23848 12173 23851
rect 12124 23820 12173 23848
rect 12124 23808 12130 23820
rect 12161 23817 12173 23820
rect 12207 23817 12219 23851
rect 12161 23811 12219 23817
rect 16114 23808 16120 23860
rect 16172 23848 16178 23860
rect 16301 23851 16359 23857
rect 16301 23848 16313 23851
rect 16172 23820 16313 23848
rect 16172 23808 16178 23820
rect 16301 23817 16313 23820
rect 16347 23817 16359 23851
rect 16301 23811 16359 23817
rect 16574 23808 16580 23860
rect 16632 23848 16638 23860
rect 17221 23851 17279 23857
rect 17221 23848 17233 23851
rect 16632 23820 17233 23848
rect 16632 23808 16638 23820
rect 17221 23817 17233 23820
rect 17267 23817 17279 23851
rect 17221 23811 17279 23817
rect 17313 23851 17371 23857
rect 17313 23817 17325 23851
rect 17359 23848 17371 23851
rect 17494 23848 17500 23860
rect 17359 23820 17500 23848
rect 17359 23817 17371 23820
rect 17313 23811 17371 23817
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 20990 23808 20996 23860
rect 21048 23848 21054 23860
rect 21453 23851 21511 23857
rect 21453 23848 21465 23851
rect 21048 23820 21465 23848
rect 21048 23808 21054 23820
rect 21453 23817 21465 23820
rect 21499 23848 21511 23851
rect 21542 23848 21548 23860
rect 21499 23820 21548 23848
rect 21499 23817 21511 23820
rect 21453 23811 21511 23817
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22373 23851 22431 23857
rect 22373 23817 22385 23851
rect 22419 23848 22431 23851
rect 23566 23848 23572 23860
rect 22419 23820 23572 23848
rect 22419 23817 22431 23820
rect 22373 23811 22431 23817
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 11146 23780 11152 23792
rect 9416 23752 10088 23780
rect 10612 23752 11152 23780
rect 4062 23672 4068 23724
rect 4120 23721 4126 23724
rect 4120 23715 4158 23721
rect 4146 23681 4158 23715
rect 4120 23675 4158 23681
rect 4120 23672 4126 23675
rect 10612 23653 10640 23752
rect 11146 23740 11152 23752
rect 11204 23740 11210 23792
rect 15933 23783 15991 23789
rect 15933 23749 15945 23783
rect 15979 23780 15991 23783
rect 18049 23783 18107 23789
rect 18049 23780 18061 23783
rect 15979 23752 18061 23780
rect 15979 23749 15991 23752
rect 15933 23743 15991 23749
rect 18049 23749 18061 23752
rect 18095 23749 18107 23783
rect 20898 23780 20904 23792
rect 20838 23752 20904 23780
rect 18049 23743 18107 23749
rect 20898 23740 20904 23752
rect 20956 23740 20962 23792
rect 21082 23740 21088 23792
rect 21140 23780 21146 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 21140 23752 22293 23780
rect 21140 23740 21146 23752
rect 22281 23749 22293 23752
rect 22327 23749 22339 23783
rect 23201 23783 23259 23789
rect 23201 23780 23213 23783
rect 22281 23743 22339 23749
rect 22388 23752 23213 23780
rect 22388 23724 22416 23752
rect 23201 23749 23213 23752
rect 23247 23749 23259 23783
rect 24670 23780 24676 23792
rect 24426 23752 24676 23780
rect 23201 23743 23259 23749
rect 24670 23740 24676 23752
rect 24728 23740 24734 23792
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 11330 23712 11336 23724
rect 10827 23684 11336 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 11330 23672 11336 23684
rect 11388 23672 11394 23724
rect 12069 23715 12127 23721
rect 12069 23681 12081 23715
rect 12115 23712 12127 23715
rect 12250 23712 12256 23724
rect 12115 23684 12256 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 12250 23672 12256 23684
rect 12308 23672 12314 23724
rect 13814 23672 13820 23724
rect 13872 23672 13878 23724
rect 15289 23715 15347 23721
rect 15289 23681 15301 23715
rect 15335 23712 15347 23715
rect 19058 23712 19064 23724
rect 15335 23684 15884 23712
rect 15335 23681 15347 23684
rect 15289 23675 15347 23681
rect 10597 23647 10655 23653
rect 10597 23613 10609 23647
rect 10643 23613 10655 23647
rect 10597 23607 10655 23613
rect 11882 23604 11888 23656
rect 11940 23604 11946 23656
rect 13722 23644 13728 23656
rect 12406 23616 13728 23644
rect 11149 23579 11207 23585
rect 11149 23545 11161 23579
rect 11195 23576 11207 23579
rect 12406 23576 12434 23616
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 15746 23604 15752 23656
rect 15804 23604 15810 23656
rect 15856 23653 15884 23684
rect 15948 23684 19064 23712
rect 15841 23647 15899 23653
rect 15841 23613 15853 23647
rect 15887 23644 15899 23647
rect 15948 23644 15976 23684
rect 19058 23672 19064 23684
rect 19116 23672 19122 23724
rect 19334 23672 19340 23724
rect 19392 23672 19398 23724
rect 21266 23672 21272 23724
rect 21324 23712 21330 23724
rect 22370 23712 22376 23724
rect 21324 23684 22376 23712
rect 21324 23672 21330 23684
rect 22370 23672 22376 23684
rect 22428 23672 22434 23724
rect 15887 23616 15976 23644
rect 15887 23613 15899 23616
rect 15841 23607 15899 23613
rect 16022 23604 16028 23656
rect 16080 23644 16086 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16080 23616 17417 23644
rect 16080 23604 16086 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 19610 23604 19616 23656
rect 19668 23604 19674 23656
rect 20622 23604 20628 23656
rect 20680 23644 20686 23656
rect 21085 23647 21143 23653
rect 21085 23644 21097 23647
rect 20680 23616 21097 23644
rect 20680 23604 20686 23616
rect 21085 23613 21097 23616
rect 21131 23613 21143 23647
rect 21085 23607 21143 23613
rect 22186 23604 22192 23656
rect 22244 23644 22250 23656
rect 22925 23647 22983 23653
rect 22925 23644 22937 23647
rect 22244 23616 22937 23644
rect 22244 23604 22250 23616
rect 22925 23613 22937 23616
rect 22971 23613 22983 23647
rect 22925 23607 22983 23613
rect 11195 23548 12434 23576
rect 12529 23579 12587 23585
rect 11195 23545 11207 23548
rect 11149 23539 11207 23545
rect 12529 23545 12541 23579
rect 12575 23576 12587 23579
rect 16574 23576 16580 23588
rect 12575 23548 16580 23576
rect 12575 23545 12587 23548
rect 12529 23539 12587 23545
rect 16574 23536 16580 23548
rect 16632 23536 16638 23588
rect 7285 23511 7343 23517
rect 7285 23477 7297 23511
rect 7331 23508 7343 23511
rect 7466 23508 7472 23520
rect 7331 23480 7472 23508
rect 7331 23477 7343 23480
rect 7285 23471 7343 23477
rect 7466 23468 7472 23480
rect 7524 23468 7530 23520
rect 13173 23511 13231 23517
rect 13173 23477 13185 23511
rect 13219 23508 13231 23511
rect 13354 23508 13360 23520
rect 13219 23480 13360 23508
rect 13219 23477 13231 23480
rect 13173 23471 13231 23477
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 16390 23468 16396 23520
rect 16448 23508 16454 23520
rect 16853 23511 16911 23517
rect 16853 23508 16865 23511
rect 16448 23480 16865 23508
rect 16448 23468 16454 23480
rect 16853 23477 16865 23480
rect 16899 23477 16911 23511
rect 22940 23508 22968 23607
rect 23290 23604 23296 23656
rect 23348 23644 23354 23656
rect 24673 23647 24731 23653
rect 24673 23644 24685 23647
rect 23348 23616 24685 23644
rect 23348 23604 23354 23616
rect 24673 23613 24685 23616
rect 24719 23613 24731 23647
rect 24673 23607 24731 23613
rect 23290 23508 23296 23520
rect 22940 23480 23296 23508
rect 16853 23471 16911 23477
rect 23290 23468 23296 23480
rect 23348 23468 23354 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 4430 23264 4436 23316
rect 4488 23264 4494 23316
rect 15194 23264 15200 23316
rect 15252 23304 15258 23316
rect 15381 23307 15439 23313
rect 15381 23304 15393 23307
rect 15252 23276 15393 23304
rect 15252 23264 15258 23276
rect 15381 23273 15393 23276
rect 15427 23304 15439 23307
rect 16758 23304 16764 23316
rect 15427 23276 16764 23304
rect 15427 23273 15439 23276
rect 15381 23267 15439 23273
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 18690 23264 18696 23316
rect 18748 23264 18754 23316
rect 19610 23264 19616 23316
rect 19668 23304 19674 23316
rect 20073 23307 20131 23313
rect 20073 23304 20085 23307
rect 19668 23276 20085 23304
rect 19668 23264 19674 23276
rect 20073 23273 20085 23276
rect 20119 23273 20131 23307
rect 20073 23267 20131 23273
rect 3418 23196 3424 23248
rect 3476 23196 3482 23248
rect 9674 23236 9680 23248
rect 8312 23208 9680 23236
rect 2774 23128 2780 23180
rect 2832 23128 2838 23180
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23168 3295 23171
rect 3436 23168 3464 23196
rect 3283 23140 3556 23168
rect 3283 23137 3295 23140
rect 3237 23131 3295 23137
rect 3418 23060 3424 23112
rect 3476 23060 3482 23112
rect 3528 23044 3556 23140
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 6641 23171 6699 23177
rect 6641 23137 6653 23171
rect 6687 23168 6699 23171
rect 7650 23168 7656 23180
rect 6687 23140 7656 23168
rect 6687 23137 6699 23140
rect 6641 23131 6699 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 8113 23171 8171 23177
rect 8113 23137 8125 23171
rect 8159 23168 8171 23171
rect 8312 23168 8340 23208
rect 9674 23196 9680 23208
rect 9732 23236 9738 23248
rect 10318 23236 10324 23248
rect 9732 23208 10324 23236
rect 9732 23196 9738 23208
rect 10318 23196 10324 23208
rect 10376 23196 10382 23248
rect 13173 23239 13231 23245
rect 13173 23205 13185 23239
rect 13219 23236 13231 23239
rect 15013 23239 15071 23245
rect 13219 23208 14964 23236
rect 13219 23205 13231 23208
rect 13173 23199 13231 23205
rect 8159 23140 8340 23168
rect 8159 23137 8171 23140
rect 8113 23131 8171 23137
rect 8386 23128 8392 23180
rect 8444 23128 8450 23180
rect 10226 23128 10232 23180
rect 10284 23128 10290 23180
rect 11330 23128 11336 23180
rect 11388 23168 11394 23180
rect 11425 23171 11483 23177
rect 11425 23168 11437 23171
rect 11388 23140 11437 23168
rect 11388 23128 11394 23140
rect 11425 23137 11437 23140
rect 11471 23137 11483 23171
rect 12621 23171 12679 23177
rect 12621 23168 12633 23171
rect 11425 23131 11483 23137
rect 12406 23140 12633 23168
rect 9766 23060 9772 23112
rect 9824 23100 9830 23112
rect 12406 23100 12434 23140
rect 12621 23137 12633 23140
rect 12667 23137 12679 23171
rect 12621 23131 12679 23137
rect 9824 23072 12434 23100
rect 9824 23060 9830 23072
rect 2774 22992 2780 23044
rect 2832 23032 2838 23044
rect 3510 23032 3516 23044
rect 2832 23004 3516 23032
rect 2832 22992 2838 23004
rect 3510 22992 3516 23004
rect 3568 22992 3574 23044
rect 5905 23035 5963 23041
rect 5905 23001 5917 23035
rect 5951 23032 5963 23035
rect 5951 23004 6868 23032
rect 5951 23001 5963 23004
rect 5905 22995 5963 23001
rect 4430 22924 4436 22976
rect 4488 22964 4494 22976
rect 5445 22967 5503 22973
rect 5445 22964 5457 22967
rect 4488 22936 5457 22964
rect 4488 22924 4494 22936
rect 5445 22933 5457 22936
rect 5491 22933 5503 22967
rect 5445 22927 5503 22933
rect 5810 22924 5816 22976
rect 5868 22924 5874 22976
rect 6840 22964 6868 23004
rect 7466 22992 7472 23044
rect 7524 22992 7530 23044
rect 9953 23035 10011 23041
rect 9953 23001 9965 23035
rect 9999 23032 10011 23035
rect 10781 23035 10839 23041
rect 10781 23032 10793 23035
rect 9999 23004 10793 23032
rect 9999 23001 10011 23004
rect 9953 22995 10011 23001
rect 10781 23001 10793 23004
rect 10827 23001 10839 23035
rect 10781 22995 10839 23001
rect 12526 22992 12532 23044
rect 12584 22992 12590 23044
rect 7834 22964 7840 22976
rect 6840 22936 7840 22964
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 8478 22924 8484 22976
rect 8536 22964 8542 22976
rect 8665 22967 8723 22973
rect 8665 22964 8677 22967
rect 8536 22936 8677 22964
rect 8536 22924 8542 22936
rect 8665 22933 8677 22936
rect 8711 22933 8723 22967
rect 8665 22927 8723 22933
rect 9582 22924 9588 22976
rect 9640 22924 9646 22976
rect 10045 22967 10103 22973
rect 10045 22933 10057 22967
rect 10091 22964 10103 22967
rect 10502 22964 10508 22976
rect 10091 22936 10508 22964
rect 10091 22933 10103 22936
rect 10045 22927 10103 22933
rect 10502 22924 10508 22936
rect 10560 22924 10566 22976
rect 11054 22924 11060 22976
rect 11112 22964 11118 22976
rect 12069 22967 12127 22973
rect 12069 22964 12081 22967
rect 11112 22936 12081 22964
rect 11112 22924 11118 22936
rect 12069 22933 12081 22936
rect 12115 22933 12127 22967
rect 12069 22927 12127 22933
rect 12437 22967 12495 22973
rect 12437 22933 12449 22967
rect 12483 22964 12495 22967
rect 13188 22964 13216 23199
rect 13814 23128 13820 23180
rect 13872 23168 13878 23180
rect 14369 23171 14427 23177
rect 14369 23168 14381 23171
rect 13872 23140 14381 23168
rect 13872 23128 13878 23140
rect 14369 23137 14381 23140
rect 14415 23137 14427 23171
rect 14369 23131 14427 23137
rect 14550 23128 14556 23180
rect 14608 23128 14614 23180
rect 14936 23168 14964 23208
rect 15013 23205 15025 23239
rect 15059 23236 15071 23239
rect 17402 23236 17408 23248
rect 15059 23208 17408 23236
rect 15059 23205 15071 23208
rect 15013 23199 15071 23205
rect 17402 23196 17408 23208
rect 17460 23196 17466 23248
rect 18708 23236 18736 23264
rect 21082 23236 21088 23248
rect 18708 23208 21088 23236
rect 21082 23196 21088 23208
rect 21140 23196 21146 23248
rect 22738 23236 22744 23248
rect 21652 23208 22744 23236
rect 17770 23168 17776 23180
rect 14936 23140 17776 23168
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 21652 23177 21680 23208
rect 22738 23196 22744 23208
rect 22796 23196 22802 23248
rect 21637 23171 21695 23177
rect 21637 23137 21649 23171
rect 21683 23137 21695 23171
rect 21637 23131 21695 23137
rect 21726 23128 21732 23180
rect 21784 23128 21790 23180
rect 22066 23140 24624 23168
rect 13722 23060 13728 23112
rect 13780 23100 13786 23112
rect 14645 23103 14703 23109
rect 14645 23100 14657 23103
rect 13780 23072 14657 23100
rect 13780 23060 13786 23072
rect 14645 23069 14657 23072
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 18598 23060 18604 23112
rect 18656 23100 18662 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 18656 23072 19441 23100
rect 18656 23060 18662 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21542 23100 21548 23112
rect 20864 23072 21548 23100
rect 20864 23060 20870 23072
rect 21542 23060 21548 23072
rect 21600 23100 21606 23112
rect 22066 23100 22094 23140
rect 21600 23072 22094 23100
rect 23109 23103 23167 23109
rect 21600 23060 21606 23072
rect 23109 23069 23121 23103
rect 23155 23100 23167 23103
rect 23382 23100 23388 23112
rect 23155 23072 23388 23100
rect 23155 23069 23167 23072
rect 23109 23063 23167 23069
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23100 24087 23103
rect 24118 23100 24124 23112
rect 24075 23072 24124 23100
rect 24075 23069 24087 23072
rect 24029 23063 24087 23069
rect 24118 23060 24124 23072
rect 24176 23060 24182 23112
rect 24596 23109 24624 23140
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 17494 22992 17500 23044
rect 17552 23032 17558 23044
rect 19058 23032 19064 23044
rect 17552 23004 19064 23032
rect 17552 22992 17558 23004
rect 19058 22992 19064 23004
rect 19116 22992 19122 23044
rect 20993 23035 21051 23041
rect 20993 23001 21005 23035
rect 21039 23032 21051 23035
rect 21821 23035 21879 23041
rect 21821 23032 21833 23035
rect 21039 23004 21833 23032
rect 21039 23001 21051 23004
rect 20993 22995 21051 23001
rect 21821 23001 21833 23004
rect 21867 23001 21879 23035
rect 21821 22995 21879 23001
rect 12483 22936 13216 22964
rect 12483 22933 12495 22936
rect 12437 22927 12495 22933
rect 15838 22924 15844 22976
rect 15896 22964 15902 22976
rect 16206 22964 16212 22976
rect 15896 22936 16212 22964
rect 15896 22924 15902 22936
rect 16206 22924 16212 22936
rect 16264 22924 16270 22976
rect 16758 22924 16764 22976
rect 16816 22924 16822 22976
rect 18690 22924 18696 22976
rect 18748 22964 18754 22976
rect 18874 22964 18880 22976
rect 18748 22936 18880 22964
rect 18748 22924 18754 22936
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 20346 22924 20352 22976
rect 20404 22924 20410 22976
rect 22186 22924 22192 22976
rect 22244 22924 22250 22976
rect 25222 22924 25228 22976
rect 25280 22924 25286 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 3510 22720 3516 22772
rect 3568 22760 3574 22772
rect 4617 22763 4675 22769
rect 4617 22760 4629 22763
rect 3568 22732 4629 22760
rect 3568 22720 3574 22732
rect 4617 22729 4629 22732
rect 4663 22729 4675 22763
rect 4617 22723 4675 22729
rect 5810 22720 5816 22772
rect 5868 22760 5874 22772
rect 7285 22763 7343 22769
rect 7285 22760 7297 22763
rect 5868 22732 7297 22760
rect 5868 22720 5874 22732
rect 7285 22729 7297 22732
rect 7331 22729 7343 22763
rect 7285 22723 7343 22729
rect 7653 22763 7711 22769
rect 7653 22729 7665 22763
rect 7699 22760 7711 22763
rect 8846 22760 8852 22772
rect 7699 22732 8852 22760
rect 7699 22729 7711 22732
rect 7653 22723 7711 22729
rect 8846 22720 8852 22732
rect 8904 22720 8910 22772
rect 10502 22720 10508 22772
rect 10560 22760 10566 22772
rect 11514 22760 11520 22772
rect 10560 22732 11520 22760
rect 10560 22720 10566 22732
rect 11514 22720 11520 22732
rect 11572 22720 11578 22772
rect 12526 22760 12532 22772
rect 12406 22732 12532 22760
rect 8386 22652 8392 22704
rect 8444 22692 8450 22704
rect 8573 22695 8631 22701
rect 8573 22692 8585 22695
rect 8444 22664 8585 22692
rect 8444 22652 8450 22664
rect 8573 22661 8585 22664
rect 8619 22661 8631 22695
rect 8573 22655 8631 22661
rect 3881 22627 3939 22633
rect 3881 22593 3893 22627
rect 3927 22624 3939 22627
rect 4430 22624 4436 22636
rect 3927 22596 4436 22624
rect 3927 22593 3939 22596
rect 3881 22587 3939 22593
rect 4430 22584 4436 22596
rect 4488 22584 4494 22636
rect 4522 22584 4528 22636
rect 4580 22624 4586 22636
rect 5077 22627 5135 22633
rect 5077 22624 5089 22627
rect 4580 22596 5089 22624
rect 4580 22584 4586 22596
rect 5077 22593 5089 22596
rect 5123 22624 5135 22627
rect 5534 22624 5540 22636
rect 5123 22596 5540 22624
rect 5123 22593 5135 22596
rect 5077 22587 5135 22593
rect 5534 22584 5540 22596
rect 5592 22584 5598 22636
rect 7745 22627 7803 22633
rect 7745 22593 7757 22627
rect 7791 22624 7803 22627
rect 8846 22624 8852 22636
rect 7791 22596 8852 22624
rect 7791 22593 7803 22596
rect 7745 22587 7803 22593
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22624 9459 22627
rect 9447 22596 9812 22624
rect 9447 22593 9459 22596
rect 9401 22587 9459 22593
rect 7650 22516 7656 22568
rect 7708 22556 7714 22568
rect 7837 22559 7895 22565
rect 7837 22556 7849 22559
rect 7708 22528 7849 22556
rect 7708 22516 7714 22528
rect 7837 22525 7849 22528
rect 7883 22556 7895 22559
rect 8202 22556 8208 22568
rect 7883 22528 8208 22556
rect 7883 22525 7895 22528
rect 7837 22519 7895 22525
rect 8202 22516 8208 22528
rect 8260 22516 8266 22568
rect 9784 22497 9812 22596
rect 9769 22491 9827 22497
rect 9769 22457 9781 22491
rect 9815 22488 9827 22491
rect 10778 22488 10784 22500
rect 9815 22460 10784 22488
rect 9815 22457 9827 22460
rect 9769 22451 9827 22457
rect 10778 22448 10784 22460
rect 10836 22448 10842 22500
rect 4065 22423 4123 22429
rect 4065 22389 4077 22423
rect 4111 22420 4123 22423
rect 4246 22420 4252 22432
rect 4111 22392 4252 22420
rect 4111 22389 4123 22392
rect 4065 22383 4123 22389
rect 4246 22380 4252 22392
rect 4304 22380 4310 22432
rect 4985 22423 5043 22429
rect 4985 22389 4997 22423
rect 5031 22420 5043 22423
rect 6270 22420 6276 22432
rect 5031 22392 6276 22420
rect 5031 22389 5043 22392
rect 4985 22383 5043 22389
rect 6270 22380 6276 22392
rect 6328 22380 6334 22432
rect 11330 22380 11336 22432
rect 11388 22420 11394 22432
rect 11885 22423 11943 22429
rect 11885 22420 11897 22423
rect 11388 22392 11897 22420
rect 11388 22380 11394 22392
rect 11885 22389 11897 22392
rect 11931 22420 11943 22423
rect 12406 22420 12434 22732
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 13906 22720 13912 22772
rect 13964 22760 13970 22772
rect 13964 22732 15424 22760
rect 13964 22720 13970 22732
rect 13081 22695 13139 22701
rect 13081 22661 13093 22695
rect 13127 22692 13139 22695
rect 13354 22692 13360 22704
rect 13127 22664 13360 22692
rect 13127 22661 13139 22664
rect 13081 22655 13139 22661
rect 13354 22652 13360 22664
rect 13412 22652 13418 22704
rect 14458 22692 14464 22704
rect 14306 22664 14464 22692
rect 14458 22652 14464 22664
rect 14516 22692 14522 22704
rect 15010 22692 15016 22704
rect 14516 22664 15016 22692
rect 14516 22652 14522 22664
rect 15010 22652 15016 22664
rect 15068 22652 15074 22704
rect 15194 22652 15200 22704
rect 15252 22692 15258 22704
rect 15289 22695 15347 22701
rect 15289 22692 15301 22695
rect 15252 22664 15301 22692
rect 15252 22652 15258 22664
rect 15289 22661 15301 22664
rect 15335 22661 15347 22695
rect 15289 22655 15347 22661
rect 15396 22633 15424 22732
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 19426 22760 19432 22772
rect 18012 22732 19432 22760
rect 18012 22720 18018 22732
rect 19426 22720 19432 22732
rect 19484 22760 19490 22772
rect 20530 22760 20536 22772
rect 19484 22732 20536 22760
rect 19484 22720 19490 22732
rect 20530 22720 20536 22732
rect 20588 22720 20594 22772
rect 16776 22664 16988 22692
rect 15381 22627 15439 22633
rect 15381 22593 15393 22627
rect 15427 22624 15439 22627
rect 15838 22624 15844 22636
rect 15427 22596 15844 22624
rect 15427 22593 15439 22596
rect 15381 22587 15439 22593
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 12802 22516 12808 22568
rect 12860 22516 12866 22568
rect 15197 22559 15255 22565
rect 15197 22525 15209 22559
rect 15243 22556 15255 22559
rect 16776 22556 16804 22664
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 15243 22528 16804 22556
rect 15243 22525 15255 22528
rect 15197 22519 15255 22525
rect 16868 22488 16896 22587
rect 16960 22556 16988 22664
rect 19334 22652 19340 22704
rect 19392 22692 19398 22704
rect 19981 22695 20039 22701
rect 19981 22692 19993 22695
rect 19392 22664 19993 22692
rect 19392 22652 19398 22664
rect 19981 22661 19993 22664
rect 20027 22692 20039 22695
rect 20070 22692 20076 22704
rect 20027 22664 20076 22692
rect 20027 22661 20039 22664
rect 19981 22655 20039 22661
rect 20070 22652 20076 22664
rect 20128 22652 20134 22704
rect 20346 22652 20352 22704
rect 20404 22692 20410 22704
rect 20809 22695 20867 22701
rect 20809 22692 20821 22695
rect 20404 22664 20821 22692
rect 20404 22652 20410 22664
rect 20809 22661 20821 22664
rect 20855 22661 20867 22695
rect 20809 22655 20867 22661
rect 22002 22652 22008 22704
rect 22060 22692 22066 22704
rect 22060 22664 22678 22692
rect 22060 22652 22066 22664
rect 24118 22652 24124 22704
rect 24176 22692 24182 22704
rect 24397 22695 24455 22701
rect 24397 22692 24409 22695
rect 24176 22664 24409 22692
rect 24176 22652 24182 22664
rect 24397 22661 24409 22664
rect 24443 22661 24455 22695
rect 24397 22655 24455 22661
rect 17126 22584 17132 22636
rect 17184 22624 17190 22636
rect 17681 22627 17739 22633
rect 17681 22624 17693 22627
rect 17184 22596 17693 22624
rect 17184 22584 17190 22596
rect 17681 22593 17693 22596
rect 17727 22593 17739 22627
rect 17681 22587 17739 22593
rect 19058 22584 19064 22636
rect 19116 22624 19122 22636
rect 20990 22624 20996 22636
rect 19116 22596 20996 22624
rect 19116 22584 19122 22596
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 21082 22584 21088 22636
rect 21140 22624 21146 22636
rect 22097 22627 22155 22633
rect 22097 22624 22109 22627
rect 21140 22596 22109 22624
rect 21140 22584 21146 22596
rect 22097 22593 22109 22596
rect 22143 22593 22155 22627
rect 22097 22587 22155 22593
rect 17957 22559 18015 22565
rect 17957 22556 17969 22559
rect 16960 22528 17969 22556
rect 17957 22525 17969 22528
rect 18003 22556 18015 22559
rect 18690 22556 18696 22568
rect 18003 22528 18696 22556
rect 18003 22525 18015 22528
rect 17957 22519 18015 22525
rect 18690 22516 18696 22528
rect 18748 22516 18754 22568
rect 23842 22516 23848 22568
rect 23900 22516 23906 22568
rect 24121 22559 24179 22565
rect 24121 22525 24133 22559
rect 24167 22556 24179 22559
rect 24762 22556 24768 22568
rect 24167 22528 24768 22556
rect 24167 22525 24179 22528
rect 24121 22519 24179 22525
rect 20622 22488 20628 22500
rect 14108 22460 16896 22488
rect 19352 22460 20628 22488
rect 11931 22392 12434 22420
rect 11931 22389 11943 22392
rect 11885 22383 11943 22389
rect 12526 22380 12532 22432
rect 12584 22380 12590 22432
rect 12710 22380 12716 22432
rect 12768 22420 12774 22432
rect 14108 22420 14136 22460
rect 12768 22392 14136 22420
rect 12768 22380 12774 22392
rect 14458 22380 14464 22432
rect 14516 22420 14522 22432
rect 14553 22423 14611 22429
rect 14553 22420 14565 22423
rect 14516 22392 14565 22420
rect 14516 22380 14522 22392
rect 14553 22389 14565 22392
rect 14599 22420 14611 22423
rect 15102 22420 15108 22432
rect 14599 22392 15108 22420
rect 14599 22389 14611 22392
rect 14553 22383 14611 22389
rect 15102 22380 15108 22392
rect 15160 22380 15166 22432
rect 15749 22423 15807 22429
rect 15749 22389 15761 22423
rect 15795 22420 15807 22423
rect 16666 22420 16672 22432
rect 15795 22392 16672 22420
rect 15795 22389 15807 22392
rect 15749 22383 15807 22389
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 17037 22423 17095 22429
rect 17037 22389 17049 22423
rect 17083 22420 17095 22423
rect 19352 22420 19380 22460
rect 20622 22448 20628 22460
rect 20680 22448 20686 22500
rect 17083 22392 19380 22420
rect 17083 22389 17095 22392
rect 17037 22383 17095 22389
rect 23290 22380 23296 22432
rect 23348 22420 23354 22432
rect 24136 22420 24164 22519
rect 24762 22516 24768 22528
rect 24820 22516 24826 22568
rect 23348 22392 24164 22420
rect 23348 22380 23354 22392
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 4614 22225 4620 22228
rect 4604 22219 4620 22225
rect 4604 22185 4616 22219
rect 4604 22179 4620 22185
rect 4614 22176 4620 22179
rect 4672 22176 4678 22228
rect 15194 22176 15200 22228
rect 15252 22216 15258 22228
rect 19337 22219 19395 22225
rect 19337 22216 19349 22219
rect 15252 22188 19349 22216
rect 15252 22176 15258 22188
rect 19337 22185 19349 22188
rect 19383 22216 19395 22219
rect 19426 22216 19432 22228
rect 19383 22188 19432 22216
rect 19383 22185 19395 22188
rect 19337 22179 19395 22185
rect 19426 22176 19432 22188
rect 19484 22216 19490 22228
rect 20346 22216 20352 22228
rect 19484 22188 20352 22216
rect 19484 22176 19490 22188
rect 20346 22176 20352 22188
rect 20404 22176 20410 22228
rect 23842 22176 23848 22228
rect 23900 22216 23906 22228
rect 24581 22219 24639 22225
rect 24581 22216 24593 22219
rect 23900 22188 24593 22216
rect 23900 22176 23906 22188
rect 24581 22185 24593 22188
rect 24627 22185 24639 22219
rect 24581 22179 24639 22185
rect 12526 22108 12532 22160
rect 12584 22148 12590 22160
rect 13722 22148 13728 22160
rect 12584 22120 13728 22148
rect 12584 22108 12590 22120
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 5350 22080 5356 22092
rect 4387 22052 5356 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 5350 22040 5356 22052
rect 5408 22080 5414 22092
rect 7006 22080 7012 22092
rect 5408 22052 7012 22080
rect 5408 22040 5414 22052
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 7098 22040 7104 22092
rect 7156 22040 7162 22092
rect 11422 22040 11428 22092
rect 11480 22080 11486 22092
rect 11517 22083 11575 22089
rect 11517 22080 11529 22083
rect 11480 22052 11529 22080
rect 11480 22040 11486 22052
rect 11517 22049 11529 22052
rect 11563 22080 11575 22083
rect 12802 22080 12808 22092
rect 11563 22052 12808 22080
rect 11563 22049 11575 22052
rect 11517 22043 11575 22049
rect 12802 22040 12808 22052
rect 12860 22040 12866 22092
rect 13464 22089 13492 22120
rect 13722 22108 13728 22120
rect 13780 22108 13786 22160
rect 14277 22151 14335 22157
rect 14277 22117 14289 22151
rect 14323 22117 14335 22151
rect 14277 22111 14335 22117
rect 13449 22083 13507 22089
rect 13449 22049 13461 22083
rect 13495 22049 13507 22083
rect 13449 22043 13507 22049
rect 9214 21972 9220 22024
rect 9272 22012 9278 22024
rect 14292 22012 14320 22111
rect 15010 22108 15016 22160
rect 15068 22148 15074 22160
rect 15289 22151 15347 22157
rect 15289 22148 15301 22151
rect 15068 22120 15301 22148
rect 15068 22108 15074 22120
rect 15289 22117 15301 22120
rect 15335 22117 15347 22151
rect 15289 22111 15347 22117
rect 15838 22108 15844 22160
rect 15896 22108 15902 22160
rect 17954 22148 17960 22160
rect 16592 22120 17960 22148
rect 14642 22040 14648 22092
rect 14700 22080 14706 22092
rect 16592 22089 16620 22120
rect 17954 22108 17960 22120
rect 18012 22108 18018 22160
rect 18322 22148 18328 22160
rect 18064 22120 18328 22148
rect 18064 22089 18092 22120
rect 18322 22108 18328 22120
rect 18380 22108 18386 22160
rect 18690 22108 18696 22160
rect 18748 22148 18754 22160
rect 19242 22148 19248 22160
rect 18748 22120 19248 22148
rect 18748 22108 18754 22120
rect 19242 22108 19248 22120
rect 19300 22108 19306 22160
rect 14829 22083 14887 22089
rect 14829 22080 14841 22083
rect 14700 22052 14841 22080
rect 14700 22040 14706 22052
rect 14829 22049 14841 22052
rect 14875 22049 14887 22083
rect 14829 22043 14887 22049
rect 16577 22083 16635 22089
rect 16577 22049 16589 22083
rect 16623 22080 16635 22083
rect 18049 22083 18107 22089
rect 16623 22052 16657 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 18049 22049 18061 22083
rect 18095 22080 18107 22083
rect 18233 22083 18291 22089
rect 18095 22052 18129 22080
rect 18095 22049 18107 22052
rect 18049 22043 18107 22049
rect 18233 22049 18245 22083
rect 18279 22080 18291 22083
rect 18414 22080 18420 22092
rect 18279 22052 18420 22080
rect 18279 22049 18291 22052
rect 18233 22043 18291 22049
rect 18414 22040 18420 22052
rect 18472 22080 18478 22092
rect 18598 22080 18604 22092
rect 18472 22052 18604 22080
rect 18472 22040 18478 22052
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 20717 22083 20775 22089
rect 20717 22049 20729 22083
rect 20763 22080 20775 22083
rect 21269 22083 21327 22089
rect 21269 22080 21281 22083
rect 20763 22052 21281 22080
rect 20763 22049 20775 22052
rect 20717 22043 20775 22049
rect 21269 22049 21281 22052
rect 21315 22080 21327 22083
rect 23198 22080 23204 22092
rect 21315 22052 23204 22080
rect 21315 22049 21327 22052
rect 21269 22043 21327 22049
rect 23198 22040 23204 22052
rect 23256 22040 23262 22092
rect 9272 21984 14320 22012
rect 9272 21972 9278 21984
rect 14366 21972 14372 22024
rect 14424 22012 14430 22024
rect 14737 22015 14795 22021
rect 14737 22012 14749 22015
rect 14424 21984 14749 22012
rect 14424 21972 14430 21984
rect 14737 21981 14749 21984
rect 14783 22012 14795 22015
rect 15654 22012 15660 22024
rect 14783 21984 15660 22012
rect 14783 21981 14795 21984
rect 14737 21975 14795 21981
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 16758 21972 16764 22024
rect 16816 21972 16822 22024
rect 16868 21984 18092 22012
rect 6362 21944 6368 21956
rect 5842 21916 6368 21944
rect 6362 21904 6368 21916
rect 6420 21944 6426 21956
rect 7466 21944 7472 21956
rect 6420 21916 7472 21944
rect 6420 21904 6426 21916
rect 7466 21904 7472 21916
rect 7524 21944 7530 21956
rect 8478 21944 8484 21956
rect 7524 21916 8484 21944
rect 7524 21904 7530 21916
rect 8478 21904 8484 21916
rect 8536 21904 8542 21956
rect 10778 21904 10784 21956
rect 10836 21944 10842 21956
rect 11790 21944 11796 21956
rect 10836 21916 11796 21944
rect 10836 21904 10842 21916
rect 11790 21904 11796 21916
rect 11848 21904 11854 21956
rect 13265 21947 13323 21953
rect 13265 21913 13277 21947
rect 13311 21944 13323 21947
rect 13311 21916 13584 21944
rect 13311 21913 13323 21916
rect 13265 21907 13323 21913
rect 6089 21879 6147 21885
rect 6089 21845 6101 21879
rect 6135 21876 6147 21879
rect 6270 21876 6276 21888
rect 6135 21848 6276 21876
rect 6135 21845 6147 21848
rect 6089 21839 6147 21845
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 6546 21836 6552 21888
rect 6604 21836 6610 21888
rect 6914 21836 6920 21888
rect 6972 21836 6978 21888
rect 7006 21836 7012 21888
rect 7064 21836 7070 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 9582 21876 9588 21888
rect 8628 21848 9588 21876
rect 8628 21836 8634 21848
rect 9582 21836 9588 21848
rect 9640 21836 9646 21888
rect 12434 21836 12440 21888
rect 12492 21836 12498 21888
rect 12710 21836 12716 21888
rect 12768 21876 12774 21888
rect 12897 21879 12955 21885
rect 12897 21876 12909 21879
rect 12768 21848 12909 21876
rect 12768 21836 12774 21848
rect 12897 21845 12909 21848
rect 12943 21845 12955 21879
rect 12897 21839 12955 21845
rect 13354 21836 13360 21888
rect 13412 21836 13418 21888
rect 13556 21876 13584 21916
rect 13630 21904 13636 21956
rect 13688 21944 13694 21956
rect 15286 21944 15292 21956
rect 13688 21916 15292 21944
rect 13688 21904 13694 21916
rect 15286 21904 15292 21916
rect 15344 21904 15350 21956
rect 15565 21947 15623 21953
rect 15565 21913 15577 21947
rect 15611 21944 15623 21947
rect 16482 21944 16488 21956
rect 15611 21916 16488 21944
rect 15611 21913 15623 21916
rect 15565 21907 15623 21913
rect 13814 21876 13820 21888
rect 13556 21848 13820 21876
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14645 21879 14703 21885
rect 14645 21845 14657 21879
rect 14691 21876 14703 21879
rect 15580 21876 15608 21907
rect 16482 21904 16488 21916
rect 16540 21944 16546 21956
rect 16868 21944 16896 21984
rect 17957 21947 18015 21953
rect 17957 21944 17969 21947
rect 16540 21916 16896 21944
rect 17144 21916 17969 21944
rect 16540 21904 16546 21916
rect 14691 21848 15608 21876
rect 14691 21845 14703 21848
rect 14645 21839 14703 21845
rect 16666 21836 16672 21888
rect 16724 21836 16730 21888
rect 17144 21885 17172 21916
rect 17957 21913 17969 21916
rect 18003 21913 18015 21947
rect 18064 21944 18092 21984
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19889 22015 19947 22021
rect 19889 22012 19901 22015
rect 19484 21984 19901 22012
rect 19484 21972 19490 21984
rect 19889 21981 19901 21984
rect 19935 21981 19947 22015
rect 19889 21975 19947 21981
rect 24946 21972 24952 22024
rect 25004 22012 25010 22024
rect 25225 22015 25283 22021
rect 25225 22012 25237 22015
rect 25004 21984 25237 22012
rect 25004 21972 25010 21984
rect 25225 21981 25237 21984
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 20714 21944 20720 21956
rect 18064 21916 20720 21944
rect 17957 21907 18015 21913
rect 20714 21904 20720 21916
rect 20772 21904 20778 21956
rect 21542 21904 21548 21956
rect 21600 21904 21606 21956
rect 22002 21944 22008 21956
rect 21652 21916 22008 21944
rect 17129 21879 17187 21885
rect 17129 21845 17141 21879
rect 17175 21845 17187 21879
rect 17129 21839 17187 21845
rect 17310 21836 17316 21888
rect 17368 21876 17374 21888
rect 17589 21879 17647 21885
rect 17589 21876 17601 21879
rect 17368 21848 17601 21876
rect 17368 21836 17374 21848
rect 17589 21845 17601 21848
rect 17635 21845 17647 21879
rect 17589 21839 17647 21845
rect 18322 21836 18328 21888
rect 18380 21876 18386 21888
rect 19058 21876 19064 21888
rect 18380 21848 19064 21876
rect 18380 21836 18386 21848
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19521 21879 19579 21885
rect 19521 21876 19533 21879
rect 19484 21848 19533 21876
rect 19484 21836 19490 21848
rect 19521 21845 19533 21848
rect 19567 21876 19579 21879
rect 20898 21876 20904 21888
rect 19567 21848 20904 21876
rect 19567 21845 19579 21848
rect 19521 21839 19579 21845
rect 20898 21836 20904 21848
rect 20956 21876 20962 21888
rect 21652 21876 21680 21916
rect 22002 21904 22008 21916
rect 22060 21904 22066 21956
rect 22830 21904 22836 21956
rect 22888 21944 22894 21956
rect 23661 21947 23719 21953
rect 23661 21944 23673 21947
rect 22888 21916 23673 21944
rect 22888 21904 22894 21916
rect 23661 21913 23673 21916
rect 23707 21913 23719 21947
rect 23661 21907 23719 21913
rect 23845 21947 23903 21953
rect 23845 21913 23857 21947
rect 23891 21944 23903 21947
rect 24302 21944 24308 21956
rect 23891 21916 24308 21944
rect 23891 21913 23903 21916
rect 23845 21907 23903 21913
rect 24302 21904 24308 21916
rect 24360 21904 24366 21956
rect 20956 21848 21680 21876
rect 20956 21836 20962 21848
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 23017 21879 23075 21885
rect 23017 21876 23029 21879
rect 22428 21848 23029 21876
rect 22428 21836 22434 21848
rect 23017 21845 23029 21848
rect 23063 21845 23075 21879
rect 23017 21839 23075 21845
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 24118 21876 24124 21888
rect 23624 21848 24124 21876
rect 23624 21836 23630 21848
rect 24118 21836 24124 21848
rect 24176 21836 24182 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 6362 21632 6368 21684
rect 6420 21632 6426 21684
rect 6914 21632 6920 21684
rect 6972 21672 6978 21684
rect 7469 21675 7527 21681
rect 7469 21672 7481 21675
rect 6972 21644 7481 21672
rect 6972 21632 6978 21644
rect 7469 21641 7481 21644
rect 7515 21641 7527 21675
rect 7469 21635 7527 21641
rect 7834 21632 7840 21684
rect 7892 21672 7898 21684
rect 8665 21675 8723 21681
rect 8665 21672 8677 21675
rect 7892 21644 8677 21672
rect 7892 21632 7898 21644
rect 8665 21641 8677 21644
rect 8711 21641 8723 21675
rect 8665 21635 8723 21641
rect 9033 21675 9091 21681
rect 9033 21641 9045 21675
rect 9079 21672 9091 21675
rect 10318 21672 10324 21684
rect 9079 21644 10324 21672
rect 9079 21641 9091 21644
rect 9033 21635 9091 21641
rect 10318 21632 10324 21644
rect 10376 21632 10382 21684
rect 10428 21644 11284 21672
rect 3326 21604 3332 21616
rect 1964 21576 3332 21604
rect 1964 21545 1992 21576
rect 3326 21564 3332 21576
rect 3384 21564 3390 21616
rect 8294 21564 8300 21616
rect 8352 21604 8358 21616
rect 8352 21576 9260 21604
rect 8352 21564 8358 21576
rect 1949 21539 2007 21545
rect 1949 21505 1961 21539
rect 1995 21505 2007 21539
rect 1949 21499 2007 21505
rect 4246 21496 4252 21548
rect 4304 21496 4310 21548
rect 7837 21539 7895 21545
rect 7837 21505 7849 21539
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 7929 21539 7987 21545
rect 7929 21505 7941 21539
rect 7975 21536 7987 21539
rect 9030 21536 9036 21548
rect 7975 21508 9036 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 2866 21428 2872 21480
rect 2924 21428 2930 21480
rect 4062 21428 4068 21480
rect 4120 21428 4126 21480
rect 7852 21468 7880 21499
rect 9030 21496 9036 21508
rect 9088 21496 9094 21548
rect 8113 21471 8171 21477
rect 7852 21440 7972 21468
rect 7944 21400 7972 21440
rect 8113 21437 8125 21471
rect 8159 21468 8171 21471
rect 8202 21468 8208 21480
rect 8159 21440 8208 21468
rect 8159 21437 8171 21440
rect 8113 21431 8171 21437
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 9232 21477 9260 21576
rect 9582 21564 9588 21616
rect 9640 21604 9646 21616
rect 10428 21604 10456 21644
rect 11146 21604 11152 21616
rect 9640 21576 10456 21604
rect 10704 21576 11152 21604
rect 9640 21564 9646 21576
rect 9125 21471 9183 21477
rect 9125 21437 9137 21471
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 9217 21471 9275 21477
rect 9217 21437 9229 21471
rect 9263 21437 9275 21471
rect 9217 21431 9275 21437
rect 8570 21400 8576 21412
rect 7944 21372 8576 21400
rect 8570 21360 8576 21372
rect 8628 21360 8634 21412
rect 1670 21292 1676 21344
rect 1728 21332 1734 21344
rect 1765 21335 1823 21341
rect 1765 21332 1777 21335
rect 1728 21304 1777 21332
rect 1728 21292 1734 21304
rect 1765 21301 1777 21304
rect 1811 21301 1823 21335
rect 9140 21332 9168 21431
rect 10134 21428 10140 21480
rect 10192 21468 10198 21480
rect 10704 21468 10732 21576
rect 11146 21564 11152 21576
rect 11204 21564 11210 21616
rect 11256 21604 11284 21644
rect 11790 21632 11796 21684
rect 11848 21672 11854 21684
rect 15194 21672 15200 21684
rect 11848 21644 15200 21672
rect 11848 21632 11854 21644
rect 15194 21632 15200 21644
rect 15252 21632 15258 21684
rect 15841 21675 15899 21681
rect 15841 21641 15853 21675
rect 15887 21672 15899 21675
rect 16850 21672 16856 21684
rect 15887 21644 16856 21672
rect 15887 21641 15899 21644
rect 15841 21635 15899 21641
rect 16850 21632 16856 21644
rect 16908 21632 16914 21684
rect 18325 21675 18383 21681
rect 18325 21641 18337 21675
rect 18371 21672 18383 21675
rect 18414 21672 18420 21684
rect 18371 21644 18420 21672
rect 18371 21641 18383 21644
rect 18325 21635 18383 21641
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 19426 21672 19432 21684
rect 18524 21644 19432 21672
rect 12161 21607 12219 21613
rect 12161 21604 12173 21607
rect 11256 21576 12173 21604
rect 12161 21573 12173 21576
rect 12207 21573 12219 21607
rect 12161 21567 12219 21573
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 11606 21536 11612 21548
rect 10827 21508 11612 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 11606 21496 11612 21508
rect 11664 21496 11670 21548
rect 12176 21536 12204 21567
rect 12434 21564 12440 21616
rect 12492 21604 12498 21616
rect 13081 21607 13139 21613
rect 13081 21604 13093 21607
rect 12492 21576 13093 21604
rect 12492 21564 12498 21576
rect 13081 21573 13093 21576
rect 13127 21573 13139 21607
rect 13081 21567 13139 21573
rect 13262 21564 13268 21616
rect 13320 21604 13326 21616
rect 13906 21604 13912 21616
rect 13320 21576 13912 21604
rect 13320 21564 13326 21576
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 15933 21607 15991 21613
rect 15933 21604 15945 21607
rect 14568 21576 15945 21604
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12176 21508 13001 21536
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 14458 21536 14464 21548
rect 12989 21499 13047 21505
rect 13372 21508 14464 21536
rect 10873 21471 10931 21477
rect 10873 21468 10885 21471
rect 10192 21440 10885 21468
rect 10192 21428 10198 21440
rect 10873 21437 10885 21440
rect 10919 21437 10931 21471
rect 10873 21431 10931 21437
rect 10962 21428 10968 21480
rect 11020 21468 11026 21480
rect 12897 21471 12955 21477
rect 11020 21440 12434 21468
rect 11020 21428 11026 21440
rect 11422 21400 11428 21412
rect 9968 21372 11428 21400
rect 9968 21332 9996 21372
rect 11422 21360 11428 21372
rect 11480 21360 11486 21412
rect 12406 21400 12434 21440
rect 12897 21437 12909 21471
rect 12943 21468 12955 21471
rect 13372 21468 13400 21508
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 14568 21468 14596 21576
rect 15933 21573 15945 21576
rect 15979 21573 15991 21607
rect 15933 21567 15991 21573
rect 17494 21564 17500 21616
rect 17552 21604 17558 21616
rect 18524 21604 18552 21644
rect 19426 21632 19432 21644
rect 19484 21672 19490 21684
rect 19702 21672 19708 21684
rect 19484 21644 19708 21672
rect 19484 21632 19490 21644
rect 19702 21632 19708 21644
rect 19760 21632 19766 21684
rect 20898 21632 20904 21684
rect 20956 21672 20962 21684
rect 21453 21675 21511 21681
rect 21453 21672 21465 21675
rect 20956 21644 21465 21672
rect 20956 21632 20962 21644
rect 21453 21641 21465 21644
rect 21499 21641 21511 21675
rect 21453 21635 21511 21641
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22373 21675 22431 21681
rect 22373 21672 22385 21675
rect 22244 21644 22385 21672
rect 22244 21632 22250 21644
rect 22373 21641 22385 21644
rect 22419 21641 22431 21675
rect 22373 21635 22431 21641
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 22554 21672 22560 21684
rect 22511 21644 22560 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 25225 21675 25283 21681
rect 25225 21672 25237 21675
rect 23860 21644 25237 21672
rect 17552 21576 18630 21604
rect 17552 21564 17558 21576
rect 20254 21564 20260 21616
rect 20312 21604 20318 21616
rect 22830 21604 22836 21616
rect 20312 21576 22836 21604
rect 20312 21564 20318 21576
rect 22830 21564 22836 21576
rect 22888 21564 22894 21616
rect 23474 21564 23480 21616
rect 23532 21564 23538 21616
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 23860 21604 23888 21644
rect 25225 21641 25237 21644
rect 25271 21641 25283 21675
rect 25225 21635 25283 21641
rect 23624 21576 23966 21604
rect 23624 21564 23630 21576
rect 14645 21539 14703 21545
rect 14645 21505 14657 21539
rect 14691 21536 14703 21539
rect 14691 21508 14964 21536
rect 14691 21505 14703 21508
rect 14645 21499 14703 21505
rect 12943 21440 13400 21468
rect 13648 21440 14596 21468
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 13262 21400 13268 21412
rect 12406 21372 13268 21400
rect 13262 21360 13268 21372
rect 13320 21360 13326 21412
rect 9140 21304 9996 21332
rect 1765 21295 1823 21301
rect 10134 21292 10140 21344
rect 10192 21292 10198 21344
rect 10410 21292 10416 21344
rect 10468 21292 10474 21344
rect 11606 21292 11612 21344
rect 11664 21292 11670 21344
rect 11790 21292 11796 21344
rect 11848 21292 11854 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 13354 21332 13360 21344
rect 12492 21304 13360 21332
rect 12492 21292 12498 21304
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 13449 21335 13507 21341
rect 13449 21301 13461 21335
rect 13495 21332 13507 21335
rect 13648 21332 13676 21440
rect 14734 21428 14740 21480
rect 14792 21428 14798 21480
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21437 14887 21471
rect 14829 21431 14887 21437
rect 13906 21360 13912 21412
rect 13964 21400 13970 21412
rect 14844 21400 14872 21431
rect 13964 21372 14872 21400
rect 14936 21400 14964 21508
rect 15286 21496 15292 21548
rect 15344 21536 15350 21548
rect 17405 21539 17463 21545
rect 17405 21536 17417 21539
rect 15344 21508 17417 21536
rect 15344 21496 15350 21508
rect 17405 21505 17417 21508
rect 17451 21505 17463 21539
rect 18322 21536 18328 21548
rect 17405 21499 17463 21505
rect 17880 21508 18328 21536
rect 15746 21428 15752 21480
rect 15804 21428 15810 21480
rect 16761 21471 16819 21477
rect 16761 21468 16773 21471
rect 15856 21440 16773 21468
rect 15856 21400 15884 21440
rect 16761 21437 16773 21440
rect 16807 21468 16819 21471
rect 17880 21468 17908 21508
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 20070 21496 20076 21548
rect 20128 21496 20134 21548
rect 20530 21496 20536 21548
rect 20588 21496 20594 21548
rect 22646 21496 22652 21548
rect 22704 21536 22710 21548
rect 23198 21536 23204 21548
rect 22704 21508 23204 21536
rect 22704 21496 22710 21508
rect 23198 21496 23204 21508
rect 23256 21496 23262 21548
rect 16807 21440 17908 21468
rect 16807 21437 16819 21440
rect 16761 21431 16819 21437
rect 17954 21428 17960 21480
rect 18012 21468 18018 21480
rect 18598 21468 18604 21480
rect 18012 21440 18604 21468
rect 18012 21428 18018 21440
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 19797 21471 19855 21477
rect 19797 21437 19809 21471
rect 19843 21468 19855 21471
rect 21177 21471 21235 21477
rect 21177 21468 21189 21471
rect 19843 21440 21189 21468
rect 19843 21437 19855 21440
rect 19797 21431 19855 21437
rect 21177 21437 21189 21440
rect 21223 21437 21235 21471
rect 21177 21431 21235 21437
rect 22557 21471 22615 21477
rect 22557 21437 22569 21471
rect 22603 21437 22615 21471
rect 22557 21431 22615 21437
rect 14936 21372 15884 21400
rect 16301 21403 16359 21409
rect 13964 21360 13970 21372
rect 16301 21369 16313 21403
rect 16347 21400 16359 21403
rect 16347 21372 18828 21400
rect 16347 21369 16359 21372
rect 16301 21363 16359 21369
rect 13495 21304 13676 21332
rect 13495 21301 13507 21304
rect 13449 21295 13507 21301
rect 13814 21292 13820 21344
rect 13872 21292 13878 21344
rect 13998 21292 14004 21344
rect 14056 21292 14062 21344
rect 14274 21292 14280 21344
rect 14332 21292 14338 21344
rect 16850 21292 16856 21344
rect 16908 21332 16914 21344
rect 17494 21332 17500 21344
rect 16908 21304 17500 21332
rect 16908 21292 16914 21304
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 17589 21335 17647 21341
rect 17589 21301 17601 21335
rect 17635 21332 17647 21335
rect 17862 21332 17868 21344
rect 17635 21304 17868 21332
rect 17635 21301 17647 21304
rect 17589 21295 17647 21301
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 18800 21332 18828 21372
rect 19242 21332 19248 21344
rect 18800 21304 19248 21332
rect 19242 21292 19248 21304
rect 19300 21292 19306 21344
rect 21634 21292 21640 21344
rect 21692 21332 21698 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21692 21304 22017 21332
rect 21692 21292 21698 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22572 21332 22600 21431
rect 24946 21332 24952 21344
rect 22572 21304 24952 21332
rect 22005 21295 22063 21301
rect 24946 21292 24952 21304
rect 25004 21292 25010 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 7098 21088 7104 21140
rect 7156 21088 7162 21140
rect 8478 21088 8484 21140
rect 8536 21128 8542 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8536 21100 8953 21128
rect 8536 21088 8542 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 9306 21088 9312 21140
rect 9364 21128 9370 21140
rect 9364 21100 10732 21128
rect 9364 21088 9370 21100
rect 1302 20952 1308 21004
rect 1360 20992 1366 21004
rect 2041 20995 2099 21001
rect 2041 20992 2053 20995
rect 1360 20964 2053 20992
rect 1360 20952 1366 20964
rect 2041 20961 2053 20964
rect 2087 20961 2099 20995
rect 2041 20955 2099 20961
rect 5350 20952 5356 21004
rect 5408 20952 5414 21004
rect 8386 20952 8392 21004
rect 8444 20992 8450 21004
rect 9401 20995 9459 21001
rect 9401 20992 9413 20995
rect 8444 20964 9413 20992
rect 8444 20952 8450 20964
rect 9401 20961 9413 20964
rect 9447 20961 9459 20995
rect 9401 20955 9459 20961
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9766 20992 9772 21004
rect 9723 20964 9772 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 10134 20952 10140 21004
rect 10192 20992 10198 21004
rect 10410 20992 10416 21004
rect 10192 20964 10416 20992
rect 10192 20952 10198 20964
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 10704 20992 10732 21100
rect 11606 21088 11612 21140
rect 11664 21128 11670 21140
rect 15286 21128 15292 21140
rect 11664 21100 15292 21128
rect 11664 21088 11670 21100
rect 15286 21088 15292 21100
rect 15344 21128 15350 21140
rect 15344 21100 15700 21128
rect 15344 21088 15350 21100
rect 15672 21060 15700 21100
rect 15746 21088 15752 21140
rect 15804 21128 15810 21140
rect 16025 21131 16083 21137
rect 16025 21128 16037 21131
rect 15804 21100 16037 21128
rect 15804 21088 15810 21100
rect 16025 21097 16037 21100
rect 16071 21097 16083 21131
rect 16025 21091 16083 21097
rect 15930 21060 15936 21072
rect 15672 21032 15936 21060
rect 15930 21020 15936 21032
rect 15988 21020 15994 21072
rect 12434 20992 12440 21004
rect 10704 20964 12440 20992
rect 12434 20952 12440 20964
rect 12492 20952 12498 21004
rect 12802 20952 12808 21004
rect 12860 20992 12866 21004
rect 14277 20995 14335 21001
rect 14277 20992 14289 20995
rect 12860 20964 14289 20992
rect 12860 20952 12866 20964
rect 14277 20961 14289 20964
rect 14323 20961 14335 20995
rect 14277 20955 14335 20961
rect 1762 20884 1768 20936
rect 1820 20884 1826 20936
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7156 20896 7573 20924
rect 7156 20884 7162 20896
rect 7561 20893 7573 20896
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 8570 20884 8576 20936
rect 8628 20924 8634 20936
rect 8938 20924 8944 20936
rect 8628 20896 8944 20924
rect 8628 20884 8634 20896
rect 8938 20884 8944 20896
rect 8996 20924 9002 20936
rect 9306 20924 9312 20936
rect 8996 20896 9312 20924
rect 8996 20884 9002 20896
rect 9306 20884 9312 20896
rect 9364 20884 9370 20936
rect 11238 20924 11244 20936
rect 10810 20910 11244 20924
rect 10796 20896 11244 20910
rect 5626 20816 5632 20868
rect 5684 20816 5690 20868
rect 6362 20816 6368 20868
rect 6420 20816 6426 20868
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 8536 20828 10166 20856
rect 8536 20816 8542 20828
rect 7834 20748 7840 20800
rect 7892 20788 7898 20800
rect 8205 20791 8263 20797
rect 8205 20788 8217 20791
rect 7892 20760 8217 20788
rect 7892 20748 7898 20760
rect 8205 20757 8217 20760
rect 8251 20757 8263 20791
rect 8205 20751 8263 20757
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 8757 20791 8815 20797
rect 8757 20788 8769 20791
rect 8720 20760 8769 20788
rect 8720 20748 8726 20760
rect 8757 20757 8769 20760
rect 8803 20788 8815 20791
rect 8938 20788 8944 20800
rect 8803 20760 8944 20788
rect 8803 20757 8815 20760
rect 8757 20751 8815 20757
rect 8938 20748 8944 20760
rect 8996 20788 9002 20800
rect 9582 20788 9588 20800
rect 8996 20760 9588 20788
rect 8996 20748 9002 20760
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 10060 20788 10088 20828
rect 10796 20788 10824 20896
rect 11238 20884 11244 20896
rect 11296 20924 11302 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11296 20896 11529 20924
rect 11296 20884 11302 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 11517 20887 11575 20893
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 12989 20927 13047 20933
rect 12989 20924 13001 20927
rect 12676 20896 13001 20924
rect 12676 20884 12682 20896
rect 12989 20893 13001 20896
rect 13035 20893 13047 20927
rect 16040 20924 16068 21091
rect 18506 21088 18512 21140
rect 18564 21128 18570 21140
rect 18877 21131 18935 21137
rect 18877 21128 18889 21131
rect 18564 21100 18889 21128
rect 18564 21088 18570 21100
rect 18877 21097 18889 21100
rect 18923 21097 18935 21131
rect 18877 21091 18935 21097
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 22097 21131 22155 21137
rect 22097 21128 22109 21131
rect 22060 21100 22109 21128
rect 22060 21088 22066 21100
rect 22097 21097 22109 21100
rect 22143 21128 22155 21131
rect 23566 21128 23572 21140
rect 22143 21100 23572 21128
rect 22143 21097 22155 21100
rect 22097 21091 22155 21097
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 18417 21063 18475 21069
rect 18417 21029 18429 21063
rect 18463 21060 18475 21063
rect 19518 21060 19524 21072
rect 18463 21032 19524 21060
rect 18463 21029 18475 21032
rect 18417 21023 18475 21029
rect 19518 21020 19524 21032
rect 19576 21020 19582 21072
rect 17865 20995 17923 21001
rect 17865 20961 17877 20995
rect 17911 20961 17923 20995
rect 17865 20955 17923 20961
rect 16485 20927 16543 20933
rect 16485 20924 16497 20927
rect 16040 20896 16497 20924
rect 12989 20887 13047 20893
rect 16485 20893 16497 20896
rect 16531 20893 16543 20927
rect 17880 20924 17908 20955
rect 17954 20952 17960 21004
rect 18012 20952 18018 21004
rect 18782 20952 18788 21004
rect 18840 20952 18846 21004
rect 20806 20992 20812 21004
rect 18892 20964 20812 20992
rect 18892 20924 18920 20964
rect 20806 20952 20812 20964
rect 20864 20952 20870 21004
rect 21821 20995 21879 21001
rect 21821 20961 21833 20995
rect 21867 20992 21879 20995
rect 22646 20992 22652 21004
rect 21867 20964 22652 20992
rect 21867 20961 21879 20964
rect 21821 20955 21879 20961
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20992 23443 20995
rect 24854 20992 24860 21004
rect 23431 20964 24860 20992
rect 23431 20961 23443 20964
rect 23385 20955 23443 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 17880 20896 18920 20924
rect 24029 20927 24087 20933
rect 16485 20887 16543 20893
rect 24029 20893 24041 20927
rect 24075 20924 24087 20927
rect 24486 20924 24492 20936
rect 24075 20896 24492 20924
rect 24075 20893 24087 20896
rect 24029 20887 24087 20893
rect 24486 20884 24492 20896
rect 24544 20884 24550 20936
rect 14458 20816 14464 20868
rect 14516 20856 14522 20868
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 14516 20828 14565 20856
rect 14516 20816 14522 20828
rect 14553 20825 14565 20828
rect 14599 20825 14611 20859
rect 16850 20856 16856 20868
rect 15778 20828 16856 20856
rect 14553 20819 14611 20825
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 18049 20859 18107 20865
rect 18049 20825 18061 20859
rect 18095 20856 18107 20859
rect 19429 20859 19487 20865
rect 19429 20856 19441 20859
rect 18095 20828 19441 20856
rect 18095 20825 18107 20828
rect 18049 20819 18107 20825
rect 19429 20825 19441 20828
rect 19475 20825 19487 20859
rect 19429 20819 19487 20825
rect 19702 20816 19708 20868
rect 19760 20856 19766 20868
rect 20162 20856 20168 20868
rect 19760 20828 20168 20856
rect 19760 20816 19766 20828
rect 20162 20816 20168 20828
rect 20220 20856 20226 20868
rect 21545 20859 21603 20865
rect 20220 20828 20378 20856
rect 20220 20816 20226 20828
rect 21545 20825 21557 20859
rect 21591 20856 21603 20859
rect 25222 20856 25228 20868
rect 21591 20828 25228 20856
rect 21591 20825 21603 20828
rect 21545 20819 21603 20825
rect 25222 20816 25228 20828
rect 25280 20816 25286 20868
rect 10060 20760 10824 20788
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11149 20791 11207 20797
rect 11149 20788 11161 20791
rect 11020 20760 11161 20788
rect 11020 20748 11026 20760
rect 11149 20757 11161 20760
rect 11195 20757 11207 20791
rect 11149 20751 11207 20757
rect 11698 20748 11704 20800
rect 11756 20748 11762 20800
rect 12526 20748 12532 20800
rect 12584 20788 12590 20800
rect 12805 20791 12863 20797
rect 12805 20788 12817 20791
rect 12584 20760 12817 20788
rect 12584 20748 12590 20760
rect 12805 20757 12817 20760
rect 12851 20757 12863 20791
rect 12805 20751 12863 20757
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 16942 20788 16948 20800
rect 13872 20760 16948 20788
rect 13872 20748 13878 20760
rect 16942 20748 16948 20760
rect 17000 20748 17006 20800
rect 17126 20748 17132 20800
rect 17184 20748 17190 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 20073 20791 20131 20797
rect 20073 20788 20085 20791
rect 19392 20760 20085 20788
rect 19392 20748 19398 20760
rect 20073 20757 20085 20760
rect 20119 20757 20131 20791
rect 20073 20751 20131 20757
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 3418 20544 3424 20596
rect 3476 20584 3482 20596
rect 3697 20587 3755 20593
rect 3697 20584 3709 20587
rect 3476 20556 3709 20584
rect 3476 20544 3482 20556
rect 3697 20553 3709 20556
rect 3743 20553 3755 20587
rect 3697 20547 3755 20553
rect 4338 20544 4344 20596
rect 4396 20544 4402 20596
rect 8846 20544 8852 20596
rect 8904 20544 8910 20596
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 10413 20587 10471 20593
rect 10413 20584 10425 20587
rect 10376 20556 10425 20584
rect 10376 20544 10382 20556
rect 10413 20553 10425 20556
rect 10459 20553 10471 20587
rect 10413 20547 10471 20553
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 11054 20584 11060 20596
rect 10827 20556 11060 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 11698 20544 11704 20596
rect 11756 20584 11762 20596
rect 12161 20587 12219 20593
rect 12161 20584 12173 20587
rect 11756 20556 12173 20584
rect 11756 20544 11762 20556
rect 12161 20553 12173 20556
rect 12207 20553 12219 20587
rect 12161 20547 12219 20553
rect 14458 20544 14464 20596
rect 14516 20584 14522 20596
rect 14734 20584 14740 20596
rect 14516 20556 14740 20584
rect 14516 20544 14522 20556
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 15105 20587 15163 20593
rect 15105 20553 15117 20587
rect 15151 20584 15163 20587
rect 16482 20584 16488 20596
rect 15151 20556 16488 20584
rect 15151 20553 15163 20556
rect 15105 20547 15163 20553
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 19518 20544 19524 20596
rect 19576 20544 19582 20596
rect 21453 20587 21511 20593
rect 21453 20553 21465 20587
rect 21499 20584 21511 20587
rect 21542 20584 21548 20596
rect 21499 20556 21548 20584
rect 21499 20553 21511 20556
rect 21453 20547 21511 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 6362 20476 6368 20528
rect 6420 20516 6426 20528
rect 6420 20488 6854 20516
rect 6420 20476 6426 20488
rect 11974 20476 11980 20528
rect 12032 20516 12038 20528
rect 12032 20488 12296 20516
rect 12032 20476 12038 20488
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20417 3939 20451
rect 3881 20411 3939 20417
rect 4525 20451 4583 20457
rect 4525 20417 4537 20451
rect 4571 20448 4583 20451
rect 6730 20448 6736 20460
rect 4571 20420 6736 20448
rect 4571 20417 4583 20420
rect 4525 20411 4583 20417
rect 3896 20380 3924 20411
rect 6730 20408 6736 20420
rect 6788 20408 6794 20460
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20448 8355 20451
rect 8386 20448 8392 20460
rect 8343 20420 8392 20448
rect 8343 20417 8355 20420
rect 8297 20411 8355 20417
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8938 20408 8944 20460
rect 8996 20448 9002 20460
rect 9217 20451 9275 20457
rect 9217 20448 9229 20451
rect 8996 20420 9229 20448
rect 8996 20408 9002 20420
rect 9217 20417 9229 20420
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 12268 20448 12296 20488
rect 14090 20476 14096 20528
rect 14148 20516 14154 20528
rect 18417 20519 18475 20525
rect 14148 20488 16068 20516
rect 14148 20476 14154 20488
rect 14550 20448 14556 20460
rect 12268 20420 14556 20448
rect 5994 20380 6000 20392
rect 3896 20352 6000 20380
rect 5994 20340 6000 20352
rect 6052 20340 6058 20392
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 9122 20380 9128 20392
rect 8067 20352 9128 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 9122 20340 9128 20352
rect 9180 20340 9186 20392
rect 9306 20340 9312 20392
rect 9364 20340 9370 20392
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20349 9551 20383
rect 9493 20343 9551 20349
rect 9508 20312 9536 20343
rect 10870 20340 10876 20392
rect 10928 20340 10934 20392
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 9674 20312 9680 20324
rect 9508 20284 9680 20312
rect 9674 20272 9680 20284
rect 9732 20312 9738 20324
rect 10980 20312 11008 20340
rect 9732 20284 11008 20312
rect 12084 20312 12112 20411
rect 12268 20389 12296 20420
rect 14550 20408 14556 20420
rect 14608 20448 14614 20460
rect 16040 20457 16068 20488
rect 18417 20485 18429 20519
rect 18463 20516 18475 20519
rect 18506 20516 18512 20528
rect 18463 20488 18512 20516
rect 18463 20485 18475 20488
rect 18417 20479 18475 20485
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 19429 20519 19487 20525
rect 19429 20485 19441 20519
rect 19475 20516 19487 20519
rect 19978 20516 19984 20528
rect 19475 20488 19984 20516
rect 19475 20485 19487 20488
rect 19429 20479 19487 20485
rect 19978 20476 19984 20488
rect 20036 20476 20042 20528
rect 16025 20451 16083 20457
rect 14608 20420 15332 20448
rect 14608 20408 14614 20420
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 14461 20383 14519 20389
rect 14461 20349 14473 20383
rect 14507 20380 14519 20383
rect 15010 20380 15016 20392
rect 14507 20352 15016 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 15010 20340 15016 20352
rect 15068 20380 15074 20392
rect 15304 20389 15332 20420
rect 16025 20417 16037 20451
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 18782 20448 18788 20460
rect 17727 20420 18788 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 19352 20420 20821 20448
rect 19352 20392 19380 20420
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 22278 20408 22284 20460
rect 22336 20408 22342 20460
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20448 23351 20451
rect 24854 20448 24860 20460
rect 23339 20420 24860 20448
rect 23339 20417 23351 20420
rect 23293 20411 23351 20417
rect 24854 20408 24860 20420
rect 24912 20408 24918 20460
rect 25130 20408 25136 20460
rect 25188 20408 25194 20460
rect 15197 20383 15255 20389
rect 15197 20380 15209 20383
rect 15068 20352 15209 20380
rect 15068 20340 15074 20352
rect 15197 20349 15209 20352
rect 15243 20349 15255 20383
rect 15197 20343 15255 20349
rect 15289 20383 15347 20389
rect 15289 20349 15301 20383
rect 15335 20349 15347 20383
rect 15289 20343 15347 20349
rect 16224 20352 19288 20380
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 12084 20284 12817 20312
rect 9732 20272 9738 20284
rect 12805 20281 12817 20284
rect 12851 20312 12863 20315
rect 15746 20312 15752 20324
rect 12851 20284 15752 20312
rect 12851 20281 12863 20284
rect 12805 20275 12863 20281
rect 15746 20272 15752 20284
rect 15804 20272 15810 20324
rect 16224 20321 16252 20352
rect 16209 20315 16267 20321
rect 16209 20281 16221 20315
rect 16255 20281 16267 20315
rect 16209 20275 16267 20281
rect 18598 20272 18604 20324
rect 18656 20272 18662 20324
rect 19260 20312 19288 20352
rect 19334 20340 19340 20392
rect 19392 20340 19398 20392
rect 24762 20340 24768 20392
rect 24820 20340 24826 20392
rect 21266 20312 21272 20324
rect 19260 20284 21272 20312
rect 21266 20272 21272 20284
rect 21324 20272 21330 20324
rect 6549 20247 6607 20253
rect 6549 20213 6561 20247
rect 6595 20244 6607 20247
rect 6914 20244 6920 20256
rect 6595 20216 6920 20244
rect 6595 20213 6607 20216
rect 6549 20207 6607 20213
rect 6914 20204 6920 20216
rect 6972 20204 6978 20256
rect 9953 20247 10011 20253
rect 9953 20213 9965 20247
rect 9999 20244 10011 20247
rect 10502 20244 10508 20256
rect 9999 20216 10508 20244
rect 9999 20213 10011 20216
rect 9953 20207 10011 20213
rect 10502 20204 10508 20216
rect 10560 20204 10566 20256
rect 10594 20204 10600 20256
rect 10652 20244 10658 20256
rect 11701 20247 11759 20253
rect 11701 20244 11713 20247
rect 10652 20216 11713 20244
rect 10652 20204 10658 20216
rect 11701 20213 11713 20216
rect 11747 20213 11759 20247
rect 11701 20207 11759 20213
rect 14734 20204 14740 20256
rect 14792 20204 14798 20256
rect 16853 20247 16911 20253
rect 16853 20213 16865 20247
rect 16899 20244 16911 20247
rect 16942 20244 16948 20256
rect 16899 20216 16948 20244
rect 16899 20213 16911 20216
rect 16853 20207 16911 20213
rect 16942 20204 16948 20216
rect 17000 20204 17006 20256
rect 17678 20204 17684 20256
rect 17736 20244 17742 20256
rect 17773 20247 17831 20253
rect 17773 20244 17785 20247
rect 17736 20216 17785 20244
rect 17736 20204 17742 20216
rect 17773 20213 17785 20216
rect 17819 20213 17831 20247
rect 17773 20207 17831 20213
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 19889 20247 19947 20253
rect 19889 20244 19901 20247
rect 19668 20216 19901 20244
rect 19668 20204 19674 20216
rect 19889 20213 19901 20216
rect 19935 20213 19947 20247
rect 19889 20207 19947 20213
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 5626 20000 5632 20052
rect 5684 20040 5690 20052
rect 6089 20043 6147 20049
rect 6089 20040 6101 20043
rect 5684 20012 6101 20040
rect 5684 20000 5690 20012
rect 6089 20009 6101 20012
rect 6135 20009 6147 20043
rect 6089 20003 6147 20009
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 7064 20012 7849 20040
rect 7064 20000 7070 20012
rect 7837 20009 7849 20012
rect 7883 20009 7895 20043
rect 7837 20003 7895 20009
rect 9030 20000 9036 20052
rect 9088 20040 9094 20052
rect 10045 20043 10103 20049
rect 10045 20040 10057 20043
rect 9088 20012 10057 20040
rect 9088 20000 9094 20012
rect 10045 20009 10057 20012
rect 10091 20009 10103 20043
rect 11698 20040 11704 20052
rect 10045 20003 10103 20009
rect 11164 20012 11704 20040
rect 5166 19932 5172 19984
rect 5224 19972 5230 19984
rect 11164 19972 11192 20012
rect 11698 20000 11704 20012
rect 11756 20000 11762 20052
rect 14277 20043 14335 20049
rect 14277 20009 14289 20043
rect 14323 20040 14335 20043
rect 14642 20040 14648 20052
rect 14323 20012 14648 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20040 17003 20043
rect 20990 20040 20996 20052
rect 16991 20012 20996 20040
rect 16991 20009 17003 20012
rect 16945 20003 17003 20009
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 23566 20000 23572 20052
rect 23624 20040 23630 20052
rect 24397 20043 24455 20049
rect 24397 20040 24409 20043
rect 23624 20012 24409 20040
rect 23624 20000 23630 20012
rect 24397 20009 24409 20012
rect 24443 20009 24455 20043
rect 24397 20003 24455 20009
rect 5224 19944 11192 19972
rect 5224 19932 5230 19944
rect 11238 19932 11244 19984
rect 11296 19972 11302 19984
rect 16393 19975 16451 19981
rect 11296 19944 12434 19972
rect 11296 19932 11302 19944
rect 8202 19864 8208 19916
rect 8260 19904 8266 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 8260 19876 8401 19904
rect 8260 19864 8266 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 10226 19864 10232 19916
rect 10284 19904 10290 19916
rect 10597 19907 10655 19913
rect 10597 19904 10609 19907
rect 10284 19876 10609 19904
rect 10284 19864 10290 19876
rect 10597 19873 10609 19876
rect 10643 19904 10655 19907
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 10643 19876 11897 19904
rect 10643 19873 10655 19876
rect 10597 19867 10655 19873
rect 11885 19873 11897 19876
rect 11931 19873 11943 19907
rect 12406 19904 12434 19944
rect 16393 19941 16405 19975
rect 16439 19972 16451 19975
rect 16482 19972 16488 19984
rect 16439 19944 16488 19972
rect 16439 19941 16451 19944
rect 16393 19935 16451 19941
rect 16482 19932 16488 19944
rect 16540 19932 16546 19984
rect 18049 19975 18107 19981
rect 18049 19941 18061 19975
rect 18095 19972 18107 19975
rect 18874 19972 18880 19984
rect 18095 19944 18880 19972
rect 18095 19941 18107 19944
rect 18049 19935 18107 19941
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 15102 19904 15108 19916
rect 12406 19876 15108 19904
rect 11885 19867 11943 19873
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 18322 19904 18328 19916
rect 16071 19876 18328 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 19794 19904 19800 19916
rect 18800 19876 19800 19904
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 6914 19836 6920 19848
rect 6779 19808 6920 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6914 19796 6920 19808
rect 6972 19836 6978 19848
rect 8220 19836 8248 19864
rect 6972 19808 8248 19836
rect 10413 19839 10471 19845
rect 6972 19796 6978 19808
rect 10413 19805 10425 19839
rect 10459 19836 10471 19839
rect 10502 19836 10508 19848
rect 10459 19808 10508 19836
rect 10459 19805 10471 19808
rect 10413 19799 10471 19805
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19836 11759 19839
rect 12710 19836 12716 19848
rect 11747 19808 12716 19836
rect 11747 19805 11759 19808
rect 11701 19799 11759 19805
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 16574 19796 16580 19848
rect 16632 19836 16638 19848
rect 16761 19839 16819 19845
rect 16761 19836 16773 19839
rect 16632 19808 16773 19836
rect 16632 19796 16638 19808
rect 16761 19805 16773 19808
rect 16807 19805 16819 19839
rect 16761 19799 16819 19805
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19836 18291 19839
rect 18800 19836 18828 19876
rect 19794 19864 19800 19876
rect 19852 19864 19858 19916
rect 23385 19907 23443 19913
rect 23385 19873 23397 19907
rect 23431 19904 23443 19907
rect 24854 19904 24860 19916
rect 23431 19876 24860 19904
rect 23431 19873 23443 19876
rect 23385 19867 23443 19873
rect 24854 19864 24860 19876
rect 24912 19864 24918 19916
rect 18279 19808 18828 19836
rect 18877 19839 18935 19845
rect 18279 19805 18291 19808
rect 18233 19799 18291 19805
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19150 19836 19156 19848
rect 18923 19808 19156 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19150 19796 19156 19808
rect 19208 19796 19214 19848
rect 21910 19796 21916 19848
rect 21968 19836 21974 19848
rect 22005 19839 22063 19845
rect 22005 19836 22017 19839
rect 21968 19808 22017 19836
rect 21968 19796 21974 19808
rect 22005 19805 22017 19808
rect 22051 19805 22063 19839
rect 22005 19799 22063 19805
rect 23750 19796 23756 19848
rect 23808 19836 23814 19848
rect 23845 19839 23903 19845
rect 23845 19836 23857 19839
rect 23808 19808 23857 19836
rect 23808 19796 23814 19808
rect 23845 19805 23857 19808
rect 23891 19805 23903 19839
rect 23845 19799 23903 19805
rect 24394 19796 24400 19848
rect 24452 19836 24458 19848
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 24452 19808 24593 19836
rect 24452 19796 24458 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 8205 19771 8263 19777
rect 8205 19737 8217 19771
rect 8251 19768 8263 19771
rect 13538 19768 13544 19780
rect 8251 19740 11376 19768
rect 8251 19737 8263 19740
rect 8205 19731 8263 19737
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 7708 19672 8309 19700
rect 7708 19660 7714 19672
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 8297 19663 8355 19669
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 10502 19660 10508 19712
rect 10560 19660 10566 19712
rect 11348 19709 11376 19740
rect 12728 19740 13544 19768
rect 12728 19712 12756 19740
rect 13538 19728 13544 19740
rect 13596 19728 13602 19780
rect 15102 19728 15108 19780
rect 15160 19728 15166 19780
rect 15749 19771 15807 19777
rect 15749 19737 15761 19771
rect 15795 19768 15807 19771
rect 17126 19768 17132 19780
rect 15795 19740 17132 19768
rect 15795 19737 15807 19740
rect 15749 19731 15807 19737
rect 17126 19728 17132 19740
rect 17184 19728 17190 19780
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 20901 19771 20959 19777
rect 20901 19768 20913 19771
rect 17920 19740 20913 19768
rect 17920 19728 17926 19740
rect 20901 19737 20913 19740
rect 20947 19737 20959 19771
rect 20901 19731 20959 19737
rect 22189 19771 22247 19777
rect 22189 19737 22201 19771
rect 22235 19768 22247 19771
rect 22370 19768 22376 19780
rect 22235 19740 22376 19768
rect 22235 19737 22247 19740
rect 22189 19731 22247 19737
rect 22370 19728 22376 19740
rect 22428 19728 22434 19780
rect 11333 19703 11391 19709
rect 11333 19669 11345 19703
rect 11379 19669 11391 19703
rect 11333 19663 11391 19669
rect 11793 19703 11851 19709
rect 11793 19669 11805 19703
rect 11839 19700 11851 19703
rect 12250 19700 12256 19712
rect 11839 19672 12256 19700
rect 11839 19669 11851 19672
rect 11793 19663 11851 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12621 19703 12679 19709
rect 12621 19669 12633 19703
rect 12667 19700 12679 19703
rect 12710 19700 12716 19712
rect 12667 19672 12716 19700
rect 12667 19669 12679 19672
rect 12621 19663 12679 19669
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 13446 19660 13452 19712
rect 13504 19660 13510 19712
rect 18693 19703 18751 19709
rect 18693 19669 18705 19703
rect 18739 19700 18751 19703
rect 18782 19700 18788 19712
rect 18739 19672 18788 19700
rect 18739 19669 18751 19672
rect 18693 19663 18751 19669
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 20993 19703 21051 19709
rect 20993 19669 21005 19703
rect 21039 19700 21051 19703
rect 22646 19700 22652 19712
rect 21039 19672 22652 19700
rect 21039 19669 21051 19672
rect 20993 19663 21051 19669
rect 22646 19660 22652 19672
rect 22704 19660 22710 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 6641 19499 6699 19505
rect 6641 19496 6653 19499
rect 4120 19468 6653 19496
rect 4120 19456 4126 19468
rect 6641 19465 6653 19468
rect 6687 19465 6699 19499
rect 6641 19459 6699 19465
rect 7742 19456 7748 19508
rect 7800 19496 7806 19508
rect 10045 19499 10103 19505
rect 10045 19496 10057 19499
rect 7800 19468 10057 19496
rect 7800 19456 7806 19468
rect 10045 19465 10057 19468
rect 10091 19465 10103 19499
rect 10045 19459 10103 19465
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10505 19499 10563 19505
rect 10505 19496 10517 19499
rect 10192 19468 10517 19496
rect 10192 19456 10198 19468
rect 10505 19465 10517 19468
rect 10551 19465 10563 19499
rect 10505 19459 10563 19465
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 13541 19499 13599 19505
rect 13541 19496 13553 19499
rect 10928 19468 13553 19496
rect 10928 19456 10934 19468
rect 13541 19465 13553 19468
rect 13587 19465 13599 19499
rect 13541 19459 13599 19465
rect 13909 19499 13967 19505
rect 13909 19465 13921 19499
rect 13955 19496 13967 19499
rect 15194 19496 15200 19508
rect 13955 19468 15200 19496
rect 13955 19465 13967 19468
rect 13909 19459 13967 19465
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 18417 19499 18475 19505
rect 18417 19465 18429 19499
rect 18463 19465 18475 19499
rect 18417 19459 18475 19465
rect 2225 19431 2283 19437
rect 2225 19397 2237 19431
rect 2271 19428 2283 19431
rect 2774 19428 2780 19440
rect 2271 19400 2780 19428
rect 2271 19397 2283 19400
rect 2225 19391 2283 19397
rect 2774 19388 2780 19400
rect 2832 19388 2838 19440
rect 8478 19388 8484 19440
rect 8536 19388 8542 19440
rect 9585 19431 9643 19437
rect 9585 19397 9597 19431
rect 9631 19428 9643 19431
rect 11974 19428 11980 19440
rect 9631 19400 11980 19428
rect 9631 19397 9643 19400
rect 9585 19391 9643 19397
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 12161 19431 12219 19437
rect 12161 19397 12173 19431
rect 12207 19428 12219 19431
rect 12710 19428 12716 19440
rect 12207 19400 12716 19428
rect 12207 19397 12219 19400
rect 12161 19391 12219 19397
rect 12710 19388 12716 19400
rect 12768 19388 12774 19440
rect 13446 19388 13452 19440
rect 13504 19428 13510 19440
rect 14001 19431 14059 19437
rect 14001 19428 14013 19431
rect 13504 19400 14013 19428
rect 13504 19388 13510 19400
rect 14001 19397 14013 19400
rect 14047 19428 14059 19431
rect 14047 19400 15056 19428
rect 14047 19397 14059 19400
rect 14001 19391 14059 19397
rect 7101 19363 7159 19369
rect 7101 19360 7113 19363
rect 6104 19332 7113 19360
rect 5534 19252 5540 19304
rect 5592 19292 5598 19304
rect 6104 19301 6132 19332
rect 7101 19329 7113 19332
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7558 19320 7564 19372
rect 7616 19320 7622 19372
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 10686 19360 10692 19372
rect 10468 19332 10692 19360
rect 10468 19320 10474 19332
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 12069 19363 12127 19369
rect 12069 19329 12081 19363
rect 12115 19360 12127 19363
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12115 19332 12909 19360
rect 12115 19329 12127 19332
rect 12069 19323 12127 19329
rect 12897 19329 12909 19332
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 14516 19332 14841 19360
rect 14516 19320 14522 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 15028 19360 15056 19400
rect 15102 19388 15108 19440
rect 15160 19428 15166 19440
rect 15565 19431 15623 19437
rect 15565 19428 15577 19431
rect 15160 19400 15577 19428
rect 15160 19388 15166 19400
rect 15565 19397 15577 19400
rect 15611 19428 15623 19431
rect 16117 19431 16175 19437
rect 16117 19428 16129 19431
rect 15611 19400 16129 19428
rect 15611 19397 15623 19400
rect 15565 19391 15623 19397
rect 16117 19397 16129 19400
rect 16163 19397 16175 19431
rect 18432 19428 18460 19459
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 19153 19499 19211 19505
rect 19153 19496 19165 19499
rect 19024 19468 19165 19496
rect 19024 19456 19030 19468
rect 19153 19465 19165 19468
rect 19199 19465 19211 19499
rect 19153 19459 19211 19465
rect 19058 19428 19064 19440
rect 18432 19400 19064 19428
rect 16117 19391 16175 19397
rect 19058 19388 19064 19400
rect 19116 19388 19122 19440
rect 20162 19388 20168 19440
rect 20220 19428 20226 19440
rect 21177 19431 21235 19437
rect 21177 19428 21189 19431
rect 20220 19400 21189 19428
rect 20220 19388 20226 19400
rect 21177 19397 21189 19400
rect 21223 19397 21235 19431
rect 23566 19428 23572 19440
rect 23506 19400 23572 19428
rect 21177 19391 21235 19397
rect 23566 19388 23572 19400
rect 23624 19428 23630 19440
rect 24118 19428 24124 19440
rect 23624 19400 24124 19428
rect 23624 19388 23630 19400
rect 24118 19388 24124 19400
rect 24176 19428 24182 19440
rect 24949 19431 25007 19437
rect 24949 19428 24961 19431
rect 24176 19400 24961 19428
rect 24176 19388 24182 19400
rect 24949 19397 24961 19400
rect 24995 19397 25007 19431
rect 24949 19391 25007 19397
rect 16666 19360 16672 19372
rect 15028 19332 16672 19360
rect 14829 19323 14887 19329
rect 6089 19295 6147 19301
rect 6089 19292 6101 19295
rect 5592 19264 6101 19292
rect 5592 19252 5598 19264
rect 6089 19261 6101 19264
rect 6135 19261 6147 19295
rect 6089 19255 6147 19261
rect 7834 19252 7840 19304
rect 7892 19252 7898 19304
rect 9398 19252 9404 19304
rect 9456 19292 9462 19304
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 9456 19264 10609 19292
rect 9456 19252 9462 19264
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 10704 19292 10732 19320
rect 11057 19295 11115 19301
rect 11057 19292 11069 19295
rect 10704 19264 11069 19292
rect 10597 19255 10655 19261
rect 11057 19261 11069 19264
rect 11103 19261 11115 19295
rect 11057 19255 11115 19261
rect 11238 19252 11244 19304
rect 11296 19252 11302 19304
rect 12342 19252 12348 19304
rect 12400 19252 12406 19304
rect 14182 19252 14188 19304
rect 14240 19252 14246 19304
rect 14844 19292 14872 19323
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 17402 19320 17408 19372
rect 17460 19360 17466 19372
rect 18233 19363 18291 19369
rect 18233 19360 18245 19363
rect 17460 19332 18245 19360
rect 17460 19320 17466 19332
rect 18233 19329 18245 19332
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 24213 19363 24271 19369
rect 24213 19329 24225 19363
rect 24259 19360 24271 19363
rect 24394 19360 24400 19372
rect 24259 19332 24400 19360
rect 24259 19329 24271 19332
rect 24213 19323 24271 19329
rect 24394 19320 24400 19332
rect 24452 19320 24458 19372
rect 16114 19292 16120 19304
rect 14844 19264 16120 19292
rect 16114 19252 16120 19264
rect 16172 19292 16178 19304
rect 16301 19295 16359 19301
rect 16301 19292 16313 19295
rect 16172 19264 16313 19292
rect 16172 19252 16178 19264
rect 16301 19261 16313 19264
rect 16347 19261 16359 19295
rect 16301 19255 16359 19261
rect 20625 19295 20683 19301
rect 20625 19261 20637 19295
rect 20671 19292 20683 19295
rect 20901 19295 20959 19301
rect 20671 19264 20852 19292
rect 20671 19261 20683 19264
rect 20625 19255 20683 19261
rect 1762 19184 1768 19236
rect 1820 19224 1826 19236
rect 2041 19227 2099 19233
rect 2041 19224 2053 19227
rect 1820 19196 2053 19224
rect 1820 19184 1826 19196
rect 2041 19193 2053 19196
rect 2087 19193 2099 19227
rect 20824 19224 20852 19264
rect 20901 19261 20913 19295
rect 20947 19292 20959 19295
rect 21082 19292 21088 19304
rect 20947 19264 21088 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 21082 19252 21088 19264
rect 21140 19292 21146 19304
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21140 19264 22017 19292
rect 21140 19252 21146 19264
rect 22005 19261 22017 19264
rect 22051 19261 22063 19295
rect 22005 19255 22063 19261
rect 22278 19252 22284 19304
rect 22336 19252 22342 19304
rect 21450 19224 21456 19236
rect 20824 19196 21456 19224
rect 2041 19187 2099 19193
rect 21450 19184 21456 19196
rect 21508 19184 21514 19236
rect 7009 19159 7067 19165
rect 7009 19125 7021 19159
rect 7055 19156 7067 19159
rect 7098 19156 7104 19168
rect 7055 19128 7104 19156
rect 7055 19125 7067 19128
rect 7009 19119 7067 19125
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 11606 19116 11612 19168
rect 11664 19156 11670 19168
rect 11701 19159 11759 19165
rect 11701 19156 11713 19159
rect 11664 19128 11713 19156
rect 11664 19116 11670 19128
rect 11701 19125 11713 19128
rect 11747 19125 11759 19159
rect 11701 19119 11759 19125
rect 16482 19116 16488 19168
rect 16540 19156 16546 19168
rect 18690 19156 18696 19168
rect 16540 19128 18696 19156
rect 16540 19116 16546 19128
rect 18690 19116 18696 19128
rect 18748 19156 18754 19168
rect 20438 19156 20444 19168
rect 18748 19128 20444 19156
rect 18748 19116 18754 19128
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 23750 19116 23756 19168
rect 23808 19116 23814 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 5994 18912 6000 18964
rect 6052 18912 6058 18964
rect 9122 18912 9128 18964
rect 9180 18912 9186 18964
rect 10229 18955 10287 18961
rect 10229 18921 10241 18955
rect 10275 18952 10287 18955
rect 10502 18952 10508 18964
rect 10275 18924 10508 18952
rect 10275 18921 10287 18924
rect 10229 18915 10287 18921
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 11422 18912 11428 18964
rect 11480 18912 11486 18964
rect 15194 18912 15200 18964
rect 15252 18952 15258 18964
rect 15289 18955 15347 18961
rect 15289 18952 15301 18955
rect 15252 18924 15301 18952
rect 15252 18912 15258 18924
rect 15289 18921 15301 18924
rect 15335 18952 15347 18955
rect 16482 18952 16488 18964
rect 15335 18924 16488 18952
rect 15335 18921 15347 18924
rect 15289 18915 15347 18921
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 16666 18912 16672 18964
rect 16724 18912 16730 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19484 18924 20300 18952
rect 19484 18912 19490 18924
rect 6270 18844 6276 18896
rect 6328 18884 6334 18896
rect 6328 18856 7972 18884
rect 6328 18844 6334 18856
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1360 18788 2053 18816
rect 1360 18776 1366 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 6638 18776 6644 18828
rect 6696 18776 6702 18828
rect 1670 18708 1676 18760
rect 1728 18708 1734 18760
rect 7944 18757 7972 18856
rect 10686 18844 10692 18896
rect 10744 18884 10750 18896
rect 12621 18887 12679 18893
rect 12621 18884 12633 18887
rect 10744 18856 12633 18884
rect 10744 18844 10750 18856
rect 12621 18853 12633 18856
rect 12667 18853 12679 18887
rect 12621 18847 12679 18853
rect 13630 18844 13636 18896
rect 13688 18884 13694 18896
rect 16206 18884 16212 18896
rect 13688 18856 16212 18884
rect 13688 18844 13694 18856
rect 16206 18844 16212 18856
rect 16264 18844 16270 18896
rect 17773 18887 17831 18893
rect 17773 18853 17785 18887
rect 17819 18884 17831 18887
rect 19886 18884 19892 18896
rect 17819 18856 19892 18884
rect 17819 18853 17831 18856
rect 17773 18847 17831 18853
rect 19886 18844 19892 18856
rect 19944 18844 19950 18896
rect 20272 18884 20300 18924
rect 20346 18912 20352 18964
rect 20404 18952 20410 18964
rect 21729 18955 21787 18961
rect 21729 18952 21741 18955
rect 20404 18924 21741 18952
rect 20404 18912 20410 18924
rect 21729 18921 21741 18924
rect 21775 18921 21787 18955
rect 21729 18915 21787 18921
rect 22278 18912 22284 18964
rect 22336 18912 22342 18964
rect 21545 18887 21603 18893
rect 21545 18884 21557 18887
rect 20272 18856 21557 18884
rect 21545 18853 21557 18856
rect 21591 18853 21603 18887
rect 21545 18847 21603 18853
rect 10502 18776 10508 18828
rect 10560 18816 10566 18828
rect 10781 18819 10839 18825
rect 10781 18816 10793 18819
rect 10560 18788 10793 18816
rect 10560 18776 10566 18788
rect 10781 18785 10793 18788
rect 10827 18785 10839 18819
rect 10781 18779 10839 18785
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11112 18788 11989 18816
rect 11112 18776 11118 18788
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 11977 18779 12035 18785
rect 12342 18776 12348 18828
rect 12400 18816 12406 18828
rect 13173 18819 13231 18825
rect 13173 18816 13185 18819
rect 12400 18788 13185 18816
rect 12400 18776 12406 18788
rect 13173 18785 13185 18788
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 14642 18776 14648 18828
rect 14700 18816 14706 18828
rect 14700 18788 14964 18816
rect 14700 18776 14706 18788
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18748 6515 18751
rect 7929 18751 7987 18757
rect 6503 18720 7880 18748
rect 6503 18717 6515 18720
rect 6457 18711 6515 18717
rect 6365 18683 6423 18689
rect 6365 18649 6377 18683
rect 6411 18680 6423 18683
rect 7282 18680 7288 18692
rect 6411 18652 7288 18680
rect 6411 18649 6423 18652
rect 6365 18643 6423 18649
rect 7282 18640 7288 18652
rect 7340 18640 7346 18692
rect 7852 18680 7880 18720
rect 7929 18717 7941 18751
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 10226 18748 10232 18760
rect 9824 18720 10232 18748
rect 9824 18708 9830 18720
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18748 10655 18751
rect 13081 18751 13139 18757
rect 10643 18720 12434 18748
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 8846 18680 8852 18692
rect 7852 18652 8852 18680
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 9490 18640 9496 18692
rect 9548 18680 9554 18692
rect 11146 18680 11152 18692
rect 9548 18652 11152 18680
rect 9548 18640 9554 18652
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 11793 18683 11851 18689
rect 11793 18649 11805 18683
rect 11839 18680 11851 18683
rect 12066 18680 12072 18692
rect 11839 18652 12072 18680
rect 11839 18649 11851 18652
rect 11793 18643 11851 18649
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 12406 18680 12434 18720
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 14734 18748 14740 18760
rect 13127 18720 14740 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 14936 18757 14964 18788
rect 17126 18776 17132 18828
rect 17184 18776 17190 18828
rect 17218 18776 17224 18828
rect 17276 18816 17282 18828
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 17276 18788 17325 18816
rect 17276 18776 17282 18788
rect 17313 18785 17325 18788
rect 17359 18816 17371 18819
rect 18049 18819 18107 18825
rect 18049 18816 18061 18819
rect 17359 18788 18061 18816
rect 17359 18785 17371 18788
rect 17313 18779 17371 18785
rect 18049 18785 18061 18788
rect 18095 18785 18107 18819
rect 18049 18779 18107 18785
rect 19613 18819 19671 18825
rect 19613 18785 19625 18819
rect 19659 18816 19671 18819
rect 19702 18816 19708 18828
rect 19659 18788 19708 18816
rect 19659 18785 19671 18788
rect 19613 18779 19671 18785
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 24026 18816 24032 18828
rect 21140 18788 24032 18816
rect 21140 18776 21146 18788
rect 24026 18776 24032 18788
rect 24084 18776 24090 18828
rect 14921 18751 14979 18757
rect 14921 18717 14933 18751
rect 14967 18717 14979 18751
rect 14921 18711 14979 18717
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 16390 18748 16396 18760
rect 16071 18720 16396 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 16666 18708 16672 18760
rect 16724 18748 16730 18760
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 16724 18720 17417 18748
rect 16724 18708 16730 18720
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18748 18383 18751
rect 18690 18748 18696 18760
rect 18371 18720 18696 18748
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19794 18708 19800 18760
rect 19852 18748 19858 18760
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 19852 18720 20637 18748
rect 19852 18708 19858 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 24578 18708 24584 18760
rect 24636 18708 24642 18760
rect 12526 18680 12532 18692
rect 12406 18652 12532 18680
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 13354 18640 13360 18692
rect 13412 18680 13418 18692
rect 14277 18683 14335 18689
rect 14277 18680 14289 18683
rect 13412 18652 14289 18680
rect 13412 18640 13418 18652
rect 14277 18649 14289 18652
rect 14323 18649 14335 18683
rect 14277 18643 14335 18649
rect 18877 18683 18935 18689
rect 18877 18649 18889 18683
rect 18923 18680 18935 18683
rect 20070 18680 20076 18692
rect 18923 18652 20076 18680
rect 18923 18649 18935 18652
rect 18877 18643 18935 18649
rect 20070 18640 20076 18652
rect 20128 18640 20134 18692
rect 23474 18680 23480 18692
rect 23322 18652 23480 18680
rect 23474 18640 23480 18652
rect 23532 18640 23538 18692
rect 23753 18683 23811 18689
rect 23753 18649 23765 18683
rect 23799 18680 23811 18683
rect 25225 18683 25283 18689
rect 25225 18680 25237 18683
rect 23799 18652 25237 18680
rect 23799 18649 23811 18652
rect 23753 18643 23811 18649
rect 25225 18649 25237 18652
rect 25271 18649 25283 18683
rect 25225 18643 25283 18649
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 7156 18584 7205 18612
rect 7156 18572 7162 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 7193 18575 7251 18581
rect 8573 18615 8631 18621
rect 8573 18581 8585 18615
rect 8619 18612 8631 18615
rect 10134 18612 10140 18624
rect 8619 18584 10140 18612
rect 8619 18581 8631 18584
rect 8573 18575 8631 18581
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 10318 18572 10324 18624
rect 10376 18612 10382 18624
rect 10689 18615 10747 18621
rect 10689 18612 10701 18615
rect 10376 18584 10701 18612
rect 10376 18572 10382 18584
rect 10689 18581 10701 18584
rect 10735 18581 10747 18615
rect 10689 18575 10747 18581
rect 11882 18572 11888 18624
rect 11940 18572 11946 18624
rect 12989 18615 13047 18621
rect 12989 18581 13001 18615
rect 13035 18612 13047 18615
rect 13998 18612 14004 18624
rect 13035 18584 14004 18612
rect 13035 18581 13047 18584
rect 12989 18575 13047 18581
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 15930 18572 15936 18624
rect 15988 18572 15994 18624
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 19705 18615 19763 18621
rect 19705 18612 19717 18615
rect 19484 18584 19717 18612
rect 19484 18572 19490 18584
rect 19705 18581 19717 18584
rect 19751 18581 19763 18615
rect 19705 18575 19763 18581
rect 19797 18615 19855 18621
rect 19797 18581 19809 18615
rect 19843 18612 19855 18615
rect 19978 18612 19984 18624
rect 19843 18584 19984 18612
rect 19843 18581 19855 18584
rect 19797 18575 19855 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 20162 18572 20168 18624
rect 20220 18572 20226 18624
rect 21174 18572 21180 18624
rect 21232 18612 21238 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 21232 18584 21281 18612
rect 21232 18572 21238 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 9030 18408 9036 18420
rect 8628 18380 9036 18408
rect 8628 18368 8634 18380
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9125 18411 9183 18417
rect 9125 18377 9137 18411
rect 9171 18408 9183 18411
rect 9766 18408 9772 18420
rect 9171 18380 9772 18408
rect 9171 18377 9183 18380
rect 9125 18371 9183 18377
rect 9766 18368 9772 18380
rect 9824 18408 9830 18420
rect 10870 18408 10876 18420
rect 9824 18380 10876 18408
rect 9824 18368 9830 18380
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 11146 18368 11152 18420
rect 11204 18368 11210 18420
rect 12066 18368 12072 18420
rect 12124 18408 12130 18420
rect 13449 18411 13507 18417
rect 13449 18408 13461 18411
rect 12124 18380 13461 18408
rect 12124 18368 12130 18380
rect 13449 18377 13461 18380
rect 13495 18377 13507 18411
rect 13449 18371 13507 18377
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14461 18411 14519 18417
rect 14461 18408 14473 18411
rect 13872 18380 14473 18408
rect 13872 18368 13878 18380
rect 14461 18377 14473 18380
rect 14507 18408 14519 18411
rect 14642 18408 14648 18420
rect 14507 18380 14648 18408
rect 14507 18377 14519 18380
rect 14461 18371 14519 18377
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 14734 18368 14740 18420
rect 14792 18368 14798 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19978 18408 19984 18420
rect 19392 18380 19984 18408
rect 19392 18368 19398 18380
rect 19978 18368 19984 18380
rect 20036 18408 20042 18420
rect 20073 18411 20131 18417
rect 20073 18408 20085 18411
rect 20036 18380 20085 18408
rect 20036 18368 20042 18380
rect 20073 18377 20085 18380
rect 20119 18377 20131 18411
rect 20073 18371 20131 18377
rect 20898 18368 20904 18420
rect 20956 18408 20962 18420
rect 22373 18411 22431 18417
rect 22373 18408 22385 18411
rect 20956 18380 22385 18408
rect 20956 18368 20962 18380
rect 22373 18377 22385 18380
rect 22419 18377 22431 18411
rect 22373 18371 22431 18377
rect 12161 18343 12219 18349
rect 12161 18309 12173 18343
rect 12207 18340 12219 18343
rect 14274 18340 14280 18352
rect 12207 18312 14280 18340
rect 12207 18309 12219 18312
rect 12161 18303 12219 18309
rect 14274 18300 14280 18312
rect 14332 18300 14338 18352
rect 18322 18340 18328 18352
rect 18064 18312 18328 18340
rect 8478 18272 8484 18284
rect 7958 18244 8484 18272
rect 8478 18232 8484 18244
rect 8536 18272 8542 18284
rect 9490 18272 9496 18284
rect 8536 18244 9496 18272
rect 8536 18232 8542 18244
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 11020 18244 12020 18272
rect 11020 18232 11026 18244
rect 6546 18164 6552 18216
rect 6604 18164 6610 18216
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 7466 18204 7472 18216
rect 6871 18176 7472 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 9858 18204 9864 18216
rect 8619 18176 9864 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 10597 18207 10655 18213
rect 10597 18204 10609 18207
rect 10560 18176 10609 18204
rect 10560 18164 10566 18176
rect 10597 18173 10609 18176
rect 10643 18173 10655 18207
rect 10597 18167 10655 18173
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 11146 18204 11152 18216
rect 10919 18176 11152 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 11992 18204 12020 18244
rect 12066 18232 12072 18284
rect 12124 18232 12130 18284
rect 12176 18244 12434 18272
rect 12176 18204 12204 18244
rect 11992 18176 12204 18204
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 12268 18136 12296 18167
rect 11072 18108 12296 18136
rect 12406 18136 12434 18244
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 15930 18272 15936 18284
rect 13872 18244 15936 18272
rect 13872 18232 13878 18244
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 18064 18281 18092 18312
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 20346 18300 20352 18352
rect 20404 18340 20410 18352
rect 20441 18343 20499 18349
rect 20441 18340 20453 18343
rect 20404 18312 20453 18340
rect 20404 18300 20410 18312
rect 20441 18309 20453 18312
rect 20487 18309 20499 18343
rect 23750 18340 23756 18352
rect 20441 18303 20499 18309
rect 22204 18312 23756 18340
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 20530 18272 20536 18284
rect 19484 18244 20536 18272
rect 19484 18232 19490 18244
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18204 13231 18207
rect 13630 18204 13636 18216
rect 13219 18176 13636 18204
rect 13219 18173 13231 18176
rect 13173 18167 13231 18173
rect 13630 18164 13636 18176
rect 13688 18204 13694 18216
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 13688 18176 13921 18204
rect 13688 18164 13694 18176
rect 13909 18173 13921 18176
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 14093 18207 14151 18213
rect 14093 18173 14105 18207
rect 14139 18204 14151 18207
rect 14182 18204 14188 18216
rect 14139 18176 14188 18204
rect 14139 18173 14151 18176
rect 14093 18167 14151 18173
rect 14108 18136 14136 18167
rect 14182 18164 14188 18176
rect 14240 18164 14246 18216
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 18012 18176 18337 18204
rect 18012 18164 18018 18176
rect 18325 18173 18337 18176
rect 18371 18173 18383 18207
rect 18325 18167 18383 18173
rect 21082 18164 21088 18216
rect 21140 18204 21146 18216
rect 22204 18213 22232 18312
rect 23750 18300 23756 18312
rect 23808 18300 23814 18352
rect 25130 18300 25136 18352
rect 25188 18300 25194 18352
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18272 22339 18275
rect 22738 18272 22744 18284
rect 22327 18244 22744 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 22738 18232 22744 18244
rect 22796 18232 22802 18284
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 21177 18207 21235 18213
rect 21177 18204 21189 18207
rect 21140 18176 21189 18204
rect 21140 18164 21146 18176
rect 21177 18173 21189 18176
rect 21223 18173 21235 18207
rect 21177 18167 21235 18173
rect 22189 18207 22247 18213
rect 22189 18173 22201 18207
rect 22235 18173 22247 18207
rect 22189 18167 22247 18173
rect 12406 18108 14136 18136
rect 9398 18028 9404 18080
rect 9456 18068 9462 18080
rect 11072 18068 11100 18108
rect 20622 18096 20628 18148
rect 20680 18136 20686 18148
rect 23308 18136 23336 18235
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 20680 18108 23336 18136
rect 20680 18096 20686 18108
rect 23474 18096 23480 18148
rect 23532 18096 23538 18148
rect 9456 18040 11100 18068
rect 9456 18028 9462 18040
rect 11698 18028 11704 18080
rect 11756 18028 11762 18080
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 13906 18068 13912 18080
rect 12032 18040 13912 18068
rect 12032 18028 12038 18040
rect 13906 18028 13912 18040
rect 13964 18028 13970 18080
rect 19794 18028 19800 18080
rect 19852 18028 19858 18080
rect 22741 18071 22799 18077
rect 22741 18037 22753 18071
rect 22787 18068 22799 18071
rect 23290 18068 23296 18080
rect 22787 18040 23296 18068
rect 22787 18037 22799 18040
rect 22741 18031 22799 18037
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 5810 17824 5816 17876
rect 5868 17864 5874 17876
rect 5868 17836 6592 17864
rect 5868 17824 5874 17836
rect 6564 17796 6592 17836
rect 6638 17824 6644 17876
rect 6696 17864 6702 17876
rect 6825 17867 6883 17873
rect 6825 17864 6837 17867
rect 6696 17836 6837 17864
rect 6696 17824 6702 17836
rect 6825 17833 6837 17836
rect 6871 17833 6883 17867
rect 6825 17827 6883 17833
rect 7282 17824 7288 17876
rect 7340 17824 7346 17876
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12124 17836 13001 17864
rect 12124 17824 12130 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 17497 17867 17555 17873
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 17954 17864 17960 17876
rect 17543 17836 17960 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 23566 17824 23572 17876
rect 23624 17864 23630 17876
rect 24578 17864 24584 17876
rect 23624 17836 24584 17864
rect 23624 17824 23630 17836
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 10318 17796 10324 17808
rect 6564 17768 10324 17796
rect 10318 17756 10324 17768
rect 10376 17796 10382 17808
rect 10505 17799 10563 17805
rect 10505 17796 10517 17799
rect 10376 17768 10517 17796
rect 10376 17756 10382 17768
rect 10505 17765 10517 17768
rect 10551 17765 10563 17799
rect 10505 17759 10563 17765
rect 12250 17756 12256 17808
rect 12308 17796 12314 17808
rect 14277 17799 14335 17805
rect 14277 17796 14289 17799
rect 12308 17768 14289 17796
rect 12308 17756 12314 17768
rect 14277 17765 14289 17768
rect 14323 17765 14335 17799
rect 14277 17759 14335 17765
rect 14642 17756 14648 17808
rect 14700 17796 14706 17808
rect 14700 17768 14872 17796
rect 14700 17756 14706 17768
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17728 5135 17731
rect 6546 17728 6552 17740
rect 5123 17700 6552 17728
rect 5123 17697 5135 17700
rect 5077 17691 5135 17697
rect 6546 17688 6552 17700
rect 6604 17728 6610 17740
rect 6604 17700 6684 17728
rect 6604 17688 6610 17700
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 6656 17660 6684 17700
rect 7742 17688 7748 17740
rect 7800 17688 7806 17740
rect 7834 17688 7840 17740
rect 7892 17688 7898 17740
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 12492 17700 13553 17728
rect 12492 17688 12498 17700
rect 13541 17697 13553 17700
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 14458 17688 14464 17740
rect 14516 17728 14522 17740
rect 14734 17728 14740 17740
rect 14516 17700 14740 17728
rect 14516 17688 14522 17700
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 14844 17737 14872 17768
rect 14918 17756 14924 17808
rect 14976 17796 14982 17808
rect 18782 17796 18788 17808
rect 14976 17768 18788 17796
rect 14976 17756 14982 17768
rect 18782 17756 18788 17768
rect 18840 17756 18846 17808
rect 24118 17756 24124 17808
rect 24176 17756 24182 17808
rect 14829 17731 14887 17737
rect 14829 17697 14841 17731
rect 14875 17697 14887 17731
rect 14829 17691 14887 17697
rect 15304 17700 18920 17728
rect 7558 17660 7564 17672
rect 6656 17632 7564 17660
rect 7558 17620 7564 17632
rect 7616 17660 7622 17672
rect 8294 17660 8300 17672
rect 7616 17632 8300 17660
rect 7616 17620 7622 17632
rect 8294 17620 8300 17632
rect 8352 17660 8358 17672
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 8352 17632 9229 17660
rect 8352 17620 8358 17632
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 11790 17660 11796 17672
rect 9217 17623 9275 17629
rect 10060 17632 11796 17660
rect 5350 17552 5356 17604
rect 5408 17552 5414 17604
rect 10060 17601 10088 17632
rect 11790 17620 11796 17632
rect 11848 17660 11854 17672
rect 12069 17663 12127 17669
rect 12069 17660 12081 17663
rect 11848 17632 12081 17660
rect 11848 17620 11854 17632
rect 12069 17629 12081 17632
rect 12115 17660 12127 17663
rect 15304 17660 15332 17700
rect 12115 17632 15332 17660
rect 12115 17629 12127 17632
rect 12069 17623 12127 17629
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 16758 17660 16764 17672
rect 15672 17632 16764 17660
rect 8757 17595 8815 17601
rect 8757 17561 8769 17595
rect 8803 17592 8815 17595
rect 10045 17595 10103 17601
rect 10045 17592 10057 17595
rect 8803 17564 10057 17592
rect 8803 17561 8815 17564
rect 8757 17555 8815 17561
rect 10045 17561 10057 17564
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 11057 17595 11115 17601
rect 11057 17561 11069 17595
rect 11103 17592 11115 17595
rect 11146 17592 11152 17604
rect 11103 17564 11152 17592
rect 11103 17561 11115 17564
rect 11057 17555 11115 17561
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 12713 17595 12771 17601
rect 12713 17561 12725 17595
rect 12759 17592 12771 17595
rect 13449 17595 13507 17601
rect 13449 17592 13461 17595
rect 12759 17564 13461 17592
rect 12759 17561 12771 17564
rect 12713 17555 12771 17561
rect 13449 17561 13461 17564
rect 13495 17592 13507 17595
rect 13630 17592 13636 17604
rect 13495 17564 13636 17592
rect 13495 17561 13507 17564
rect 13449 17555 13507 17561
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 15672 17592 15700 17632
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 16850 17620 16856 17672
rect 16908 17660 16914 17672
rect 17126 17660 17132 17672
rect 16908 17632 17132 17660
rect 16908 17620 16914 17632
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 17310 17620 17316 17672
rect 17368 17620 17374 17672
rect 18141 17663 18199 17669
rect 18141 17629 18153 17663
rect 18187 17660 18199 17663
rect 18322 17660 18328 17672
rect 18187 17632 18328 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18892 17669 18920 17700
rect 21082 17688 21088 17740
rect 21140 17728 21146 17740
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 21140 17700 21373 17728
rect 21140 17688 21146 17700
rect 21361 17697 21373 17700
rect 21407 17728 21419 17731
rect 21821 17731 21879 17737
rect 21821 17728 21833 17731
rect 21407 17700 21833 17728
rect 21407 17697 21419 17700
rect 21361 17691 21419 17697
rect 21821 17697 21833 17700
rect 21867 17697 21879 17731
rect 21821 17691 21879 17697
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17660 18935 17663
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18923 17632 19257 17660
rect 18923 17629 18935 17632
rect 18877 17623 18935 17629
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 23750 17620 23756 17672
rect 23808 17660 23814 17672
rect 24581 17663 24639 17669
rect 24581 17660 24593 17663
rect 23808 17632 24593 17660
rect 23808 17620 23814 17632
rect 24581 17629 24593 17632
rect 24627 17629 24639 17663
rect 24581 17623 24639 17629
rect 14568 17564 15700 17592
rect 16301 17595 16359 17601
rect 7650 17484 7656 17536
rect 7708 17484 7714 17536
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 8478 17524 8484 17536
rect 8435 17496 8484 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 8573 17527 8631 17533
rect 8573 17493 8585 17527
rect 8619 17524 8631 17527
rect 8938 17524 8944 17536
rect 8619 17496 8944 17524
rect 8619 17493 8631 17496
rect 8573 17487 8631 17493
rect 8938 17484 8944 17496
rect 8996 17524 9002 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 8996 17496 10333 17524
rect 8996 17484 9002 17496
rect 10321 17493 10333 17496
rect 10367 17524 10379 17527
rect 10502 17524 10508 17536
rect 10367 17496 10508 17524
rect 10367 17493 10379 17496
rect 10321 17487 10379 17493
rect 10502 17484 10508 17496
rect 10560 17524 10566 17536
rect 12618 17524 12624 17536
rect 10560 17496 12624 17524
rect 10560 17484 10566 17496
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17524 13415 17527
rect 14568 17524 14596 17564
rect 16301 17561 16313 17595
rect 16347 17592 16359 17595
rect 17328 17592 17356 17620
rect 16347 17564 17356 17592
rect 16347 17561 16359 17564
rect 16301 17555 16359 17561
rect 20622 17552 20628 17604
rect 20680 17552 20686 17604
rect 21085 17595 21143 17601
rect 21085 17561 21097 17595
rect 21131 17592 21143 17595
rect 21174 17592 21180 17604
rect 21131 17564 21180 17592
rect 21131 17561 21143 17564
rect 21085 17555 21143 17561
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 22094 17552 22100 17604
rect 22152 17552 22158 17604
rect 22480 17564 22586 17592
rect 22480 17536 22508 17564
rect 13403 17496 14596 17524
rect 14645 17527 14703 17533
rect 13403 17493 13415 17496
rect 13357 17487 13415 17493
rect 14645 17493 14657 17527
rect 14691 17524 14703 17527
rect 14918 17524 14924 17536
rect 14691 17496 14924 17524
rect 14691 17493 14703 17496
rect 14645 17487 14703 17493
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 15194 17484 15200 17536
rect 15252 17524 15258 17536
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15252 17496 15669 17524
rect 15252 17484 15258 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 16209 17527 16267 17533
rect 16209 17493 16221 17527
rect 16255 17524 16267 17527
rect 16666 17524 16672 17536
rect 16255 17496 16672 17524
rect 16255 17493 16267 17496
rect 16209 17487 16267 17493
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17862 17484 17868 17536
rect 17920 17524 17926 17536
rect 19426 17524 19432 17536
rect 17920 17496 19432 17524
rect 17920 17484 17926 17496
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 19613 17527 19671 17533
rect 19613 17493 19625 17527
rect 19659 17524 19671 17527
rect 19702 17524 19708 17536
rect 19659 17496 19708 17524
rect 19659 17493 19671 17496
rect 19613 17487 19671 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 22462 17484 22468 17536
rect 22520 17484 22526 17536
rect 25222 17484 25228 17536
rect 25280 17484 25286 17536
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 5350 17280 5356 17332
rect 5408 17280 5414 17332
rect 7466 17280 7472 17332
rect 7524 17280 7530 17332
rect 7650 17280 7656 17332
rect 7708 17320 7714 17332
rect 9125 17323 9183 17329
rect 9125 17320 9137 17323
rect 7708 17292 9137 17320
rect 7708 17280 7714 17292
rect 9125 17289 9137 17292
rect 9171 17289 9183 17323
rect 9125 17283 9183 17289
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 9582 17320 9588 17332
rect 9539 17292 9588 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10962 17320 10968 17332
rect 9916 17292 10968 17320
rect 9916 17280 9922 17292
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 11422 17280 11428 17332
rect 11480 17320 11486 17332
rect 12253 17323 12311 17329
rect 12253 17320 12265 17323
rect 11480 17292 12265 17320
rect 11480 17280 11486 17292
rect 12253 17289 12265 17292
rect 12299 17289 12311 17323
rect 12253 17283 12311 17289
rect 2409 17255 2467 17261
rect 2409 17221 2421 17255
rect 2455 17252 2467 17255
rect 4062 17252 4068 17264
rect 2455 17224 4068 17252
rect 2455 17221 2467 17224
rect 2409 17215 2467 17221
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 8297 17255 8355 17261
rect 8297 17221 8309 17255
rect 8343 17252 8355 17255
rect 11606 17252 11612 17264
rect 8343 17224 11612 17252
rect 8343 17221 8355 17224
rect 8297 17215 8355 17221
rect 11606 17212 11612 17224
rect 11664 17212 11670 17264
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6696 17156 6837 17184
rect 6696 17144 6702 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17184 9643 17187
rect 10042 17184 10048 17196
rect 9631 17156 10048 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17184 10839 17187
rect 10827 17156 11652 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 8386 17076 8392 17128
rect 8444 17076 8450 17128
rect 8570 17076 8576 17128
rect 8628 17076 8634 17128
rect 9398 17076 9404 17128
rect 9456 17116 9462 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9456 17088 9689 17116
rect 9456 17076 9462 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 9677 17079 9735 17085
rect 10502 17076 10508 17128
rect 10560 17116 10566 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10560 17088 10885 17116
rect 10560 17076 10566 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 8478 17048 8484 17060
rect 6656 17020 8484 17048
rect 6656 16992 6684 17020
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 9306 17008 9312 17060
rect 9364 17048 9370 17060
rect 10413 17051 10471 17057
rect 10413 17048 10425 17051
rect 9364 17020 10425 17048
rect 9364 17008 9370 17020
rect 10413 17017 10425 17020
rect 10459 17017 10471 17051
rect 10413 17011 10471 17017
rect 2317 16983 2375 16989
rect 2317 16949 2329 16983
rect 2363 16980 2375 16983
rect 2774 16980 2780 16992
rect 2363 16952 2780 16980
rect 2363 16949 2375 16952
rect 2317 16943 2375 16949
rect 2774 16940 2780 16952
rect 2832 16940 2838 16992
rect 6454 16940 6460 16992
rect 6512 16980 6518 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6512 16952 6561 16980
rect 6512 16940 6518 16952
rect 6549 16949 6561 16952
rect 6595 16980 6607 16983
rect 6638 16980 6644 16992
rect 6595 16952 6644 16980
rect 6595 16949 6607 16952
rect 6549 16943 6607 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 7742 16940 7748 16992
rect 7800 16980 7806 16992
rect 7929 16983 7987 16989
rect 7929 16980 7941 16983
rect 7800 16952 7941 16980
rect 7800 16940 7806 16952
rect 7929 16949 7941 16952
rect 7975 16949 7987 16983
rect 10888 16980 10916 17079
rect 10962 17076 10968 17128
rect 11020 17076 11026 17128
rect 11624 17057 11652 17156
rect 12268 17116 12296 17283
rect 12802 17280 12808 17332
rect 12860 17280 12866 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 13814 17320 13820 17332
rect 13219 17292 13820 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 13998 17280 14004 17332
rect 14056 17280 14062 17332
rect 16850 17280 16856 17332
rect 16908 17280 16914 17332
rect 18414 17320 18420 17332
rect 17052 17292 18420 17320
rect 13265 17255 13323 17261
rect 13265 17252 13277 17255
rect 12452 17224 13277 17252
rect 12452 17116 12480 17224
rect 13265 17221 13277 17224
rect 13311 17252 13323 17255
rect 13538 17252 13544 17264
rect 13311 17224 13544 17252
rect 13311 17221 13323 17224
rect 13265 17215 13323 17221
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 14369 17255 14427 17261
rect 14369 17221 14381 17255
rect 14415 17252 14427 17255
rect 15105 17255 15163 17261
rect 15105 17252 15117 17255
rect 14415 17224 15117 17252
rect 14415 17221 14427 17224
rect 14369 17215 14427 17221
rect 15105 17221 15117 17224
rect 15151 17252 15163 17255
rect 17052 17252 17080 17292
rect 18414 17280 18420 17292
rect 18472 17320 18478 17332
rect 18966 17320 18972 17332
rect 18472 17292 18972 17320
rect 18472 17280 18478 17292
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 21450 17280 21456 17332
rect 21508 17280 21514 17332
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 22649 17323 22707 17329
rect 22649 17320 22661 17323
rect 22152 17292 22661 17320
rect 22152 17280 22158 17292
rect 22649 17289 22661 17292
rect 22695 17289 22707 17323
rect 22649 17283 22707 17289
rect 15151 17224 17080 17252
rect 15151 17221 15163 17224
rect 15105 17215 15163 17221
rect 17862 17212 17868 17264
rect 17920 17212 17926 17264
rect 18325 17255 18383 17261
rect 18325 17221 18337 17255
rect 18371 17252 18383 17255
rect 18690 17252 18696 17264
rect 18371 17224 18696 17252
rect 18371 17221 18383 17224
rect 18325 17215 18383 17221
rect 18690 17212 18696 17224
rect 18748 17212 18754 17264
rect 19702 17212 19708 17264
rect 19760 17252 19766 17264
rect 19760 17224 22048 17252
rect 19760 17212 19766 17224
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17153 12587 17187
rect 15197 17187 15255 17193
rect 15197 17184 15209 17187
rect 12529 17147 12587 17153
rect 14476 17156 15209 17184
rect 12268 17088 12480 17116
rect 12544 17116 12572 17147
rect 12618 17116 12624 17128
rect 12544 17088 12624 17116
rect 12618 17076 12624 17088
rect 12676 17116 12682 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 12676 17088 13461 17116
rect 12676 17076 12682 17088
rect 13449 17085 13461 17088
rect 13495 17116 13507 17119
rect 13722 17116 13728 17128
rect 13495 17088 13728 17116
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 14476 17125 14504 17156
rect 15197 17153 15209 17156
rect 15243 17184 15255 17187
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15243 17156 15945 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 19242 17144 19248 17196
rect 19300 17184 19306 17196
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19300 17156 20177 17184
rect 19300 17144 19306 17156
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 22020 17193 22048 17224
rect 25130 17212 25136 17264
rect 25188 17212 25194 17264
rect 20809 17187 20867 17193
rect 20809 17184 20821 17187
rect 20772 17156 20821 17184
rect 20772 17144 20778 17156
rect 20809 17153 20821 17156
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 23201 17187 23259 17193
rect 23201 17153 23213 17187
rect 23247 17153 23259 17187
rect 23201 17147 23259 17153
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 13872 17088 14473 17116
rect 13872 17076 13878 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14550 17076 14556 17128
rect 14608 17076 14614 17128
rect 15654 17076 15660 17128
rect 15712 17076 15718 17128
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17116 15899 17119
rect 16390 17116 16396 17128
rect 15887 17088 16396 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 18601 17119 18659 17125
rect 18601 17085 18613 17119
rect 18647 17116 18659 17119
rect 21082 17116 21088 17128
rect 18647 17088 21088 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 21082 17076 21088 17088
rect 21140 17076 21146 17128
rect 21266 17076 21272 17128
rect 21324 17116 21330 17128
rect 23216 17116 23244 17147
rect 23658 17144 23664 17196
rect 23716 17184 23722 17196
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 23716 17156 23949 17184
rect 23716 17144 23722 17156
rect 23937 17153 23949 17156
rect 23983 17153 23995 17187
rect 23937 17147 23995 17153
rect 21324 17088 23244 17116
rect 21324 17076 21330 17088
rect 11609 17051 11667 17057
rect 11609 17017 11621 17051
rect 11655 17048 11667 17051
rect 11974 17048 11980 17060
rect 11655 17020 11980 17048
rect 11655 17017 11667 17020
rect 11609 17011 11667 17017
rect 11974 17008 11980 17020
rect 12032 17008 12038 17060
rect 18782 17008 18788 17060
rect 18840 17048 18846 17060
rect 20254 17048 20260 17060
rect 18840 17020 20260 17048
rect 18840 17008 18846 17020
rect 20254 17008 20260 17020
rect 20312 17008 20318 17060
rect 20349 17051 20407 17057
rect 20349 17017 20361 17051
rect 20395 17048 20407 17051
rect 20395 17020 22094 17048
rect 20395 17017 20407 17020
rect 20349 17011 20407 17017
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 10888 16952 11713 16980
rect 7929 16943 7987 16949
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 16301 16983 16359 16989
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 18598 16980 18604 16992
rect 16347 16952 18604 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 22066 16980 22094 17020
rect 23382 17008 23388 17060
rect 23440 17008 23446 17060
rect 22830 16980 22836 16992
rect 22066 16952 22836 16980
rect 22830 16940 22836 16952
rect 22888 16940 22894 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 5994 16736 6000 16788
rect 6052 16776 6058 16788
rect 6181 16779 6239 16785
rect 6181 16776 6193 16779
rect 6052 16748 6193 16776
rect 6052 16736 6058 16748
rect 6181 16745 6193 16748
rect 6227 16776 6239 16779
rect 7834 16776 7840 16788
rect 6227 16748 7840 16776
rect 6227 16745 6239 16748
rect 6181 16739 6239 16745
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 8297 16779 8355 16785
rect 8297 16745 8309 16779
rect 8343 16776 8355 16779
rect 8478 16776 8484 16788
rect 8343 16748 8484 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 16390 16736 16396 16788
rect 16448 16736 16454 16788
rect 18690 16736 18696 16788
rect 18748 16736 18754 16788
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 22462 16776 22468 16788
rect 20680 16748 22468 16776
rect 20680 16736 20686 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 25222 16776 25228 16788
rect 23400 16748 25228 16776
rect 8662 16708 8668 16720
rect 7852 16680 8668 16708
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 7852 16640 7880 16680
rect 8662 16668 8668 16680
rect 8720 16708 8726 16720
rect 9490 16708 9496 16720
rect 8720 16680 9496 16708
rect 8720 16668 8726 16680
rect 9490 16668 9496 16680
rect 9548 16668 9554 16720
rect 10796 16680 11008 16708
rect 6972 16612 7880 16640
rect 7929 16643 7987 16649
rect 6972 16600 6978 16612
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 8294 16640 8300 16652
rect 7975 16612 8300 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 9214 16600 9220 16652
rect 9272 16600 9278 16652
rect 10796 16649 10824 16680
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16640 9367 16643
rect 10781 16643 10839 16649
rect 9355 16612 10732 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 1762 16532 1768 16584
rect 1820 16532 1826 16584
rect 9232 16572 9260 16600
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 9232 16544 9413 16572
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9401 16535 9459 16541
rect 9490 16532 9496 16584
rect 9548 16532 9554 16584
rect 10704 16572 10732 16612
rect 10781 16609 10793 16643
rect 10827 16609 10839 16643
rect 10781 16603 10839 16609
rect 10870 16600 10876 16652
rect 10928 16600 10934 16652
rect 10980 16640 11008 16680
rect 12618 16640 12624 16652
rect 10980 16612 12624 16640
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 13354 16640 13360 16652
rect 13035 16612 13360 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 13814 16600 13820 16652
rect 13872 16600 13878 16652
rect 17586 16600 17592 16652
rect 17644 16640 17650 16652
rect 17862 16640 17868 16652
rect 17644 16612 17868 16640
rect 17644 16600 17650 16612
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 21269 16643 21327 16649
rect 21269 16609 21281 16643
rect 21315 16640 21327 16643
rect 22186 16640 22192 16652
rect 21315 16612 22192 16640
rect 21315 16609 21327 16612
rect 21269 16603 21327 16609
rect 22186 16600 22192 16612
rect 22244 16600 22250 16652
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16640 23259 16643
rect 23400 16640 23428 16748
rect 25222 16736 25228 16748
rect 25280 16736 25286 16788
rect 24026 16708 24032 16720
rect 23492 16680 24032 16708
rect 23492 16649 23520 16680
rect 24026 16668 24032 16680
rect 24084 16668 24090 16720
rect 23247 16612 23428 16640
rect 23477 16643 23535 16649
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 23477 16609 23489 16643
rect 23523 16609 23535 16643
rect 23477 16603 23535 16609
rect 11514 16572 11520 16584
rect 10704 16544 11520 16572
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16572 13323 16575
rect 13446 16572 13452 16584
rect 13311 16544 13452 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16572 18107 16575
rect 18506 16572 18512 16584
rect 18095 16544 18512 16572
rect 18095 16541 18107 16544
rect 18049 16535 18107 16541
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 20806 16532 20812 16584
rect 20864 16532 20870 16584
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 21048 16544 21097 16572
rect 21048 16532 21054 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 2501 16467 2559 16473
rect 6914 16464 6920 16516
rect 6972 16464 6978 16516
rect 7650 16464 7656 16516
rect 7708 16464 7714 16516
rect 10689 16507 10747 16513
rect 8128 16476 10364 16504
rect 7558 16396 7564 16448
rect 7616 16436 7622 16448
rect 8128 16436 8156 16476
rect 7616 16408 8156 16436
rect 7616 16396 7622 16408
rect 9858 16396 9864 16448
rect 9916 16396 9922 16448
rect 10336 16445 10364 16476
rect 10689 16473 10701 16507
rect 10735 16504 10747 16507
rect 16482 16504 16488 16516
rect 10735 16476 11652 16504
rect 12558 16476 16488 16504
rect 10735 16473 10747 16476
rect 10689 16467 10747 16473
rect 10321 16439 10379 16445
rect 10321 16405 10333 16439
rect 10367 16405 10379 16439
rect 10321 16399 10379 16405
rect 11514 16396 11520 16448
rect 11572 16396 11578 16448
rect 11624 16436 11652 16476
rect 16482 16464 16488 16476
rect 16540 16464 16546 16516
rect 20824 16504 20852 16532
rect 21174 16504 21180 16516
rect 20824 16476 21180 16504
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 22462 16464 22468 16516
rect 22520 16464 22526 16516
rect 12802 16436 12808 16448
rect 11624 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 19334 16396 19340 16448
rect 19392 16396 19398 16448
rect 19978 16396 19984 16448
rect 20036 16436 20042 16448
rect 20073 16439 20131 16445
rect 20073 16436 20085 16439
rect 20036 16408 20085 16436
rect 20036 16396 20042 16408
rect 20073 16405 20085 16408
rect 20119 16405 20131 16439
rect 20073 16399 20131 16405
rect 20806 16396 20812 16448
rect 20864 16436 20870 16448
rect 21729 16439 21787 16445
rect 21729 16436 21741 16439
rect 20864 16408 21741 16436
rect 20864 16396 20870 16408
rect 21729 16405 21741 16408
rect 21775 16405 21787 16439
rect 21729 16399 21787 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 7377 16235 7435 16241
rect 7377 16232 7389 16235
rect 6788 16204 7389 16232
rect 6788 16192 6794 16204
rect 7377 16201 7389 16204
rect 7423 16201 7435 16235
rect 7377 16195 7435 16201
rect 7742 16192 7748 16244
rect 7800 16192 7806 16244
rect 7837 16235 7895 16241
rect 7837 16201 7849 16235
rect 7883 16232 7895 16235
rect 10321 16235 10379 16241
rect 10321 16232 10333 16235
rect 7883 16204 10333 16232
rect 7883 16201 7895 16204
rect 7837 16195 7895 16201
rect 10321 16201 10333 16204
rect 10367 16201 10379 16235
rect 10321 16195 10379 16201
rect 10686 16192 10692 16244
rect 10744 16192 10750 16244
rect 19886 16192 19892 16244
rect 19944 16192 19950 16244
rect 19978 16192 19984 16244
rect 20036 16192 20042 16244
rect 20162 16192 20168 16244
rect 20220 16232 20226 16244
rect 22281 16235 22339 16241
rect 22281 16232 22293 16235
rect 20220 16204 22293 16232
rect 20220 16192 20226 16204
rect 22281 16201 22293 16204
rect 22327 16201 22339 16235
rect 22281 16195 22339 16201
rect 9309 16167 9367 16173
rect 9309 16133 9321 16167
rect 9355 16164 9367 16167
rect 11790 16164 11796 16176
rect 9355 16136 11796 16164
rect 9355 16133 9367 16136
rect 9309 16127 9367 16133
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 15102 16124 15108 16176
rect 15160 16164 15166 16176
rect 15657 16167 15715 16173
rect 15657 16164 15669 16167
rect 15160 16136 15669 16164
rect 15160 16124 15166 16136
rect 15657 16133 15669 16136
rect 15703 16164 15715 16167
rect 17494 16164 17500 16176
rect 15703 16136 17500 16164
rect 15703 16133 15715 16136
rect 15657 16127 15715 16133
rect 17494 16124 17500 16136
rect 17552 16164 17558 16176
rect 20990 16164 20996 16176
rect 17552 16136 20996 16164
rect 17552 16124 17558 16136
rect 20990 16124 20996 16136
rect 21048 16124 21054 16176
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 9217 16099 9275 16105
rect 7892 16068 8616 16096
rect 7892 16056 7898 16068
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 16028 8079 16031
rect 8478 16028 8484 16040
rect 8067 16000 8484 16028
rect 8067 15997 8079 16000
rect 8021 15991 8079 15997
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 8588 16028 8616 16068
rect 9217 16065 9229 16099
rect 9263 16096 9275 16099
rect 9263 16068 9996 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 9401 16031 9459 16037
rect 9401 16028 9413 16031
rect 8588 16000 9413 16028
rect 9401 15997 9413 16000
rect 9447 15997 9459 16031
rect 9968 16028 9996 16068
rect 10042 16056 10048 16108
rect 10100 16056 10106 16108
rect 11698 16096 11704 16108
rect 10704 16068 11704 16096
rect 10704 16028 10732 16068
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12342 16056 12348 16108
rect 12400 16056 12406 16108
rect 20806 16056 20812 16108
rect 20864 16056 20870 16108
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16096 22431 16099
rect 23201 16099 23259 16105
rect 23201 16096 23213 16099
rect 22419 16068 23213 16096
rect 22419 16065 22431 16068
rect 22373 16059 22431 16065
rect 23201 16065 23213 16068
rect 23247 16065 23259 16099
rect 23201 16059 23259 16065
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16096 24179 16099
rect 24302 16096 24308 16108
rect 24167 16068 24308 16096
rect 24167 16065 24179 16068
rect 24121 16059 24179 16065
rect 24302 16056 24308 16068
rect 24360 16056 24366 16108
rect 9968 16000 10732 16028
rect 10781 16031 10839 16037
rect 9401 15991 9459 15997
rect 10781 15997 10793 16031
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 8846 15920 8852 15972
rect 8904 15920 8910 15972
rect 10796 15960 10824 15991
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 12360 16028 12388 16056
rect 11664 16000 12388 16028
rect 18141 16031 18199 16037
rect 11664 15988 11670 16000
rect 18141 15997 18153 16031
rect 18187 16028 18199 16031
rect 18414 16028 18420 16040
rect 18187 16000 18420 16028
rect 18187 15997 18199 16000
rect 18141 15991 18199 15997
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 19150 15988 19156 16040
rect 19208 15988 19214 16040
rect 19794 15988 19800 16040
rect 19852 15988 19858 16040
rect 21450 16028 21456 16040
rect 20364 16000 21456 16028
rect 12802 15960 12808 15972
rect 10796 15932 12808 15960
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 14090 15920 14096 15972
rect 14148 15960 14154 15972
rect 20364 15969 20392 16000
rect 21450 15988 21456 16000
rect 21508 15988 21514 16040
rect 22189 16031 22247 16037
rect 22189 15997 22201 16031
rect 22235 15997 22247 16031
rect 22189 15991 22247 15997
rect 20349 15963 20407 15969
rect 14148 15932 18736 15960
rect 14148 15920 14154 15932
rect 18708 15904 18736 15932
rect 20349 15929 20361 15963
rect 20395 15929 20407 15963
rect 22204 15960 22232 15991
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 23566 15960 23572 15972
rect 22204 15932 23572 15960
rect 20349 15923 20407 15929
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 11701 15895 11759 15901
rect 11701 15892 11713 15895
rect 10100 15864 11713 15892
rect 10100 15852 10106 15864
rect 11701 15861 11713 15864
rect 11747 15861 11759 15895
rect 11701 15855 11759 15861
rect 16482 15852 16488 15904
rect 16540 15892 16546 15904
rect 17586 15892 17592 15904
rect 16540 15864 17592 15892
rect 16540 15852 16546 15864
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 18690 15852 18696 15904
rect 18748 15852 18754 15904
rect 21358 15852 21364 15904
rect 21416 15892 21422 15904
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 21416 15864 21465 15892
rect 21416 15852 21422 15864
rect 21453 15861 21465 15864
rect 21499 15861 21511 15895
rect 21453 15855 21511 15861
rect 22646 15852 22652 15904
rect 22704 15892 22710 15904
rect 22741 15895 22799 15901
rect 22741 15892 22753 15895
rect 22704 15864 22753 15892
rect 22704 15852 22710 15864
rect 22741 15861 22753 15864
rect 22787 15861 22799 15895
rect 22741 15855 22799 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7708 15660 7941 15688
rect 7708 15648 7714 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 7929 15651 7987 15657
rect 8386 15648 8392 15700
rect 8444 15688 8450 15700
rect 9585 15691 9643 15697
rect 9585 15688 9597 15691
rect 8444 15660 9597 15688
rect 8444 15648 8450 15660
rect 9585 15657 9597 15660
rect 9631 15657 9643 15691
rect 9585 15651 9643 15657
rect 13191 15691 13249 15697
rect 13191 15657 13203 15691
rect 13237 15688 13249 15691
rect 14550 15688 14556 15700
rect 13237 15660 14556 15688
rect 13237 15657 13249 15660
rect 13191 15651 13249 15657
rect 14550 15648 14556 15660
rect 14608 15688 14614 15700
rect 17218 15688 17224 15700
rect 14608 15660 17224 15688
rect 14608 15648 14614 15660
rect 8570 15620 8576 15632
rect 7484 15592 8576 15620
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7484 15493 7512 15592
rect 8570 15580 8576 15592
rect 8628 15620 8634 15632
rect 10870 15620 10876 15632
rect 8628 15592 10876 15620
rect 8628 15580 8634 15592
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 11698 15552 11704 15564
rect 10275 15524 11704 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 13446 15552 13452 15564
rect 12492 15524 13452 15552
rect 12492 15512 12498 15524
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 15381 15555 15439 15561
rect 15381 15521 15393 15555
rect 15427 15552 15439 15555
rect 15488 15552 15516 15660
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 17681 15691 17739 15697
rect 17681 15657 17693 15691
rect 17727 15688 17739 15691
rect 18506 15688 18512 15700
rect 17727 15660 18512 15688
rect 17727 15657 17739 15660
rect 17681 15651 17739 15657
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 20165 15691 20223 15697
rect 20165 15657 20177 15691
rect 20211 15688 20223 15691
rect 20898 15688 20904 15700
rect 20211 15660 20904 15688
rect 20211 15657 20223 15660
rect 20165 15651 20223 15657
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 22278 15648 22284 15700
rect 22336 15648 22342 15700
rect 22296 15620 22324 15648
rect 19628 15592 22324 15620
rect 15427 15524 15516 15552
rect 15933 15555 15991 15561
rect 15427 15521 15439 15524
rect 15381 15515 15439 15521
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 18233 15555 18291 15561
rect 15979 15524 17724 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 7340 15456 7481 15484
rect 7340 15444 7346 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15484 8631 15487
rect 9398 15484 9404 15496
rect 8619 15456 9404 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10594 15484 10600 15496
rect 10091 15456 10600 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 15197 15487 15255 15493
rect 15197 15484 15209 15487
rect 14608 15456 15209 15484
rect 14608 15444 14614 15456
rect 15197 15453 15209 15456
rect 15243 15453 15255 15487
rect 17586 15484 17592 15496
rect 17342 15456 17592 15484
rect 15197 15447 15255 15453
rect 14277 15419 14335 15425
rect 11256 15388 12006 15416
rect 11256 15360 11284 15388
rect 6825 15351 6883 15357
rect 6825 15317 6837 15351
rect 6871 15348 6883 15351
rect 7006 15348 7012 15360
rect 6871 15320 7012 15348
rect 6871 15317 6883 15320
rect 6825 15311 6883 15317
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 9217 15351 9275 15357
rect 9217 15348 9229 15351
rect 7616 15320 9229 15348
rect 7616 15308 7622 15320
rect 9217 15317 9229 15320
rect 9263 15348 9275 15351
rect 9953 15351 10011 15357
rect 9953 15348 9965 15351
rect 9263 15320 9965 15348
rect 9263 15317 9275 15320
rect 9217 15311 9275 15317
rect 9953 15317 9965 15320
rect 9999 15348 10011 15351
rect 11054 15348 11060 15360
rect 9999 15320 11060 15348
rect 9999 15317 10011 15320
rect 9953 15311 10011 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11238 15308 11244 15360
rect 11296 15308 11302 15360
rect 11698 15308 11704 15360
rect 11756 15308 11762 15360
rect 11900 15348 11928 15388
rect 14277 15385 14289 15419
rect 14323 15416 14335 15419
rect 15010 15416 15016 15428
rect 14323 15388 15016 15416
rect 14323 15385 14335 15388
rect 14277 15379 14335 15385
rect 15010 15376 15016 15388
rect 15068 15376 15074 15428
rect 15102 15376 15108 15428
rect 15160 15376 15166 15428
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 11900 15320 13737 15348
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 14461 15351 14519 15357
rect 14461 15317 14473 15351
rect 14507 15348 14519 15351
rect 14550 15348 14556 15360
rect 14507 15320 14556 15348
rect 14507 15317 14519 15320
rect 14461 15311 14519 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 15212 15348 15240 15447
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 17696 15484 17724 15524
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 18782 15552 18788 15564
rect 18279 15524 18788 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 19628 15561 19656 15592
rect 19613 15555 19671 15561
rect 19613 15521 19625 15555
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 20806 15512 20812 15564
rect 20864 15512 20870 15564
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15552 20959 15555
rect 21174 15552 21180 15564
rect 20947 15524 21180 15552
rect 20947 15521 20959 15524
rect 20901 15515 20959 15521
rect 21174 15512 21180 15524
rect 21232 15552 21238 15564
rect 22281 15555 22339 15561
rect 22281 15552 22293 15555
rect 21232 15524 22293 15552
rect 21232 15512 21238 15524
rect 22281 15521 22293 15524
rect 22327 15521 22339 15555
rect 22281 15515 22339 15521
rect 18322 15484 18328 15496
rect 17696 15456 18328 15484
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 18690 15484 18696 15496
rect 18555 15456 18696 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 19208 15456 19809 15484
rect 19208 15444 19214 15456
rect 19797 15453 19809 15456
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 21600 15456 22017 15484
rect 21600 15444 21606 15456
rect 22005 15453 22017 15456
rect 22051 15453 22063 15487
rect 22005 15447 22063 15453
rect 22738 15444 22744 15496
rect 22796 15444 22802 15496
rect 16206 15376 16212 15428
rect 16264 15376 16270 15428
rect 19334 15416 19340 15428
rect 17512 15388 19340 15416
rect 17512 15348 17540 15388
rect 19334 15376 19340 15388
rect 19392 15416 19398 15428
rect 19705 15419 19763 15425
rect 19705 15416 19717 15419
rect 19392 15388 19717 15416
rect 19392 15376 19398 15388
rect 19705 15385 19717 15388
rect 19751 15385 19763 15419
rect 19705 15379 19763 15385
rect 23845 15419 23903 15425
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 25498 15416 25504 15428
rect 23891 15388 25504 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 25498 15376 25504 15388
rect 25556 15376 25562 15428
rect 15212 15320 17540 15348
rect 18417 15351 18475 15357
rect 18417 15317 18429 15351
rect 18463 15348 18475 15351
rect 18690 15348 18696 15360
rect 18463 15320 18696 15348
rect 18463 15317 18475 15320
rect 18417 15311 18475 15317
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 18877 15351 18935 15357
rect 18877 15317 18889 15351
rect 18923 15348 18935 15351
rect 19518 15348 19524 15360
rect 18923 15320 19524 15348
rect 18923 15317 18935 15320
rect 18877 15311 18935 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 20990 15308 20996 15360
rect 21048 15308 21054 15360
rect 21361 15351 21419 15357
rect 21361 15317 21373 15351
rect 21407 15348 21419 15351
rect 21726 15348 21732 15360
rect 21407 15320 21732 15348
rect 21407 15317 21419 15320
rect 21361 15311 21419 15317
rect 21726 15308 21732 15320
rect 21784 15308 21790 15360
rect 21821 15351 21879 15357
rect 21821 15317 21833 15351
rect 21867 15348 21879 15351
rect 21910 15348 21916 15360
rect 21867 15320 21916 15348
rect 21867 15317 21879 15320
rect 21821 15311 21879 15317
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 8757 15147 8815 15153
rect 8757 15144 8769 15147
rect 6880 15116 8769 15144
rect 6880 15104 6886 15116
rect 7006 15036 7012 15088
rect 7064 15036 7070 15088
rect 7392 15076 7420 15116
rect 8757 15113 8769 15116
rect 8803 15113 8815 15147
rect 8757 15107 8815 15113
rect 8772 15076 8800 15107
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 13633 15147 13691 15153
rect 13633 15144 13645 15147
rect 11940 15116 13645 15144
rect 11940 15104 11946 15116
rect 13633 15113 13645 15116
rect 13679 15113 13691 15147
rect 13633 15107 13691 15113
rect 14090 15104 14096 15156
rect 14148 15104 14154 15156
rect 16206 15104 16212 15156
rect 16264 15144 16270 15156
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 16264 15116 16313 15144
rect 16264 15104 16270 15116
rect 16301 15113 16313 15116
rect 16347 15113 16359 15147
rect 17494 15144 17500 15156
rect 16301 15107 16359 15113
rect 17052 15116 17500 15144
rect 7392 15048 7498 15076
rect 8772 15048 9706 15076
rect 10778 15036 10784 15088
rect 10836 15076 10842 15088
rect 10873 15079 10931 15085
rect 10873 15076 10885 15079
rect 10836 15048 10885 15076
rect 10836 15036 10842 15048
rect 10873 15045 10885 15048
rect 10919 15045 10931 15079
rect 10873 15039 10931 15045
rect 12434 15036 12440 15088
rect 12492 15076 12498 15088
rect 12710 15076 12716 15088
rect 12492 15048 12716 15076
rect 12492 15036 12498 15048
rect 12710 15036 12716 15048
rect 12768 15036 12774 15088
rect 13357 15079 13415 15085
rect 13357 15045 13369 15079
rect 13403 15076 13415 15079
rect 13446 15076 13452 15088
rect 13403 15048 13452 15076
rect 13403 15045 13415 15048
rect 13357 15039 13415 15045
rect 13446 15036 13452 15048
rect 13504 15076 13510 15088
rect 14108 15076 14136 15104
rect 13504 15048 14136 15076
rect 13504 15036 13510 15048
rect 15010 15036 15016 15088
rect 15068 15036 15074 15088
rect 17052 15085 17080 15116
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 18141 15147 18199 15153
rect 18141 15113 18153 15147
rect 18187 15144 18199 15147
rect 18414 15144 18420 15156
rect 18187 15116 18420 15144
rect 18187 15113 18199 15116
rect 18141 15107 18199 15113
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 19058 15104 19064 15156
rect 19116 15144 19122 15156
rect 19116 15116 20668 15144
rect 19116 15104 19122 15116
rect 17037 15079 17095 15085
rect 17037 15045 17049 15079
rect 17083 15045 17095 15079
rect 18506 15076 18512 15088
rect 17037 15039 17095 15045
rect 17972 15048 18512 15076
rect 11514 14968 11520 15020
rect 11572 15008 11578 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11572 14980 11713 15008
rect 11572 14968 11578 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14056 14980 14320 15008
rect 14056 14968 14062 14980
rect 6733 14943 6791 14949
rect 6733 14909 6745 14943
rect 6779 14909 6791 14943
rect 6733 14903 6791 14909
rect 6748 14804 6776 14903
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 7650 14940 7656 14952
rect 7156 14912 7656 14940
rect 7156 14900 7162 14912
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 11146 14900 11152 14952
rect 11204 14940 11210 14952
rect 12342 14940 12348 14952
rect 11204 14912 12348 14940
rect 11204 14900 11210 14912
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 14182 14900 14188 14952
rect 14240 14900 14246 14952
rect 14292 14940 14320 14980
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 16666 14940 16672 14952
rect 14292 14912 16672 14940
rect 16666 14900 16672 14912
rect 16724 14940 16730 14952
rect 17218 14940 17224 14952
rect 16724 14912 17224 14940
rect 16724 14900 16730 14912
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 17972 14949 18000 15048
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 19794 15036 19800 15088
rect 19852 15036 19858 15088
rect 20640 15076 20668 15116
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 20809 15147 20867 15153
rect 20809 15144 20821 15147
rect 20772 15116 20821 15144
rect 20772 15104 20778 15116
rect 20809 15113 20821 15116
rect 20855 15113 20867 15147
rect 20809 15107 20867 15113
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 24394 15144 24400 15156
rect 21876 15116 24400 15144
rect 21876 15104 21882 15116
rect 24394 15104 24400 15116
rect 24452 15104 24458 15156
rect 20640 15048 22094 15076
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 19061 15011 19119 15017
rect 19061 15008 19073 15011
rect 18380 14980 19073 15008
rect 18380 14968 18386 14980
rect 19061 14977 19073 14980
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 15008 21511 15011
rect 21634 15008 21640 15020
rect 21499 14980 21640 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 21634 14968 21640 14980
rect 21692 14968 21698 15020
rect 22066 15008 22094 15048
rect 22370 15036 22376 15088
rect 22428 15076 22434 15088
rect 22428 15048 23980 15076
rect 22428 15036 22434 15048
rect 23952 15017 23980 15048
rect 22741 15011 22799 15017
rect 22741 15008 22753 15011
rect 22066 14980 22753 15008
rect 22741 14977 22753 14980
rect 22787 14977 22799 15011
rect 22741 14971 22799 14977
rect 23937 15011 23995 15017
rect 23937 14977 23949 15011
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 17957 14943 18015 14949
rect 17957 14909 17969 14943
rect 18003 14909 18015 14943
rect 17957 14903 18015 14909
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 18598 14940 18604 14952
rect 18095 14912 18604 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 19337 14943 19395 14949
rect 19337 14909 19349 14943
rect 19383 14940 19395 14943
rect 19426 14940 19432 14952
rect 19383 14912 19432 14940
rect 19383 14909 19395 14912
rect 19337 14903 19395 14909
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 19794 14900 19800 14952
rect 19852 14940 19858 14952
rect 21818 14940 21824 14952
rect 19852 14912 21824 14940
rect 19852 14900 19858 14912
rect 21818 14900 21824 14912
rect 21876 14900 21882 14952
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 14826 14832 14832 14884
rect 14884 14832 14890 14884
rect 16574 14832 16580 14884
rect 16632 14872 16638 14884
rect 16853 14875 16911 14881
rect 16853 14872 16865 14875
rect 16632 14844 16865 14872
rect 16632 14832 16638 14844
rect 16853 14841 16865 14844
rect 16899 14841 16911 14875
rect 18690 14872 18696 14884
rect 16853 14835 16911 14841
rect 18432 14844 18696 14872
rect 8294 14804 8300 14816
rect 6748 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 8478 14764 8484 14816
rect 8536 14764 8542 14816
rect 9398 14764 9404 14816
rect 9456 14764 9462 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 12345 14807 12403 14813
rect 12345 14804 12357 14807
rect 9732 14776 12357 14804
rect 9732 14764 9738 14776
rect 12345 14773 12357 14776
rect 12391 14773 12403 14807
rect 12345 14767 12403 14773
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 18432 14804 18460 14844
rect 18690 14832 18696 14844
rect 18748 14832 18754 14884
rect 21174 14872 21180 14884
rect 20548 14844 21180 14872
rect 15620 14776 18460 14804
rect 18509 14807 18567 14813
rect 15620 14764 15626 14776
rect 18509 14773 18521 14807
rect 18555 14804 18567 14807
rect 20548 14804 20576 14844
rect 21174 14832 21180 14844
rect 21232 14832 21238 14884
rect 22925 14875 22983 14881
rect 22925 14841 22937 14875
rect 22971 14872 22983 14875
rect 23842 14872 23848 14884
rect 22971 14844 23848 14872
rect 22971 14841 22983 14844
rect 22925 14835 22983 14841
rect 23842 14832 23848 14844
rect 23900 14832 23906 14884
rect 18555 14776 20576 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 21269 14807 21327 14813
rect 21269 14804 21281 14807
rect 20680 14776 21281 14804
rect 20680 14764 20686 14776
rect 21269 14773 21281 14776
rect 21315 14773 21327 14807
rect 21269 14767 21327 14773
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 6825 14603 6883 14609
rect 6825 14569 6837 14603
rect 6871 14600 6883 14603
rect 7282 14600 7288 14612
rect 6871 14572 7288 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7708 14572 11192 14600
rect 7708 14560 7714 14572
rect 11164 14532 11192 14572
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11977 14603 12035 14609
rect 11977 14600 11989 14603
rect 11296 14572 11989 14600
rect 11296 14560 11302 14572
rect 11977 14569 11989 14572
rect 12023 14569 12035 14603
rect 11977 14563 12035 14569
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12676 14572 13001 14600
rect 12676 14560 12682 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15654 14600 15660 14612
rect 15611 14572 15660 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16298 14560 16304 14612
rect 16356 14600 16362 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 16356 14572 20453 14600
rect 16356 14560 16362 14572
rect 20441 14569 20453 14572
rect 20487 14600 20499 14603
rect 20990 14600 20996 14612
rect 20487 14572 20996 14600
rect 20487 14569 20499 14572
rect 20441 14563 20499 14569
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 12713 14535 12771 14541
rect 11164 14504 11652 14532
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8352 14436 8585 14464
rect 8352 14424 8358 14436
rect 8573 14433 8585 14436
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 9861 14467 9919 14473
rect 9861 14433 9873 14467
rect 9907 14464 9919 14467
rect 11146 14464 11152 14476
rect 9907 14436 11152 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 6270 14288 6276 14340
rect 6328 14328 6334 14340
rect 6822 14328 6828 14340
rect 6328 14300 6828 14328
rect 6328 14288 6334 14300
rect 6822 14288 6828 14300
rect 6880 14328 6886 14340
rect 8297 14331 8355 14337
rect 6880 14300 7130 14328
rect 6880 14288 6886 14300
rect 8297 14297 8309 14331
rect 8343 14328 8355 14331
rect 10042 14328 10048 14340
rect 8343 14300 10048 14328
rect 8343 14297 8355 14300
rect 8297 14291 8355 14297
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 10134 14288 10140 14340
rect 10192 14288 10198 14340
rect 10244 14300 10626 14328
rect 8938 14220 8944 14272
rect 8996 14260 9002 14272
rect 10244 14260 10272 14300
rect 11624 14269 11652 14504
rect 12713 14501 12725 14535
rect 12759 14532 12771 14535
rect 13722 14532 13728 14544
rect 12759 14504 13728 14532
rect 12759 14501 12771 14504
rect 12713 14495 12771 14501
rect 12529 14467 12587 14473
rect 12529 14433 12541 14467
rect 12575 14464 12587 14467
rect 13446 14464 13452 14476
rect 12575 14436 13452 14464
rect 12575 14433 12587 14436
rect 12529 14427 12587 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 13556 14473 13584 14504
rect 13722 14492 13728 14504
rect 13780 14492 13786 14544
rect 18690 14492 18696 14544
rect 18748 14532 18754 14544
rect 18969 14535 19027 14541
rect 18969 14532 18981 14535
rect 18748 14504 18981 14532
rect 18748 14492 18754 14504
rect 18969 14501 18981 14504
rect 19015 14501 19027 14535
rect 18969 14495 19027 14501
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 14553 14467 14611 14473
rect 13587 14436 13621 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 16022 14464 16028 14476
rect 14599 14436 16028 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 17402 14464 17408 14476
rect 17359 14436 17408 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 17402 14424 17408 14436
rect 17460 14464 17466 14476
rect 18322 14464 18328 14476
rect 17460 14436 18328 14464
rect 17460 14424 17466 14436
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 21358 14424 21364 14476
rect 21416 14424 21422 14476
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 14737 14399 14795 14405
rect 14737 14396 14749 14399
rect 14700 14368 14749 14396
rect 14700 14356 14706 14368
rect 14737 14365 14749 14368
rect 14783 14365 14795 14399
rect 15562 14396 15568 14408
rect 14737 14359 14795 14365
rect 14936 14368 15568 14396
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13998 14328 14004 14340
rect 13403 14300 14004 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 8996 14232 10272 14260
rect 11609 14263 11667 14269
rect 8996 14220 9002 14232
rect 11609 14229 11621 14263
rect 11655 14260 11667 14263
rect 11882 14260 11888 14272
rect 11655 14232 11888 14260
rect 11655 14229 11667 14232
rect 11609 14223 11667 14229
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 14645 14263 14703 14269
rect 14645 14229 14657 14263
rect 14691 14260 14703 14263
rect 14936 14260 14964 14368
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 17770 14356 17776 14408
rect 17828 14356 17834 14408
rect 19610 14356 19616 14408
rect 19668 14356 19674 14408
rect 21082 14356 21088 14408
rect 21140 14356 21146 14408
rect 22830 14356 22836 14408
rect 22888 14396 22894 14408
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 22888 14368 23397 14396
rect 22888 14356 22894 14368
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 16482 14288 16488 14340
rect 16540 14288 16546 14340
rect 17037 14331 17095 14337
rect 17037 14297 17049 14331
rect 17083 14328 17095 14331
rect 18417 14331 18475 14337
rect 18417 14328 18429 14331
rect 17083 14300 18429 14328
rect 17083 14297 17095 14300
rect 17037 14291 17095 14297
rect 18417 14297 18429 14300
rect 18463 14297 18475 14331
rect 18417 14291 18475 14297
rect 22370 14288 22376 14340
rect 22428 14288 22434 14340
rect 23569 14331 23627 14337
rect 23569 14297 23581 14331
rect 23615 14328 23627 14331
rect 23934 14328 23940 14340
rect 23615 14300 23940 14328
rect 23615 14297 23627 14300
rect 23569 14291 23627 14297
rect 23934 14288 23940 14300
rect 23992 14288 23998 14340
rect 14691 14232 14964 14260
rect 15105 14263 15163 14269
rect 14691 14229 14703 14232
rect 14645 14223 14703 14229
rect 15105 14229 15117 14263
rect 15151 14260 15163 14263
rect 16390 14260 16396 14272
rect 15151 14232 16396 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 19429 14263 19487 14269
rect 19429 14229 19441 14263
rect 19475 14260 19487 14263
rect 19702 14260 19708 14272
rect 19475 14232 19708 14260
rect 19475 14229 19487 14232
rect 19429 14223 19487 14229
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 22830 14220 22836 14272
rect 22888 14220 22894 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 8938 14056 8944 14068
rect 6880 14028 8944 14056
rect 6880 14016 6886 14028
rect 8294 13988 8300 14000
rect 7944 13960 8300 13988
rect 2774 13880 2780 13932
rect 2832 13880 2838 13932
rect 7944 13929 7972 13960
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 8588 13988 8616 14028
rect 8938 14016 8944 14028
rect 8996 14056 9002 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 8996 14028 10241 14056
rect 8996 14016 9002 14028
rect 10229 14025 10241 14028
rect 10275 14056 10287 14059
rect 11238 14056 11244 14068
rect 10275 14028 11244 14056
rect 10275 14025 10287 14028
rect 10229 14019 10287 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11790 14016 11796 14068
rect 11848 14016 11854 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 12989 14059 13047 14065
rect 12989 14056 13001 14059
rect 12860 14028 13001 14056
rect 12860 14016 12866 14028
rect 12989 14025 13001 14028
rect 13035 14025 13047 14059
rect 12989 14019 13047 14025
rect 13357 14059 13415 14065
rect 13357 14025 13369 14059
rect 13403 14056 13415 14059
rect 14734 14056 14740 14068
rect 13403 14028 14740 14056
rect 13403 14025 13415 14028
rect 13357 14019 13415 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 19426 14016 19432 14068
rect 19484 14016 19490 14068
rect 19518 14016 19524 14068
rect 19576 14056 19582 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 19576 14028 20545 14056
rect 19576 14016 19582 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 20533 14019 20591 14025
rect 20993 14059 21051 14065
rect 20993 14025 21005 14059
rect 21039 14056 21051 14059
rect 22002 14056 22008 14068
rect 21039 14028 22008 14056
rect 21039 14025 21051 14028
rect 20993 14019 21051 14025
rect 22002 14016 22008 14028
rect 22060 14016 22066 14068
rect 9953 13991 10011 13997
rect 8588 13960 8694 13988
rect 9953 13957 9965 13991
rect 9999 13988 10011 13991
rect 10778 13988 10784 14000
rect 9999 13960 10784 13988
rect 9999 13957 10011 13960
rect 9953 13951 10011 13957
rect 10778 13948 10784 13960
rect 10836 13948 10842 14000
rect 12253 13991 12311 13997
rect 12253 13957 12265 13991
rect 12299 13988 12311 13991
rect 15286 13988 15292 14000
rect 12299 13960 15292 13988
rect 12299 13957 12311 13960
rect 12253 13951 12311 13957
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 15746 13948 15752 14000
rect 15804 13988 15810 14000
rect 16209 13991 16267 13997
rect 16209 13988 16221 13991
rect 15804 13960 16221 13988
rect 15804 13948 15810 13960
rect 16209 13957 16221 13960
rect 16255 13957 16267 13991
rect 16209 13951 16267 13957
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 17920 13960 18337 13988
rect 17920 13948 17926 13960
rect 18325 13957 18337 13960
rect 18371 13957 18383 13991
rect 18325 13951 18383 13957
rect 20625 13991 20683 13997
rect 20625 13957 20637 13991
rect 20671 13988 20683 13991
rect 23293 13991 23351 13997
rect 23293 13988 23305 13991
rect 20671 13960 23305 13988
rect 20671 13957 20683 13960
rect 20625 13951 20683 13957
rect 23293 13957 23305 13960
rect 23339 13957 23351 13991
rect 23293 13951 23351 13957
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 13354 13920 13360 13932
rect 12207 13892 13360 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13920 13507 13923
rect 14274 13920 14280 13932
rect 13495 13892 14280 13920
rect 13495 13889 13507 13892
rect 13449 13883 13507 13889
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 14366 13880 14372 13932
rect 14424 13880 14430 13932
rect 18782 13880 18788 13932
rect 18840 13880 18846 13932
rect 22094 13880 22100 13932
rect 22152 13920 22158 13932
rect 22830 13920 22836 13932
rect 22152 13892 22836 13920
rect 22152 13880 22158 13892
rect 22830 13880 22836 13892
rect 22888 13880 22894 13932
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 23532 13892 23949 13920
rect 23532 13880 23538 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 934 13812 940 13864
rect 992 13852 998 13864
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 992 13824 1777 13852
rect 992 13812 998 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 8202 13812 8208 13864
rect 8260 13812 8266 13864
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 8938 13852 8944 13864
rect 8812 13824 8944 13852
rect 8812 13812 8818 13824
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 12345 13855 12403 13861
rect 12345 13852 12357 13855
rect 11624 13824 12357 13852
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 11624 13784 11652 13824
rect 12345 13821 12357 13824
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 9456 13756 11652 13784
rect 9456 13744 9462 13756
rect 11698 13744 11704 13796
rect 11756 13784 11762 13796
rect 13556 13784 13584 13815
rect 14182 13812 14188 13864
rect 14240 13812 14246 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15562 13852 15568 13864
rect 15335 13824 15568 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15896 13824 15945 13852
rect 15896 13812 15902 13824
rect 15933 13821 15945 13824
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13852 18107 13855
rect 18322 13852 18328 13864
rect 18095 13824 18328 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 11756 13756 13584 13784
rect 11756 13744 11762 13756
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 19334 13784 19340 13796
rect 14700 13756 19340 13784
rect 14700 13744 14706 13756
rect 19334 13744 19340 13756
rect 19392 13744 19398 13796
rect 20456 13784 20484 13815
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 22189 13855 22247 13861
rect 22189 13852 22201 13855
rect 21508 13824 22201 13852
rect 21508 13812 21514 13824
rect 22189 13821 22201 13824
rect 22235 13821 22247 13855
rect 22189 13815 22247 13821
rect 20714 13784 20720 13796
rect 20456 13756 20720 13784
rect 20714 13744 20720 13756
rect 20772 13744 20778 13796
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 14734 13716 14740 13728
rect 10560 13688 14740 13716
rect 10560 13676 10566 13688
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 16114 13676 16120 13728
rect 16172 13716 16178 13728
rect 19518 13716 19524 13728
rect 16172 13688 19524 13716
rect 16172 13676 16178 13688
rect 19518 13676 19524 13688
rect 19576 13716 19582 13728
rect 19794 13716 19800 13728
rect 19576 13688 19800 13716
rect 19576 13676 19582 13688
rect 19794 13676 19800 13688
rect 19852 13676 19858 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 9769 13515 9827 13521
rect 9769 13512 9781 13515
rect 8260 13484 9781 13512
rect 8260 13472 8266 13484
rect 9769 13481 9781 13484
rect 9815 13481 9827 13515
rect 9769 13475 9827 13481
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 11112 13484 12265 13512
rect 11112 13472 11118 13484
rect 12253 13481 12265 13484
rect 12299 13512 12311 13515
rect 14185 13515 14243 13521
rect 12299 13484 12434 13512
rect 12299 13481 12311 13484
rect 12253 13475 12311 13481
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8536 13280 9137 13308
rect 8536 13268 8542 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 12406 13308 12434 13484
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 14366 13512 14372 13524
rect 14231 13484 14372 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 15197 13515 15255 13521
rect 15197 13481 15209 13515
rect 15243 13512 15255 13515
rect 17770 13512 17776 13524
rect 15243 13484 17776 13512
rect 15243 13481 15255 13484
rect 15197 13475 15255 13481
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 20990 13472 20996 13524
rect 21048 13512 21054 13524
rect 22281 13515 22339 13521
rect 22281 13512 22293 13515
rect 21048 13484 22293 13512
rect 21048 13472 21054 13484
rect 22281 13481 22293 13484
rect 22327 13481 22339 13515
rect 22281 13475 22339 13481
rect 13357 13447 13415 13453
rect 13357 13413 13369 13447
rect 13403 13444 13415 13447
rect 15378 13444 15384 13456
rect 13403 13416 15384 13444
rect 13403 13413 13415 13416
rect 13357 13407 13415 13413
rect 15378 13404 15384 13416
rect 15436 13404 15442 13456
rect 17402 13444 17408 13456
rect 17236 13416 17408 13444
rect 12710 13336 12716 13388
rect 12768 13336 12774 13388
rect 12894 13336 12900 13388
rect 12952 13376 12958 13388
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 12952 13348 13645 13376
rect 12952 13336 12958 13348
rect 13633 13345 13645 13348
rect 13679 13376 13691 13379
rect 13722 13376 13728 13388
rect 13679 13348 13728 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 14918 13376 14924 13388
rect 14424 13348 14924 13376
rect 14424 13336 14430 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 12406 13280 13001 13308
rect 9125 13271 9183 13277
rect 12989 13277 13001 13280
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 13998 13308 14004 13320
rect 13955 13280 14004 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 13998 13268 14004 13280
rect 14056 13308 14062 13320
rect 14642 13308 14648 13320
rect 14056 13280 14648 13308
rect 14056 13268 14062 13280
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13308 17003 13311
rect 17236 13308 17264 13416
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 17310 13336 17316 13388
rect 17368 13376 17374 13388
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 17368 13348 19257 13376
rect 17368 13336 17374 13348
rect 16991 13280 17264 13308
rect 17405 13311 17463 13317
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 17405 13277 17417 13311
rect 17451 13308 17463 13311
rect 17494 13308 17500 13320
rect 17451 13280 17500 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 18616 13317 18644 13348
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 22370 13376 22376 13388
rect 19245 13339 19303 13345
rect 22066 13348 22376 13376
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13308 18843 13311
rect 20714 13308 20720 13320
rect 18831 13280 20720 13308
rect 18831 13277 18843 13280
rect 18785 13271 18843 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 20898 13268 20904 13320
rect 20956 13308 20962 13320
rect 21821 13311 21879 13317
rect 21821 13308 21833 13311
rect 20956 13280 21833 13308
rect 20956 13268 20962 13280
rect 21821 13277 21833 13280
rect 21867 13308 21879 13311
rect 22066 13308 22094 13348
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 21867 13280 22094 13308
rect 21867 13277 21879 13280
rect 21821 13271 21879 13277
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22649 13311 22707 13317
rect 22649 13308 22661 13311
rect 22244 13280 22661 13308
rect 22244 13268 22250 13280
rect 22649 13277 22661 13280
rect 22695 13277 22707 13311
rect 22649 13271 22707 13277
rect 16669 13243 16727 13249
rect 16238 13212 16528 13240
rect 16500 13184 16528 13212
rect 16669 13209 16681 13243
rect 16715 13240 16727 13243
rect 18049 13243 18107 13249
rect 18049 13240 18061 13243
rect 16715 13212 18061 13240
rect 16715 13209 16727 13212
rect 16669 13203 16727 13209
rect 18049 13209 18061 13212
rect 18095 13209 18107 13243
rect 18049 13203 18107 13209
rect 19150 13200 19156 13252
rect 19208 13240 19214 13252
rect 20165 13243 20223 13249
rect 20165 13240 20177 13243
rect 19208 13212 20177 13240
rect 19208 13200 19214 13212
rect 20165 13209 20177 13212
rect 20211 13209 20223 13243
rect 20165 13203 20223 13209
rect 16482 13132 16488 13184
rect 16540 13132 16546 13184
rect 20180 13172 20208 13203
rect 20346 13200 20352 13252
rect 20404 13200 20410 13252
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 21085 13243 21143 13249
rect 21085 13240 21097 13243
rect 21048 13212 21097 13240
rect 21048 13200 21054 13212
rect 21085 13209 21097 13212
rect 21131 13209 21143 13243
rect 21085 13203 21143 13209
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 25498 13240 25504 13252
rect 23891 13212 25504 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 25498 13200 25504 13212
rect 25556 13200 25562 13252
rect 20625 13175 20683 13181
rect 20625 13172 20637 13175
rect 20180 13144 20637 13172
rect 20625 13141 20637 13144
rect 20671 13141 20683 13175
rect 20625 13135 20683 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 11238 12928 11244 12980
rect 11296 12928 11302 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12216 12940 12434 12968
rect 12216 12928 12222 12940
rect 12406 12900 12434 12940
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 14001 12971 14059 12977
rect 14001 12968 14013 12971
rect 13412 12940 14013 12968
rect 13412 12928 13418 12940
rect 14001 12937 14013 12940
rect 14047 12937 14059 12971
rect 14001 12931 14059 12937
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 15194 12968 15200 12980
rect 14415 12940 15200 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 15194 12928 15200 12940
rect 15252 12968 15258 12980
rect 15470 12968 15476 12980
rect 15252 12940 15476 12968
rect 15252 12928 15258 12940
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 17184 12940 17233 12968
rect 17184 12928 17190 12940
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 17221 12931 17279 12937
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 18782 12968 18788 12980
rect 18187 12940 18788 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 21726 12928 21732 12980
rect 21784 12968 21790 12980
rect 22281 12971 22339 12977
rect 22281 12968 22293 12971
rect 21784 12940 22293 12968
rect 21784 12928 21790 12940
rect 22281 12937 22293 12940
rect 22327 12937 22339 12971
rect 22281 12931 22339 12937
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 12406 12872 12633 12900
rect 12621 12869 12633 12872
rect 12667 12869 12679 12903
rect 12621 12863 12679 12869
rect 14461 12903 14519 12909
rect 14461 12869 14473 12903
rect 14507 12900 14519 12903
rect 14642 12900 14648 12912
rect 14507 12872 14648 12900
rect 14507 12869 14519 12872
rect 14461 12863 14519 12869
rect 14642 12860 14648 12872
rect 14700 12860 14706 12912
rect 15562 12860 15568 12912
rect 15620 12900 15626 12912
rect 16025 12903 16083 12909
rect 16025 12900 16037 12903
rect 15620 12872 16037 12900
rect 15620 12860 15626 12872
rect 16025 12869 16037 12872
rect 16071 12869 16083 12903
rect 19518 12900 19524 12912
rect 19182 12872 19524 12900
rect 16025 12863 16083 12869
rect 19518 12860 19524 12872
rect 19576 12900 19582 12912
rect 20165 12903 20223 12909
rect 20165 12900 20177 12903
rect 19576 12872 20177 12900
rect 19576 12860 19582 12872
rect 20165 12869 20177 12872
rect 20211 12869 20223 12903
rect 20165 12863 20223 12869
rect 20717 12903 20775 12909
rect 20717 12869 20729 12903
rect 20763 12900 20775 12903
rect 21361 12903 21419 12909
rect 21361 12900 21373 12903
rect 20763 12872 21373 12900
rect 20763 12869 20775 12872
rect 20717 12863 20775 12869
rect 21361 12869 21373 12872
rect 21407 12900 21419 12903
rect 24210 12900 24216 12912
rect 21407 12872 24216 12900
rect 21407 12869 21419 12872
rect 21361 12863 21419 12869
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12832 13415 12835
rect 14366 12832 14372 12844
rect 13403 12804 14372 12832
rect 13403 12801 13415 12804
rect 13357 12795 13415 12801
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 16390 12792 16396 12844
rect 16448 12832 16454 12844
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 16448 12804 17141 12832
rect 16448 12792 16454 12804
rect 17129 12801 17141 12804
rect 17175 12801 17187 12835
rect 20180 12832 20208 12863
rect 24210 12860 24216 12872
rect 24268 12900 24274 12912
rect 24578 12900 24584 12912
rect 24268 12872 24584 12900
rect 24268 12860 24274 12872
rect 24578 12860 24584 12872
rect 24636 12860 24642 12912
rect 20990 12832 20996 12844
rect 20180 12804 20996 12832
rect 17129 12795 17187 12801
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 22370 12792 22376 12844
rect 22428 12792 22434 12844
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12832 23259 12835
rect 23290 12832 23296 12844
rect 23247 12804 23296 12832
rect 23247 12801 23259 12804
rect 23201 12795 23259 12801
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 23440 12804 23949 12832
rect 23440 12792 23446 12804
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 10778 12724 10784 12776
rect 10836 12764 10842 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 10836 12736 14657 12764
rect 10836 12724 10842 12736
rect 14645 12733 14657 12736
rect 14691 12764 14703 12767
rect 15562 12764 15568 12776
rect 14691 12736 15568 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12764 17095 12767
rect 17770 12764 17776 12776
rect 17083 12736 17776 12764
rect 17083 12733 17095 12736
rect 17037 12727 17095 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12764 19671 12767
rect 19889 12767 19947 12773
rect 19659 12736 19840 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 12802 12656 12808 12708
rect 12860 12656 12866 12708
rect 15749 12699 15807 12705
rect 15749 12665 15761 12699
rect 15795 12696 15807 12699
rect 16850 12696 16856 12708
rect 15795 12668 16856 12696
rect 15795 12665 15807 12668
rect 15749 12659 15807 12665
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 18046 12696 18052 12708
rect 17512 12668 18052 12696
rect 13446 12588 13452 12640
rect 13504 12588 13510 12640
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 17512 12628 17540 12668
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 19812 12696 19840 12736
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 21082 12764 21088 12776
rect 19935 12736 21088 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 21082 12724 21088 12736
rect 21140 12764 21146 12776
rect 21140 12736 21404 12764
rect 21140 12724 21146 12736
rect 21376 12708 21404 12736
rect 22094 12724 22100 12776
rect 22152 12724 22158 12776
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 20990 12696 20996 12708
rect 19812 12668 20996 12696
rect 20990 12656 20996 12668
rect 21048 12656 21054 12708
rect 21358 12656 21364 12708
rect 21416 12656 21422 12708
rect 22830 12656 22836 12708
rect 22888 12696 22894 12708
rect 23385 12699 23443 12705
rect 23385 12696 23397 12699
rect 22888 12668 23397 12696
rect 22888 12656 22894 12668
rect 23385 12665 23397 12668
rect 23431 12665 23443 12699
rect 23385 12659 23443 12665
rect 13780 12600 17540 12628
rect 17589 12631 17647 12637
rect 13780 12588 13786 12600
rect 17589 12597 17601 12631
rect 17635 12628 17647 12631
rect 20438 12628 20444 12640
rect 17635 12600 20444 12628
rect 17635 12597 17647 12600
rect 17589 12591 17647 12597
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 22741 12631 22799 12637
rect 22741 12597 22753 12631
rect 22787 12628 22799 12631
rect 23290 12628 23296 12640
rect 22787 12600 23296 12628
rect 22787 12597 22799 12600
rect 22741 12591 22799 12597
rect 23290 12588 23296 12600
rect 23348 12588 23354 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 16022 12384 16028 12436
rect 16080 12384 16086 12436
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 5902 12356 5908 12368
rect 2832 12328 5908 12356
rect 2832 12316 2838 12328
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 19889 12359 19947 12365
rect 19889 12356 19901 12359
rect 17972 12328 19901 12356
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 8352 12260 9413 12288
rect 8352 12248 8358 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 11238 12288 11244 12300
rect 10796 12260 11244 12288
rect 10796 12206 10824 12260
rect 11238 12248 11244 12260
rect 11296 12288 11302 12300
rect 11296 12260 11744 12288
rect 11296 12248 11302 12260
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11164 12192 11621 12220
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 11164 12093 11192 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11716 12220 11744 12260
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 17972 12297 18000 12328
rect 19889 12325 19901 12328
rect 19935 12356 19947 12359
rect 20070 12356 20076 12368
rect 19935 12328 20076 12356
rect 19935 12325 19947 12328
rect 19889 12319 19947 12325
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 23385 12359 23443 12365
rect 23385 12325 23397 12359
rect 23431 12356 23443 12359
rect 25038 12356 25044 12368
rect 23431 12328 25044 12356
rect 23431 12325 23443 12328
rect 23385 12319 23443 12325
rect 25038 12316 25044 12328
rect 25096 12316 25102 12368
rect 14277 12291 14335 12297
rect 14277 12288 14289 12291
rect 12216 12260 14289 12288
rect 12216 12248 12222 12260
rect 14277 12257 14289 12260
rect 14323 12257 14335 12291
rect 14277 12251 14335 12257
rect 17957 12291 18015 12297
rect 17957 12257 17969 12291
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18104 12260 18797 12288
rect 18104 12248 18110 12260
rect 18785 12257 18797 12260
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 21637 12291 21695 12297
rect 21637 12288 21649 12291
rect 21416 12260 21649 12288
rect 21416 12248 21422 12260
rect 21637 12257 21649 12260
rect 21683 12257 21695 12291
rect 21637 12251 21695 12257
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12288 22339 12291
rect 22370 12288 22376 12300
rect 22327 12260 22376 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 22370 12248 22376 12260
rect 22428 12248 22434 12300
rect 22646 12248 22652 12300
rect 22704 12288 22710 12300
rect 22704 12260 23888 12288
rect 22704 12248 22710 12260
rect 12250 12220 12256 12232
rect 11716 12192 12256 12220
rect 11609 12183 11667 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 13722 12180 13728 12232
rect 13780 12180 13786 12232
rect 15654 12180 15660 12232
rect 15712 12220 15718 12232
rect 16482 12220 16488 12232
rect 15712 12192 16488 12220
rect 15712 12180 15718 12192
rect 16482 12180 16488 12192
rect 16540 12220 16546 12232
rect 18874 12220 18880 12232
rect 16540 12192 18880 12220
rect 16540 12180 16546 12192
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 21726 12180 21732 12232
rect 21784 12220 21790 12232
rect 23860 12229 23888 12260
rect 23201 12223 23259 12229
rect 23201 12220 23213 12223
rect 21784 12192 23213 12220
rect 21784 12180 21790 12192
rect 23201 12189 23213 12192
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 13081 12155 13139 12161
rect 13081 12121 13093 12155
rect 13127 12152 13139 12155
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 13127 12124 14565 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 14553 12121 14565 12124
rect 14599 12121 14611 12155
rect 14553 12115 14611 12121
rect 17310 12112 17316 12164
rect 17368 12152 17374 12164
rect 18141 12155 18199 12161
rect 18141 12152 18153 12155
rect 17368 12124 18153 12152
rect 17368 12112 17374 12124
rect 18141 12121 18153 12124
rect 18187 12121 18199 12155
rect 18141 12115 18199 12121
rect 20898 12112 20904 12164
rect 20956 12112 20962 12164
rect 21361 12155 21419 12161
rect 21361 12121 21373 12155
rect 21407 12152 21419 12155
rect 21450 12152 21456 12164
rect 21407 12124 21456 12152
rect 21407 12121 21419 12124
rect 21361 12115 21419 12121
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10652 12056 11161 12084
rect 10652 12044 10658 12056
rect 11149 12053 11161 12056
rect 11195 12053 11207 12087
rect 11149 12047 11207 12053
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 11296 12056 12265 12084
rect 11296 12044 11302 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 18509 12087 18567 12093
rect 18509 12053 18521 12087
rect 18555 12084 18567 12087
rect 19518 12084 19524 12096
rect 18555 12056 19524 12084
rect 18555 12053 18567 12056
rect 18509 12047 18567 12053
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 24029 12087 24087 12093
rect 24029 12053 24041 12087
rect 24075 12084 24087 12087
rect 24854 12084 24860 12096
rect 24075 12056 24860 12084
rect 24075 12053 24087 12056
rect 24029 12047 24087 12053
rect 24854 12044 24860 12056
rect 24912 12044 24918 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 9916 11852 10701 11880
rect 9916 11840 9922 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12032 11852 13768 11880
rect 12032 11840 12038 11852
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 7892 11716 10793 11744
rect 7892 11704 7898 11716
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11422 11744 11428 11756
rect 11112 11716 11428 11744
rect 11112 11704 11118 11716
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 13740 11744 13768 11852
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 16853 11883 16911 11889
rect 16853 11880 16865 11883
rect 14332 11852 16865 11880
rect 14332 11840 14338 11852
rect 16853 11849 16865 11852
rect 16899 11849 16911 11883
rect 16853 11843 16911 11849
rect 17221 11883 17279 11889
rect 17221 11849 17233 11883
rect 17267 11880 17279 11883
rect 19702 11880 19708 11892
rect 17267 11852 19708 11880
rect 17267 11849 17279 11852
rect 17221 11843 17279 11849
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 20990 11840 20996 11892
rect 21048 11840 21054 11892
rect 15289 11815 15347 11821
rect 15289 11781 15301 11815
rect 15335 11812 15347 11815
rect 15654 11812 15660 11824
rect 15335 11784 15660 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 15654 11772 15660 11784
rect 15712 11772 15718 11824
rect 15841 11815 15899 11821
rect 15841 11781 15853 11815
rect 15887 11812 15899 11815
rect 16301 11815 16359 11821
rect 16301 11812 16313 11815
rect 15887 11784 16313 11812
rect 15887 11781 15899 11784
rect 15841 11775 15899 11781
rect 16301 11781 16313 11784
rect 16347 11781 16359 11815
rect 16301 11775 16359 11781
rect 15856 11744 15884 11775
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 17000 11784 17448 11812
rect 17000 11772 17006 11784
rect 10594 11636 10600 11688
rect 10652 11636 10658 11688
rect 12158 11636 12164 11688
rect 12216 11636 12222 11688
rect 12434 11636 12440 11688
rect 12492 11636 12498 11688
rect 13556 11676 13584 11730
rect 13740 11716 15884 11744
rect 13906 11676 13912 11688
rect 13556 11648 13912 11676
rect 13906 11636 13912 11648
rect 13964 11676 13970 11688
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 13964 11648 14473 11676
rect 13964 11636 13970 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 17310 11636 17316 11688
rect 17368 11636 17374 11688
rect 17420 11685 17448 11784
rect 18874 11772 18880 11824
rect 18932 11772 18938 11824
rect 20530 11772 20536 11824
rect 20588 11812 20594 11824
rect 21269 11815 21327 11821
rect 21269 11812 21281 11815
rect 20588 11784 21281 11812
rect 20588 11772 20594 11784
rect 21269 11781 21281 11784
rect 21315 11781 21327 11815
rect 21269 11775 21327 11781
rect 22094 11772 22100 11824
rect 22152 11812 22158 11824
rect 23201 11815 23259 11821
rect 23201 11812 23213 11815
rect 22152 11784 23213 11812
rect 22152 11772 22158 11784
rect 23201 11781 23213 11784
rect 23247 11781 23259 11815
rect 23201 11775 23259 11781
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 18141 11747 18199 11753
rect 18141 11744 18153 11747
rect 17552 11716 18153 11744
rect 17552 11704 17558 11716
rect 18141 11713 18153 11716
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 19944 11716 20361 11744
rect 19944 11704 19950 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 21174 11704 21180 11756
rect 21232 11744 21238 11756
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 21232 11716 22753 11744
rect 21232 11704 21238 11716
rect 22741 11713 22753 11716
rect 22787 11713 22799 11747
rect 22741 11707 22799 11713
rect 23842 11704 23848 11756
rect 23900 11744 23906 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23900 11716 23949 11744
rect 23900 11704 23906 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 19426 11676 19432 11688
rect 18463 11648 19432 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 16025 11611 16083 11617
rect 16025 11577 16037 11611
rect 16071 11608 16083 11611
rect 16482 11608 16488 11620
rect 16071 11580 16488 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 22281 11611 22339 11617
rect 22281 11577 22293 11611
rect 22327 11608 22339 11611
rect 22554 11608 22560 11620
rect 22327 11580 22560 11608
rect 22327 11577 22339 11580
rect 22281 11571 22339 11577
rect 22554 11568 22560 11580
rect 22612 11568 22618 11620
rect 22925 11611 22983 11617
rect 22925 11577 22937 11611
rect 22971 11608 22983 11611
rect 23382 11608 23388 11620
rect 22971 11580 23388 11608
rect 22971 11577 22983 11580
rect 22925 11571 22983 11577
rect 23382 11568 23388 11580
rect 23440 11568 23446 11620
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 13538 11540 13544 11552
rect 11195 11512 13544 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13780 11512 13921 11540
rect 13780 11500 13786 11512
rect 13909 11509 13921 11512
rect 13955 11540 13967 11543
rect 15194 11540 15200 11552
rect 13955 11512 15200 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 19886 11500 19892 11552
rect 19944 11500 19950 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12492 11308 12909 11336
rect 12492 11296 12498 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13906 11336 13912 11348
rect 13044 11308 13912 11336
rect 13044 11296 13050 11308
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 15197 11339 15255 11345
rect 15197 11305 15209 11339
rect 15243 11336 15255 11339
rect 15286 11336 15292 11348
rect 15243 11308 15292 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 18969 11339 19027 11345
rect 18969 11305 18981 11339
rect 19015 11336 19027 11339
rect 19058 11336 19064 11348
rect 19015 11308 19064 11336
rect 19015 11305 19027 11308
rect 18969 11299 19027 11305
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 19426 11296 19432 11348
rect 19484 11296 19490 11348
rect 12526 11228 12532 11280
rect 12584 11268 12590 11280
rect 14829 11271 14887 11277
rect 14829 11268 14841 11271
rect 12584 11240 14841 11268
rect 12584 11228 12590 11240
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11200 10747 11203
rect 12158 11200 12164 11212
rect 10735 11172 12164 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 12710 11200 12716 11212
rect 12483 11172 12716 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 12710 11160 12716 11172
rect 12768 11200 12774 11212
rect 12768 11172 13584 11200
rect 12768 11160 12774 11172
rect 13556 11141 13584 11172
rect 14476 11141 14504 11240
rect 14829 11237 14841 11240
rect 14875 11237 14887 11271
rect 20622 11268 20628 11280
rect 14829 11231 14887 11237
rect 15580 11240 20628 11268
rect 15580 11141 15608 11240
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 15749 11203 15807 11209
rect 15749 11200 15761 11203
rect 15712 11172 15761 11200
rect 15712 11160 15718 11172
rect 15749 11169 15761 11172
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 20864 11172 21404 11200
rect 20864 11160 20870 11172
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11132 18475 11135
rect 19058 11132 19064 11144
rect 18463 11104 19064 11132
rect 18463 11101 18475 11104
rect 18417 11095 18475 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 20070 11092 20076 11144
rect 20128 11092 20134 11144
rect 20530 11092 20536 11144
rect 20588 11132 20594 11144
rect 21376 11141 21404 11172
rect 20625 11135 20683 11141
rect 20625 11132 20637 11135
rect 20588 11104 20637 11132
rect 20588 11092 20594 11104
rect 20625 11101 20637 11104
rect 20671 11101 20683 11135
rect 20625 11095 20683 11101
rect 21361 11135 21419 11141
rect 21361 11101 21373 11135
rect 21407 11132 21419 11135
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 21407 11104 21833 11132
rect 21407 11101 21419 11104
rect 21361 11095 21419 11101
rect 21821 11101 21833 11104
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 10965 11067 11023 11073
rect 10965 11033 10977 11067
rect 11011 11064 11023 11067
rect 11238 11064 11244 11076
rect 11011 11036 11244 11064
rect 11011 11033 11023 11036
rect 10965 11027 11023 11033
rect 11238 11024 11244 11036
rect 11296 11024 11302 11076
rect 12250 11064 12256 11076
rect 12190 11036 12256 11064
rect 12250 11024 12256 11036
rect 12308 11064 12314 11076
rect 12986 11064 12992 11076
rect 12308 11036 12992 11064
rect 12308 11024 12314 11036
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 14274 11024 14280 11076
rect 14332 11024 14338 11076
rect 15657 11067 15715 11073
rect 15657 11033 15669 11067
rect 15703 11064 15715 11067
rect 16114 11064 16120 11076
rect 15703 11036 16120 11064
rect 15703 11033 15715 11036
rect 15657 11027 15715 11033
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 15672 10996 15700 11027
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 18601 11067 18659 11073
rect 18601 11033 18613 11067
rect 18647 11064 18659 11067
rect 19610 11064 19616 11076
rect 18647 11036 19616 11064
rect 18647 11033 18659 11036
rect 18601 11027 18659 11033
rect 19610 11024 19616 11036
rect 19668 11024 19674 11076
rect 20809 11067 20867 11073
rect 20809 11033 20821 11067
rect 20855 11064 20867 11067
rect 21266 11064 21272 11076
rect 20855 11036 21272 11064
rect 20855 11033 20867 11036
rect 20809 11027 20867 11033
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 21542 11024 21548 11076
rect 21600 11024 21606 11076
rect 15620 10968 15700 10996
rect 15620 10956 15626 10968
rect 16390 10956 16396 11008
rect 16448 10956 16454 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 10008 10764 11529 10792
rect 10008 10752 10014 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 12621 10795 12679 10801
rect 12621 10761 12633 10795
rect 12667 10792 12679 10795
rect 12986 10792 12992 10804
rect 12667 10764 12992 10792
rect 12667 10761 12679 10764
rect 12621 10755 12679 10761
rect 11532 10724 11560 10755
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 15562 10792 15568 10804
rect 14568 10764 15568 10792
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 11532 10696 11989 10724
rect 11977 10693 11989 10696
rect 12023 10693 12035 10727
rect 11977 10687 12035 10693
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 14568 10597 14596 10764
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 15657 10795 15715 10801
rect 15657 10761 15669 10795
rect 15703 10792 15715 10795
rect 15703 10764 16574 10792
rect 15703 10761 15715 10764
rect 15657 10755 15715 10761
rect 15194 10684 15200 10736
rect 15252 10684 15258 10736
rect 15289 10727 15347 10733
rect 15289 10693 15301 10727
rect 15335 10724 15347 10727
rect 16390 10724 16396 10736
rect 15335 10696 16396 10724
rect 15335 10693 15347 10696
rect 15289 10687 15347 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 15212 10656 15240 10684
rect 15120 10628 15240 10656
rect 16117 10659 16175 10665
rect 15120 10597 15148 10628
rect 16117 10625 16129 10659
rect 16163 10625 16175 10659
rect 16546 10656 16574 10764
rect 19518 10752 19524 10804
rect 19576 10752 19582 10804
rect 20625 10795 20683 10801
rect 20625 10761 20637 10795
rect 20671 10792 20683 10795
rect 20671 10764 22140 10792
rect 20671 10761 20683 10764
rect 20625 10755 20683 10761
rect 19613 10727 19671 10733
rect 19613 10693 19625 10727
rect 19659 10724 19671 10727
rect 21085 10727 21143 10733
rect 21085 10724 21097 10727
rect 19659 10696 21097 10724
rect 19659 10693 19671 10696
rect 19613 10687 19671 10693
rect 21085 10693 21097 10696
rect 21131 10693 21143 10727
rect 21085 10687 21143 10693
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 16546 10628 18613 10656
rect 16117 10619 16175 10625
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 19886 10656 19892 10668
rect 18601 10619 18659 10625
rect 19444 10628 19892 10656
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 12032 10560 14565 10588
rect 12032 10548 12038 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10588 15255 10591
rect 15378 10588 15384 10600
rect 15243 10560 15384 10588
rect 15243 10557 15255 10560
rect 15197 10551 15255 10557
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 16132 10520 16160 10619
rect 19444 10597 19472 10628
rect 19886 10616 19892 10628
rect 19944 10616 19950 10668
rect 20438 10616 20444 10668
rect 20496 10616 20502 10668
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10625 22063 10659
rect 22112 10656 22140 10764
rect 23293 10659 23351 10665
rect 23293 10656 23305 10659
rect 22112 10628 23305 10656
rect 22005 10619 22063 10625
rect 23293 10625 23305 10628
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 19429 10591 19487 10597
rect 19429 10557 19441 10591
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 13596 10492 16160 10520
rect 16301 10523 16359 10529
rect 13596 10480 13602 10492
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 22020 10520 22048 10619
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 16347 10492 22048 10520
rect 22189 10523 22247 10529
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 22189 10489 22201 10523
rect 22235 10520 22247 10523
rect 23934 10520 23940 10532
rect 22235 10492 23940 10520
rect 22235 10489 22247 10492
rect 22189 10483 22247 10489
rect 23934 10480 23940 10492
rect 23992 10480 23998 10532
rect 12066 10412 12072 10464
rect 12124 10412 12130 10464
rect 18785 10455 18843 10461
rect 18785 10421 18797 10455
rect 18831 10452 18843 10455
rect 19886 10452 19892 10464
rect 18831 10424 19892 10452
rect 18831 10421 18843 10424
rect 18785 10415 18843 10421
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 19981 10455 20039 10461
rect 19981 10421 19993 10455
rect 20027 10452 20039 10455
rect 21450 10452 21456 10464
rect 20027 10424 21456 10452
rect 20027 10421 20039 10424
rect 19981 10415 20039 10421
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 23474 10412 23480 10464
rect 23532 10412 23538 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 18966 10044 18972 10056
rect 16899 10016 18972 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 22002 10004 22008 10056
rect 22060 10004 22066 10056
rect 22830 10004 22836 10056
rect 22888 10004 22894 10056
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 24946 10044 24952 10056
rect 23891 10016 24952 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 17034 9936 17040 9988
rect 17092 9936 17098 9988
rect 22922 9936 22928 9988
rect 22980 9976 22986 9988
rect 24765 9979 24823 9985
rect 24765 9976 24777 9979
rect 22980 9948 24777 9976
rect 22980 9936 22986 9948
rect 24765 9945 24777 9948
rect 24811 9945 24823 9979
rect 24765 9939 24823 9945
rect 22186 9868 22192 9920
rect 22244 9868 22250 9920
rect 23198 9868 23204 9920
rect 23256 9908 23262 9920
rect 24673 9911 24731 9917
rect 24673 9908 24685 9911
rect 23256 9880 24685 9908
rect 23256 9868 23262 9880
rect 24673 9877 24685 9880
rect 24719 9877 24731 9911
rect 24673 9871 24731 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 22830 9664 22836 9716
rect 22888 9664 22894 9716
rect 12618 9596 12624 9648
rect 12676 9636 12682 9648
rect 14553 9639 14611 9645
rect 14553 9636 14565 9639
rect 12676 9608 14565 9636
rect 12676 9596 12682 9608
rect 14553 9605 14565 9608
rect 14599 9605 14611 9639
rect 14553 9599 14611 9605
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 13722 9568 13728 9580
rect 13504 9540 13728 9568
rect 13504 9528 13510 9540
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 19944 9540 22661 9568
rect 19944 9528 19950 9540
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 23290 9528 23296 9580
rect 23348 9528 23354 9580
rect 23934 9528 23940 9580
rect 23992 9528 23998 9580
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 5718 9500 5724 9512
rect 2924 9472 5724 9500
rect 2924 9460 2930 9472
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 14645 9367 14703 9373
rect 14645 9333 14657 9367
rect 14691 9364 14703 9367
rect 19426 9364 19432 9376
rect 14691 9336 19432 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 24578 9364 24584 9376
rect 23523 9336 24584 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 24578 9324 24584 9336
rect 24636 9324 24642 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8956 16635 8959
rect 16758 8956 16764 8968
rect 16623 8928 16764 8956
rect 16623 8925 16635 8928
rect 16577 8919 16635 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 19521 8959 19579 8965
rect 19521 8925 19533 8959
rect 19567 8956 19579 8959
rect 20346 8956 20352 8968
rect 19567 8928 20352 8956
rect 19567 8925 19579 8928
rect 19521 8919 19579 8925
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 23382 8916 23388 8968
rect 23440 8956 23446 8968
rect 23753 8959 23811 8965
rect 23753 8956 23765 8959
rect 23440 8928 23765 8956
rect 23440 8916 23446 8928
rect 23753 8925 23765 8928
rect 23799 8925 23811 8959
rect 23753 8919 23811 8925
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8956 24915 8959
rect 25038 8956 25044 8968
rect 24903 8928 25044 8956
rect 24903 8925 24915 8928
rect 24857 8919 24915 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 19705 8891 19763 8897
rect 19705 8857 19717 8891
rect 19751 8888 19763 8891
rect 21818 8888 21824 8900
rect 19751 8860 21824 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 7800 8792 7849 8820
rect 7800 8780 7806 8792
rect 7837 8789 7849 8792
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 16669 8823 16727 8829
rect 16669 8789 16681 8823
rect 16715 8820 16727 8823
rect 17770 8820 17776 8832
rect 16715 8792 17776 8820
rect 16715 8789 16727 8792
rect 16669 8783 16727 8789
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 23934 8780 23940 8832
rect 23992 8780 23998 8832
rect 24026 8780 24032 8832
rect 24084 8820 24090 8832
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 24084 8792 24685 8820
rect 24084 8780 24090 8792
rect 24673 8789 24685 8792
rect 24719 8789 24731 8823
rect 24673 8783 24731 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 7742 8576 7748 8628
rect 7800 8576 7806 8628
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 7892 8588 8125 8616
rect 7892 8576 7898 8588
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 8113 8579 8171 8585
rect 20901 8551 20959 8557
rect 20901 8517 20913 8551
rect 20947 8548 20959 8551
rect 21910 8548 21916 8560
rect 20947 8520 21916 8548
rect 20947 8517 20959 8520
rect 20901 8511 20959 8517
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 5592 8452 7665 8480
rect 5592 8440 5598 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 11514 8412 11520 8424
rect 7607 8384 11520 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 21545 8415 21603 8421
rect 21545 8412 21557 8415
rect 11940 8384 21557 8412
rect 11940 8372 11946 8384
rect 21545 8381 21557 8384
rect 21591 8412 21603 8415
rect 22112 8412 22140 8443
rect 23474 8440 23480 8492
rect 23532 8480 23538 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23532 8452 23949 8480
rect 23532 8440 23538 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 21591 8384 22140 8412
rect 21591 8381 21603 8384
rect 21545 8375 21603 8381
rect 22646 8372 22652 8424
rect 22704 8372 22710 8424
rect 20717 8347 20775 8353
rect 20717 8313 20729 8347
rect 20763 8344 20775 8347
rect 20990 8344 20996 8356
rect 20763 8316 20996 8344
rect 20763 8313 20775 8316
rect 20717 8307 20775 8313
rect 20990 8304 20996 8316
rect 21048 8304 21054 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 3973 7939 4031 7945
rect 3973 7905 3985 7939
rect 4019 7936 4031 7939
rect 8294 7936 8300 7948
rect 4019 7908 8300 7936
rect 4019 7905 4031 7908
rect 3973 7899 4031 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 23290 7896 23296 7948
rect 23348 7896 23354 7948
rect 6270 7868 6276 7880
rect 5382 7840 6276 7868
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 21450 7828 21456 7880
rect 21508 7868 21514 7880
rect 21545 7871 21603 7877
rect 21545 7868 21557 7871
rect 21508 7840 21557 7868
rect 21508 7828 21514 7840
rect 21545 7837 21557 7840
rect 21591 7837 21603 7871
rect 21545 7831 21603 7837
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 22649 7871 22707 7877
rect 22649 7868 22661 7871
rect 21692 7840 22661 7868
rect 21692 7828 21698 7840
rect 22649 7837 22661 7840
rect 22695 7837 22707 7871
rect 22649 7831 22707 7837
rect 24854 7828 24860 7880
rect 24912 7828 24918 7880
rect 4246 7760 4252 7812
rect 4304 7760 4310 7812
rect 5997 7803 6055 7809
rect 5997 7769 6009 7803
rect 6043 7800 6055 7803
rect 8570 7800 8576 7812
rect 6043 7772 8576 7800
rect 6043 7769 6055 7772
rect 5997 7763 6055 7769
rect 8570 7760 8576 7772
rect 8628 7760 8634 7812
rect 15930 7760 15936 7812
rect 15988 7800 15994 7812
rect 19521 7803 19579 7809
rect 19521 7800 19533 7803
rect 15988 7772 19533 7800
rect 15988 7760 15994 7772
rect 19521 7769 19533 7772
rect 19567 7769 19579 7803
rect 19521 7763 19579 7769
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 22002 7800 22008 7812
rect 19751 7772 22008 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 21726 7692 21732 7744
rect 21784 7692 21790 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24673 7735 24731 7741
rect 24673 7732 24685 7735
rect 24176 7704 24685 7732
rect 24176 7692 24182 7704
rect 24673 7701 24685 7704
rect 24719 7701 24731 7735
rect 24673 7695 24731 7701
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4304 7500 4629 7528
rect 4304 7488 4310 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 4617 7491 4675 7497
rect 15470 7420 15476 7472
rect 15528 7460 15534 7472
rect 18417 7463 18475 7469
rect 18417 7460 18429 7463
rect 15528 7432 18429 7460
rect 15528 7420 15534 7432
rect 18417 7429 18429 7432
rect 18463 7429 18475 7463
rect 18417 7423 18475 7429
rect 23382 7420 23388 7472
rect 23440 7420 23446 7472
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 20622 7352 20628 7404
rect 20680 7352 20686 7404
rect 23293 7395 23351 7401
rect 23293 7361 23305 7395
rect 23339 7392 23351 7395
rect 23400 7392 23428 7420
rect 23339 7364 23428 7392
rect 23937 7395 23995 7401
rect 23339 7361 23351 7364
rect 23293 7355 23351 7361
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 23017 7327 23075 7333
rect 23017 7293 23029 7327
rect 23063 7324 23075 7327
rect 23382 7324 23388 7336
rect 23063 7296 23388 7324
rect 23063 7293 23075 7296
rect 23017 7287 23075 7293
rect 23382 7284 23388 7296
rect 23440 7284 23446 7336
rect 16298 7216 16304 7268
rect 16356 7256 16362 7268
rect 23952 7256 23980 7355
rect 16356 7228 23980 7256
rect 16356 7216 16362 7228
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 20254 7188 20260 7200
rect 18555 7160 20260 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 20346 7148 20352 7200
rect 20404 7188 20410 7200
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 20404 7160 20453 7188
rect 20404 7148 20410 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 20441 7151 20499 7157
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 23385 6851 23443 6857
rect 23385 6817 23397 6851
rect 23431 6848 23443 6851
rect 24854 6848 24860 6860
rect 23431 6820 24860 6848
rect 23431 6817 23443 6820
rect 23385 6811 23443 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 17276 6752 19625 6780
rect 17276 6740 17282 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 6178 6644 6184 6656
rect 3200 6616 6184 6644
rect 3200 6604 3206 6616
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 19797 6647 19855 6653
rect 19797 6613 19809 6647
rect 19843 6644 19855 6647
rect 20824 6644 20852 6743
rect 24026 6740 24032 6792
rect 24084 6740 24090 6792
rect 24578 6740 24584 6792
rect 24636 6780 24642 6792
rect 24765 6783 24823 6789
rect 24765 6780 24777 6783
rect 24636 6752 24777 6780
rect 24636 6740 24642 6752
rect 24765 6749 24777 6752
rect 24811 6749 24823 6783
rect 24765 6743 24823 6749
rect 21910 6672 21916 6724
rect 21968 6672 21974 6724
rect 19843 6616 20852 6644
rect 19843 6613 19855 6616
rect 19797 6607 19855 6613
rect 21450 6604 21456 6656
rect 21508 6644 21514 6656
rect 24581 6647 24639 6653
rect 24581 6644 24593 6647
rect 21508 6616 24593 6644
rect 21508 6604 21514 6616
rect 24581 6613 24593 6616
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 3697 6443 3755 6449
rect 3697 6409 3709 6443
rect 3743 6440 3755 6443
rect 3970 6440 3976 6452
rect 3743 6412 3976 6440
rect 3743 6409 3755 6412
rect 3697 6403 3755 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 19521 6443 19579 6449
rect 19521 6409 19533 6443
rect 19567 6440 19579 6443
rect 21634 6440 21640 6452
rect 19567 6412 21640 6440
rect 19567 6409 19579 6412
rect 19521 6403 19579 6409
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 19429 6375 19487 6381
rect 19429 6341 19441 6375
rect 19475 6372 19487 6375
rect 19702 6372 19708 6384
rect 19475 6344 19708 6372
rect 19475 6341 19487 6344
rect 19429 6335 19487 6341
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2832 6276 3065 6304
rect 2832 6264 2838 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 21450 6264 21456 6316
rect 21508 6264 21514 6316
rect 22002 6264 22008 6316
rect 22060 6304 22066 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 22060 6276 22109 6304
rect 22060 6264 22066 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 23934 6264 23940 6316
rect 23992 6264 23998 6316
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6205 21051 6239
rect 20993 6199 21051 6205
rect 21008 6168 21036 6199
rect 22278 6196 22284 6248
rect 22336 6236 22342 6248
rect 22557 6239 22615 6245
rect 22557 6236 22569 6239
rect 22336 6208 22569 6236
rect 22336 6196 22342 6208
rect 22557 6205 22569 6208
rect 22603 6205 22615 6239
rect 22557 6199 22615 6205
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 22830 6168 22836 6180
rect 21008 6140 22836 6168
rect 22830 6128 22836 6140
rect 22888 6128 22894 6180
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 21910 5720 21916 5772
rect 21968 5760 21974 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 21968 5732 22477 5760
rect 21968 5720 21974 5732
rect 22465 5729 22477 5732
rect 22511 5729 22523 5763
rect 22465 5723 22523 5729
rect 20346 5652 20352 5704
rect 20404 5652 20410 5704
rect 21542 5652 21548 5704
rect 21600 5692 21606 5704
rect 22005 5695 22063 5701
rect 22005 5692 22017 5695
rect 21600 5664 22017 5692
rect 21600 5652 21606 5664
rect 22005 5661 22017 5664
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 22186 5652 22192 5704
rect 22244 5692 22250 5704
rect 24765 5695 24823 5701
rect 24765 5692 24777 5695
rect 22244 5664 24777 5692
rect 22244 5652 22250 5664
rect 24765 5661 24777 5664
rect 24811 5661 24823 5695
rect 24765 5655 24823 5661
rect 21358 5584 21364 5636
rect 21416 5584 21422 5636
rect 23014 5584 23020 5636
rect 23072 5624 23078 5636
rect 24581 5627 24639 5633
rect 24581 5624 24593 5627
rect 23072 5596 24593 5624
rect 23072 5584 23078 5596
rect 24581 5593 24593 5596
rect 24627 5593 24639 5627
rect 24581 5587 24639 5593
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 21450 5556 21456 5568
rect 20036 5528 21456 5556
rect 20036 5516 20042 5528
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 2774 5352 2780 5364
rect 2547 5324 2780 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 23014 5284 23020 5296
rect 19260 5256 23020 5284
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1728 5188 1777 5216
rect 1728 5176 1734 5188
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3970 5216 3976 5228
rect 3191 5188 3976 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 19260 5225 19288 5256
rect 23014 5244 23020 5256
rect 23072 5244 23078 5296
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5185 19303 5219
rect 19245 5179 19303 5185
rect 20990 5176 20996 5228
rect 21048 5176 21054 5228
rect 21818 5176 21824 5228
rect 21876 5216 21882 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21876 5188 22017 5216
rect 21876 5176 21882 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 24118 5176 24124 5228
rect 24176 5176 24182 5228
rect 18877 5151 18935 5157
rect 18877 5117 18889 5151
rect 18923 5117 18935 5151
rect 18877 5111 18935 5117
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 5534 5080 5540 5092
rect 1995 5052 5540 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 5534 5040 5540 5052
rect 5592 5040 5598 5092
rect 18892 5080 18920 5111
rect 19702 5108 19708 5160
rect 19760 5148 19766 5160
rect 19981 5151 20039 5157
rect 19981 5148 19993 5151
rect 19760 5120 19993 5148
rect 19760 5108 19766 5120
rect 19981 5117 19993 5120
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 22462 5108 22468 5160
rect 22520 5108 22526 5160
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 21818 5080 21824 5092
rect 18892 5052 21824 5080
rect 21818 5040 21824 5052
rect 21876 5040 21882 5092
rect 1489 5015 1547 5021
rect 1489 4981 1501 5015
rect 1535 5012 1547 5015
rect 1670 5012 1676 5024
rect 1535 4984 1676 5012
rect 1535 4981 1547 4984
rect 1489 4975 1547 4981
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 13354 5012 13360 5024
rect 9548 4984 13360 5012
rect 9548 4972 9554 4984
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 3970 4768 3976 4820
rect 4028 4768 4034 4820
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 9122 4740 9128 4752
rect 2915 4712 9128 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 9122 4700 9128 4712
rect 9180 4700 9186 4752
rect 22094 4740 22100 4752
rect 18432 4712 22100 4740
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 8294 4672 8300 4684
rect 1995 4644 8300 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 13446 4632 13452 4684
rect 13504 4672 13510 4684
rect 13630 4672 13636 4684
rect 13504 4644 13636 4672
rect 13504 4632 13510 4644
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 18432 4681 18460 4712
rect 22094 4700 22100 4712
rect 22152 4700 22158 4752
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4641 18475 4675
rect 23477 4675 23535 4681
rect 23477 4672 23489 4675
rect 18417 4635 18475 4641
rect 18892 4644 23489 4672
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2685 4607 2743 4613
rect 2685 4604 2697 4607
rect 2556 4576 2697 4604
rect 2556 4564 2562 4576
rect 2685 4573 2697 4576
rect 2731 4604 2743 4607
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 2731 4576 3249 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 18892 4613 18920 4644
rect 23477 4641 23489 4644
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 19610 4564 19616 4616
rect 19668 4564 19674 4616
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 21726 4564 21732 4616
rect 21784 4604 21790 4616
rect 23201 4607 23259 4613
rect 23201 4604 23213 4607
rect 21784 4576 23213 4604
rect 21784 4564 21790 4576
rect 23201 4573 23213 4576
rect 23247 4573 23259 4607
rect 23201 4567 23259 4573
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4505 1823 4539
rect 1765 4499 1823 4505
rect 1780 4468 1808 4499
rect 20346 4496 20352 4548
rect 20404 4496 20410 4548
rect 22189 4539 22247 4545
rect 22189 4505 22201 4539
rect 22235 4505 22247 4539
rect 22189 4499 22247 4505
rect 2038 4468 2044 4480
rect 1780 4440 2044 4468
rect 2038 4428 2044 4440
rect 2096 4468 2102 4480
rect 2225 4471 2283 4477
rect 2225 4468 2237 4471
rect 2096 4440 2237 4468
rect 2096 4428 2102 4440
rect 2225 4437 2237 4440
rect 2271 4437 2283 4471
rect 2225 4431 2283 4437
rect 20070 4428 20076 4480
rect 20128 4468 20134 4480
rect 22204 4468 22232 4499
rect 20128 4440 22232 4468
rect 20128 4428 20134 4440
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 22112 4168 22324 4196
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1452 4100 1593 4128
rect 1452 4088 1458 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 7558 4128 7564 4140
rect 3375 4100 7564 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 11974 4088 11980 4140
rect 12032 4088 12038 4140
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16408 4100 16865 4128
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 3476 4032 3617 4060
rect 3476 4020 3482 4032
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 3620 3992 3648 4023
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 4065 4063 4123 4069
rect 4065 4060 4077 4063
rect 3936 4032 4077 4060
rect 3936 4020 3942 4032
rect 4065 4029 4077 4032
rect 4111 4029 4123 4063
rect 4065 4023 4123 4029
rect 7466 4020 7472 4072
rect 7524 4060 7530 4072
rect 10410 4060 10416 4072
rect 7524 4032 10416 4060
rect 7524 4020 7530 4032
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11606 4060 11612 4072
rect 11379 4032 11612 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11606 4020 11612 4032
rect 11664 4060 11670 4072
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11664 4032 11713 4060
rect 11664 4020 11670 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13504 4032 14013 4060
rect 13504 4020 13510 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 15838 4020 15844 4072
rect 15896 4060 15902 4072
rect 16408 4060 16436 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 18782 4088 18788 4140
rect 18840 4088 18846 4140
rect 20254 4088 20260 4140
rect 20312 4128 20318 4140
rect 22112 4128 22140 4168
rect 20312 4100 22140 4128
rect 20312 4088 20318 4100
rect 22186 4088 22192 4140
rect 22244 4088 22250 4140
rect 22296 4128 22324 4168
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 22296 4100 23857 4128
rect 23845 4097 23857 4100
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 15896 4032 16436 4060
rect 16546 4032 17325 4060
rect 15896 4020 15902 4032
rect 3973 3995 4031 4001
rect 3973 3992 3985 3995
rect 3620 3964 3985 3992
rect 3973 3961 3985 3964
rect 4019 3961 4031 3995
rect 4798 3992 4804 4004
rect 3973 3955 4031 3961
rect 4080 3964 4804 3992
rect 4080 3936 4108 3964
rect 4798 3952 4804 3964
rect 4856 3952 4862 4004
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 9953 3995 10011 4001
rect 9953 3992 9965 3995
rect 9640 3964 9965 3992
rect 9640 3952 9646 3964
rect 9953 3961 9965 3964
rect 9999 3961 10011 3995
rect 9953 3955 10011 3961
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 16546 3992 16574 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 17552 4032 19165 4060
rect 17552 4020 17558 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20438 4020 20444 4072
rect 20496 4060 20502 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 20496 4032 22477 4060
rect 20496 4020 20502 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 16448 3964 16574 3992
rect 16448 3952 16454 3964
rect 21542 3952 21548 4004
rect 21600 3992 21606 4004
rect 24320 3992 24348 4023
rect 21600 3964 24348 3992
rect 21600 3952 21606 3964
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 2682 3924 2688 3936
rect 2271 3896 2688 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 4062 3884 4068 3936
rect 4120 3884 4126 3936
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 4304 3896 4353 3924
rect 4304 3884 4310 3896
rect 4341 3893 4353 3896
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6144 3896 6377 3924
rect 6144 3884 6150 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 8754 3924 8760 3936
rect 6788 3896 8760 3924
rect 6788 3884 6794 3896
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9456 3896 9505 3924
rect 9456 3884 9462 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 9766 3884 9772 3936
rect 9824 3884 9830 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 11020 3896 11069 3924
rect 11020 3884 11026 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 8938 3720 8944 3732
rect 8251 3692 8944 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9214 3680 9220 3732
rect 9272 3680 9278 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 22646 3680 22652 3732
rect 22704 3720 22710 3732
rect 24946 3720 24952 3732
rect 22704 3692 24952 3720
rect 22704 3680 22710 3692
rect 24946 3680 24952 3692
rect 25004 3680 25010 3732
rect 4157 3655 4215 3661
rect 4157 3621 4169 3655
rect 4203 3621 4215 3655
rect 4157 3615 4215 3621
rect 4172 3584 4200 3615
rect 5258 3612 5264 3664
rect 5316 3612 5322 3664
rect 6089 3655 6147 3661
rect 6089 3621 6101 3655
rect 6135 3652 6147 3655
rect 16114 3652 16120 3664
rect 6135 3624 16120 3652
rect 6135 3621 6147 3624
rect 6089 3615 6147 3621
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 7466 3584 7472 3596
rect 4172 3556 7472 3584
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 8294 3584 8300 3596
rect 7607 3556 8300 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 14642 3584 14648 3596
rect 11287 3556 14648 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 14642 3544 14648 3556
rect 14700 3544 14706 3596
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 16080 3556 17325 3584
rect 16080 3544 16086 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17920 3556 19901 3584
rect 17920 3544 17926 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 2406 3476 2412 3528
rect 2464 3476 2470 3528
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 3145 3519 3203 3525
rect 3145 3516 3157 3519
rect 2915 3488 3157 3516
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 3145 3485 3157 3488
rect 3191 3516 3203 3519
rect 3510 3516 3516 3528
rect 3191 3488 3516 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 3973 3479 4031 3485
rect 5000 3488 5089 3516
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 3988 3448 4016 3479
rect 4525 3451 4583 3457
rect 4525 3448 4537 3451
rect 2832 3420 4537 3448
rect 2832 3408 2838 3420
rect 4525 3417 4537 3420
rect 4571 3417 4583 3451
rect 4525 3411 4583 3417
rect 5000 3392 5028 3488
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 6086 3516 6092 3528
rect 5951 3488 6092 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6512 3488 6561 3516
rect 6512 3476 6518 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 6549 3479 6607 3485
rect 7852 3488 8033 3516
rect 7852 3392 7880 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 9398 3476 9404 3528
rect 9456 3476 9462 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10870 3516 10876 3528
rect 10551 3488 10876 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10928 3488 10977 3516
rect 10928 3476 10934 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14182 3516 14188 3528
rect 13771 3488 14188 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3516 16451 3519
rect 16574 3516 16580 3528
rect 16439 3488 16580 3516
rect 16439 3485 16451 3488
rect 16393 3479 16451 3485
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16850 3476 16856 3528
rect 16908 3476 16914 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18380 3488 19441 3516
rect 18380 3476 18386 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20864 3488 21281 3516
rect 20864 3476 20870 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 12710 3408 12716 3460
rect 12768 3408 12774 3460
rect 14918 3408 14924 3460
rect 14976 3448 14982 3460
rect 15197 3451 15255 3457
rect 15197 3448 15209 3451
rect 14976 3420 15209 3448
rect 14976 3408 14982 3420
rect 15197 3417 15209 3420
rect 15243 3417 15255 3451
rect 15197 3411 15255 3417
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 21744 3448 21772 3547
rect 19024 3420 21772 3448
rect 19024 3408 19030 3420
rect 1394 3340 1400 3392
rect 1452 3340 1458 3392
rect 1762 3340 1768 3392
rect 1820 3340 1826 3392
rect 3326 3340 3332 3392
rect 3384 3340 3390 3392
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 4982 3380 4988 3392
rect 4847 3352 4988 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 6880 3352 7205 3380
rect 6880 3340 6886 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7193 3343 7251 3349
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 7834 3380 7840 3392
rect 7791 3352 7840 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8662 3340 8668 3392
rect 8720 3340 8726 3392
rect 10689 3383 10747 3389
rect 10689 3349 10701 3383
rect 10735 3380 10747 3383
rect 11238 3380 11244 3392
rect 10735 3352 11244 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 23382 3380 23388 3392
rect 22060 3352 23388 3380
rect 22060 3340 22066 3352
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 3513 3179 3571 3185
rect 3513 3176 3525 3179
rect 2464 3148 3525 3176
rect 2464 3136 2470 3148
rect 3513 3145 3525 3148
rect 3559 3145 3571 3179
rect 3513 3139 3571 3145
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 5902 3136 5908 3188
rect 5960 3136 5966 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7432 3148 7757 3176
rect 7432 3136 7438 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8386 3136 8392 3188
rect 8444 3136 8450 3188
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11112 3148 11897 3176
rect 11112 3136 11118 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19392 3148 22968 3176
rect 19392 3136 19398 3148
rect 4249 3111 4307 3117
rect 4249 3077 4261 3111
rect 4295 3108 4307 3111
rect 7190 3108 7196 3120
rect 4295 3080 7196 3108
rect 4295 3077 4307 3080
rect 4249 3071 4307 3077
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 9582 3068 9588 3120
rect 9640 3068 9646 3120
rect 14826 3108 14832 3120
rect 13740 3080 14832 3108
rect 1762 3000 1768 3052
rect 1820 3000 1826 3052
rect 2866 3000 2872 3052
rect 2924 3000 2930 3052
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 3936 3012 4077 3040
rect 3936 3000 3942 3012
rect 4065 3009 4077 3012
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4755 3012 4997 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5350 3040 5356 3052
rect 5031 3012 5356 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8294 3040 8300 3052
rect 7607 3012 8300 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8662 3040 8668 3052
rect 8619 3012 8668 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9600 3040 9628 3068
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9088 3012 9873 3040
rect 9088 3000 9094 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 10962 3040 10968 3052
rect 10560 3012 10968 3040
rect 10560 3000 10566 3012
rect 10962 3000 10968 3012
rect 11020 3040 11026 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 11020 3012 11161 3040
rect 11020 3000 11026 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 13740 3049 13768 3080
rect 14826 3068 14832 3080
rect 14884 3068 14890 3120
rect 18598 3068 18604 3120
rect 18656 3108 18662 3120
rect 20346 3108 20352 3120
rect 18656 3080 20352 3108
rect 18656 3068 18662 3080
rect 20346 3068 20352 3080
rect 20404 3068 20410 3120
rect 21450 3068 21456 3120
rect 21508 3108 21514 3120
rect 22940 3117 22968 3148
rect 21545 3111 21603 3117
rect 21545 3108 21557 3111
rect 21508 3080 21557 3108
rect 21508 3068 21514 3080
rect 21545 3077 21557 3080
rect 21591 3108 21603 3111
rect 22925 3111 22983 3117
rect 21591 3080 22048 3108
rect 21591 3077 21603 3080
rect 21545 3071 21603 3077
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11296 3012 11713 3040
rect 11296 3000 11302 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16540 3012 16865 3040
rect 16540 3000 16546 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 18506 3040 18512 3052
rect 17736 3012 18512 3040
rect 17736 3000 17742 3012
rect 18506 3000 18512 3012
rect 18564 3040 18570 3052
rect 18693 3043 18751 3049
rect 18693 3040 18705 3043
rect 18564 3012 18705 3040
rect 18564 3000 18570 3012
rect 18693 3009 18705 3012
rect 18739 3009 18751 3043
rect 20714 3040 20720 3052
rect 18693 3003 18751 3009
rect 18800 3012 20720 3040
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 4154 2972 4160 2984
rect 2455 2944 4160 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 9490 2932 9496 2984
rect 9548 2972 9554 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 9548 2944 9597 2972
rect 9548 2932 9554 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2941 10931 2975
rect 10873 2935 10931 2941
rect 10888 2904 10916 2935
rect 13354 2932 13360 2984
rect 13412 2932 13418 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14240 2944 14749 2972
rect 14240 2932 14246 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15712 2944 17325 2972
rect 15712 2932 15718 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 18322 2932 18328 2984
rect 18380 2972 18386 2984
rect 18800 2972 18828 3012
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 22020 3049 22048 3080
rect 22925 3077 22937 3111
rect 22971 3077 22983 3111
rect 22925 3071 22983 3077
rect 22005 3043 22063 3049
rect 22005 3009 22017 3043
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 22612 3012 23857 3040
rect 22612 3000 22618 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 18380 2944 18828 2972
rect 19153 2975 19211 2981
rect 18380 2932 18386 2944
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 13906 2904 13912 2916
rect 10888 2876 13912 2904
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 19168 2904 19196 2935
rect 21174 2932 21180 2984
rect 21232 2972 21238 2984
rect 22462 2972 22468 2984
rect 21232 2944 22468 2972
rect 21232 2932 21238 2944
rect 22462 2932 22468 2944
rect 22520 2932 22526 2984
rect 24305 2975 24363 2981
rect 24305 2941 24317 2975
rect 24351 2941 24363 2975
rect 24305 2935 24363 2941
rect 17184 2876 19196 2904
rect 17184 2864 17190 2876
rect 21358 2864 21364 2916
rect 21416 2904 21422 2916
rect 22646 2904 22652 2916
rect 21416 2876 22652 2904
rect 21416 2864 21422 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 6454 2796 6460 2848
rect 6512 2796 6518 2848
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 11330 2836 11336 2848
rect 7055 2808 11336 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 19886 2836 19892 2848
rect 16816 2808 19892 2836
rect 16816 2796 16822 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 24320 2836 24348 2935
rect 20864 2808 24348 2836
rect 20864 2796 20870 2808
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2866 2632 2872 2644
rect 1627 2604 2872 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4062 2592 4068 2644
rect 4120 2592 4126 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 14458 2632 14464 2644
rect 9815 2604 14464 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 18506 2592 18512 2644
rect 18564 2592 18570 2644
rect 24670 2592 24676 2644
rect 24728 2592 24734 2644
rect 13630 2564 13636 2576
rect 10888 2536 13636 2564
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 2240 2468 3341 2496
rect 2240 2437 2268 2468
rect 3329 2465 3341 2468
rect 3375 2465 3387 2499
rect 3329 2459 3387 2465
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 10594 2496 10600 2508
rect 5307 2468 10600 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 10888 2505 10916 2536
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 10873 2499 10931 2505
rect 10873 2465 10885 2499
rect 10919 2465 10931 2499
rect 11974 2496 11980 2508
rect 10873 2459 10931 2465
rect 11716 2468 11980 2496
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2682 2388 2688 2440
rect 2740 2388 2746 2440
rect 4246 2388 4252 2440
rect 4304 2388 4310 2440
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 4672 2400 5549 2428
rect 4672 2388 4678 2400
rect 5537 2397 5549 2400
rect 5583 2428 5595 2431
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 5583 2400 5825 2428
rect 5583 2397 5595 2400
rect 5537 2391 5595 2397
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6503 2400 6929 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6917 2397 6929 2400
rect 6963 2428 6975 2431
rect 7190 2428 7196 2440
rect 6963 2400 7196 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8938 2428 8944 2440
rect 7975 2400 8944 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9171 2400 9597 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9585 2397 9597 2400
rect 9631 2428 9643 2431
rect 10134 2428 10140 2440
rect 9631 2400 10140 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11716 2437 11744 2468
rect 11974 2456 11980 2468
rect 12032 2496 12038 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 12032 2468 14105 2496
rect 12032 2456 12038 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14608 2468 15209 2496
rect 14608 2456 14614 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15344 2468 17325 2496
rect 15344 2456 15350 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17770 2456 17776 2508
rect 17828 2496 17834 2508
rect 17828 2468 19564 2496
rect 17828 2456 17834 2468
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12124 2400 12357 2428
rect 12124 2388 12130 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 14645 2431 14703 2437
rect 14645 2428 14657 2431
rect 12860 2400 14657 2428
rect 12860 2388 12866 2400
rect 14645 2397 14657 2400
rect 14691 2397 14703 2431
rect 14645 2391 14703 2397
rect 17034 2388 17040 2440
rect 17092 2388 17098 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19536 2428 19564 2468
rect 19886 2456 19892 2508
rect 19944 2456 19950 2508
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 20772 2468 22477 2496
rect 20772 2456 20778 2468
rect 22465 2465 22477 2468
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 19536 2400 22017 2428
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 24029 2431 24087 2437
rect 24029 2397 24041 2431
rect 24075 2428 24087 2431
rect 25038 2428 25044 2440
rect 24075 2400 25044 2428
rect 24075 2397 24087 2400
rect 24029 2391 24087 2397
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 5718 2320 5724 2372
rect 5776 2360 5782 2372
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 5776 2332 6101 2360
rect 5776 2320 5782 2332
rect 6089 2329 6101 2332
rect 6135 2329 6147 2363
rect 6089 2323 6147 2329
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 7576 2360 7604 2388
rect 6687 2332 7604 2360
rect 9309 2363 9367 2369
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 11164 2360 11192 2388
rect 9355 2332 11192 2360
rect 13541 2363 13599 2369
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 13814 2360 13820 2372
rect 13587 2332 13820 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 24118 2320 24124 2372
rect 24176 2360 24182 2372
rect 24765 2363 24823 2369
rect 24765 2360 24777 2363
rect 24176 2332 24777 2360
rect 24176 2320 24182 2332
rect 24765 2329 24777 2332
rect 24811 2360 24823 2363
rect 25133 2363 25191 2369
rect 25133 2360 25145 2363
rect 24811 2332 25145 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 25133 2329 25145 2332
rect 25179 2329 25191 2363
rect 25133 2323 25191 2329
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2292 11943 2295
rect 12250 2292 12256 2304
rect 11931 2264 12256 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 8938 2048 8944 2100
rect 8996 2088 9002 2100
rect 13906 2088 13912 2100
rect 8996 2060 13912 2088
rect 8996 2048 9002 2060
rect 13906 2048 13912 2060
rect 13964 2048 13970 2100
rect 12250 1980 12256 2032
rect 12308 2020 12314 2032
rect 17310 2020 17316 2032
rect 12308 1992 17316 2020
rect 12308 1980 12314 1992
rect 17310 1980 17316 1992
rect 17368 1980 17374 2032
rect 7098 1912 7104 1964
rect 7156 1952 7162 1964
rect 13722 1952 13728 1964
rect 7156 1924 13728 1952
rect 7156 1912 7162 1924
rect 13722 1912 13728 1924
rect 13780 1912 13786 1964
rect 11146 1844 11152 1896
rect 11204 1884 11210 1896
rect 12342 1884 12348 1896
rect 11204 1856 12348 1884
rect 11204 1844 11210 1856
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 14740 54272 14792 54324
rect 16212 54272 16264 54324
rect 5632 54136 5684 54188
rect 6000 54179 6052 54188
rect 6000 54145 6009 54179
rect 6009 54145 6043 54179
rect 6043 54145 6052 54179
rect 6000 54136 6052 54145
rect 3976 54068 4028 54120
rect 7840 54136 7892 54188
rect 9956 54179 10008 54188
rect 9956 54145 9965 54179
rect 9965 54145 9999 54179
rect 9999 54145 10008 54179
rect 9956 54136 10008 54145
rect 11428 54204 11480 54256
rect 11520 54136 11572 54188
rect 12900 54204 12952 54256
rect 12532 54179 12584 54188
rect 12532 54145 12541 54179
rect 12541 54145 12575 54179
rect 12575 54145 12584 54179
rect 12532 54136 12584 54145
rect 15200 54136 15252 54188
rect 24492 54315 24544 54324
rect 24492 54281 24501 54315
rect 24501 54281 24535 54315
rect 24535 54281 24544 54315
rect 24492 54272 24544 54281
rect 24676 54315 24728 54324
rect 24676 54281 24685 54315
rect 24685 54281 24719 54315
rect 24719 54281 24728 54315
rect 24676 54272 24728 54281
rect 16948 54136 17000 54188
rect 19524 54204 19576 54256
rect 17960 54136 18012 54188
rect 18512 54179 18564 54188
rect 18512 54145 18521 54179
rect 18521 54145 18555 54179
rect 18555 54145 18564 54179
rect 18512 54136 18564 54145
rect 18604 54136 18656 54188
rect 19708 54179 19760 54188
rect 19708 54145 19717 54179
rect 19717 54145 19751 54179
rect 19751 54145 19760 54179
rect 19708 54136 19760 54145
rect 20720 54136 20772 54188
rect 21180 54179 21232 54188
rect 21180 54145 21189 54179
rect 21189 54145 21223 54179
rect 21223 54145 21232 54179
rect 21180 54136 21232 54145
rect 21364 54136 21416 54188
rect 22468 54136 22520 54188
rect 25320 54179 25372 54188
rect 25320 54145 25329 54179
rect 25329 54145 25363 54179
rect 25363 54145 25372 54179
rect 25320 54136 25372 54145
rect 9864 54068 9916 54120
rect 12624 54068 12676 54120
rect 16764 54000 16816 54052
rect 12716 53932 12768 53984
rect 15016 53975 15068 53984
rect 15016 53941 15025 53975
rect 15025 53941 15059 53975
rect 15059 53941 15068 53975
rect 15016 53932 15068 53941
rect 15752 53932 15804 53984
rect 17040 53975 17092 53984
rect 17040 53941 17049 53975
rect 17049 53941 17083 53975
rect 17083 53941 17092 53975
rect 17040 53932 17092 53941
rect 18420 53975 18472 53984
rect 18420 53941 18429 53975
rect 18429 53941 18463 53975
rect 18463 53941 18472 53975
rect 18420 53932 18472 53941
rect 19340 53932 19392 53984
rect 20444 53932 20496 53984
rect 21640 53932 21692 53984
rect 22192 53932 22244 53984
rect 22284 53932 22336 53984
rect 24584 53932 24636 53984
rect 25964 53932 26016 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 3976 53728 4028 53780
rect 5908 53728 5960 53780
rect 16580 53728 16632 53780
rect 18512 53728 18564 53780
rect 2412 53388 2464 53440
rect 20628 53660 20680 53712
rect 22284 53660 22336 53712
rect 5540 53524 5592 53576
rect 8852 53592 8904 53644
rect 11060 53635 11112 53644
rect 11060 53601 11069 53635
rect 11069 53601 11103 53635
rect 11103 53601 11112 53635
rect 11060 53592 11112 53601
rect 12164 53592 12216 53644
rect 6736 53567 6788 53576
rect 6736 53533 6745 53567
rect 6745 53533 6779 53567
rect 6779 53533 6788 53567
rect 6736 53524 6788 53533
rect 8576 53567 8628 53576
rect 8576 53533 8585 53567
rect 8585 53533 8619 53567
rect 8619 53533 8628 53567
rect 8576 53524 8628 53533
rect 9128 53567 9180 53576
rect 9128 53533 9137 53567
rect 9137 53533 9171 53567
rect 9171 53533 9180 53567
rect 9128 53524 9180 53533
rect 12072 53524 12124 53576
rect 12624 53524 12676 53576
rect 14004 53524 14056 53576
rect 15476 53524 15528 53576
rect 16580 53524 16632 53576
rect 17316 53524 17368 53576
rect 18328 53567 18380 53576
rect 18328 53533 18337 53567
rect 18337 53533 18371 53567
rect 18371 53533 18380 53567
rect 18328 53524 18380 53533
rect 19156 53524 19208 53576
rect 19892 53524 19944 53576
rect 20996 53524 21048 53576
rect 21732 53524 21784 53576
rect 22100 53524 22152 53576
rect 22836 53524 22888 53576
rect 24492 53524 24544 53576
rect 24768 53524 24820 53576
rect 7380 53456 7432 53508
rect 7288 53388 7340 53440
rect 14648 53388 14700 53440
rect 15844 53388 15896 53440
rect 17040 53388 17092 53440
rect 17592 53431 17644 53440
rect 17592 53397 17601 53431
rect 17601 53397 17635 53431
rect 17635 53397 17644 53431
rect 17592 53388 17644 53397
rect 18328 53388 18380 53440
rect 19616 53431 19668 53440
rect 19616 53397 19625 53431
rect 19625 53397 19659 53431
rect 19659 53397 19668 53431
rect 19616 53388 19668 53397
rect 20536 53388 20588 53440
rect 21272 53431 21324 53440
rect 21272 53397 21281 53431
rect 21281 53397 21315 53431
rect 21315 53397 21324 53431
rect 21272 53388 21324 53397
rect 21916 53388 21968 53440
rect 23848 53431 23900 53440
rect 23848 53397 23857 53431
rect 23857 53397 23891 53431
rect 23891 53397 23900 53431
rect 23848 53388 23900 53397
rect 25136 53431 25188 53440
rect 25136 53397 25145 53431
rect 25145 53397 25179 53431
rect 25179 53397 25188 53431
rect 25136 53388 25188 53397
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 17316 53227 17368 53236
rect 17316 53193 17325 53227
rect 17325 53193 17359 53227
rect 17359 53193 17368 53227
rect 17316 53184 17368 53193
rect 19156 53184 19208 53236
rect 19708 53227 19760 53236
rect 19708 53193 19717 53227
rect 19717 53193 19751 53227
rect 19751 53193 19760 53227
rect 19708 53184 19760 53193
rect 20996 53227 21048 53236
rect 20996 53193 21005 53227
rect 21005 53193 21039 53227
rect 21039 53193 21048 53227
rect 20996 53184 21048 53193
rect 21180 53227 21232 53236
rect 21180 53193 21189 53227
rect 21189 53193 21223 53227
rect 21223 53193 21232 53227
rect 21180 53184 21232 53193
rect 21732 53184 21784 53236
rect 22100 53184 22152 53236
rect 22468 53184 22520 53236
rect 23296 53184 23348 53236
rect 13636 53116 13688 53168
rect 2412 53048 2464 53100
rect 4252 53048 4304 53100
rect 6184 53048 6236 53100
rect 7196 53091 7248 53100
rect 7196 53057 7205 53091
rect 7205 53057 7239 53091
rect 7239 53057 7248 53091
rect 7196 53048 7248 53057
rect 8392 53048 8444 53100
rect 9496 53048 9548 53100
rect 11888 53091 11940 53100
rect 11888 53057 11897 53091
rect 11897 53057 11931 53091
rect 11931 53057 11940 53091
rect 11888 53048 11940 53057
rect 14372 53048 14424 53100
rect 15936 53091 15988 53100
rect 15936 53057 15945 53091
rect 15945 53057 15979 53091
rect 15979 53057 15988 53091
rect 15936 53048 15988 53057
rect 18788 53048 18840 53100
rect 20260 53048 20312 53100
rect 23572 53048 23624 53100
rect 25320 53091 25372 53100
rect 25320 53057 25329 53091
rect 25329 53057 25363 53091
rect 25363 53057 25372 53091
rect 25320 53048 25372 53057
rect 4436 52980 4488 53032
rect 6276 52980 6328 53032
rect 9220 52980 9272 53032
rect 10324 53023 10376 53032
rect 10324 52989 10333 53023
rect 10333 52989 10367 53023
rect 10367 52989 10376 53023
rect 10324 52980 10376 52989
rect 11796 52980 11848 53032
rect 2964 52912 3016 52964
rect 7840 52912 7892 52964
rect 14004 52955 14056 52964
rect 14004 52921 14013 52955
rect 14013 52921 14047 52955
rect 14047 52921 14056 52955
rect 14004 52912 14056 52921
rect 15568 52912 15620 52964
rect 1584 52844 1636 52896
rect 6552 52887 6604 52896
rect 6552 52853 6561 52887
rect 6561 52853 6595 52887
rect 6595 52853 6604 52887
rect 6552 52844 6604 52853
rect 16120 52887 16172 52896
rect 16120 52853 16129 52887
rect 16129 52853 16163 52887
rect 16163 52853 16172 52887
rect 16120 52844 16172 52853
rect 18880 52887 18932 52896
rect 18880 52853 18889 52887
rect 18889 52853 18923 52887
rect 18923 52853 18932 52887
rect 18880 52844 18932 52853
rect 20076 52844 20128 52896
rect 23296 52887 23348 52896
rect 23296 52853 23305 52887
rect 23305 52853 23339 52887
rect 23339 52853 23348 52887
rect 23296 52844 23348 52853
rect 23388 52844 23440 52896
rect 25688 52844 25740 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 3700 52640 3752 52692
rect 4252 52640 4304 52692
rect 12624 52683 12676 52692
rect 12624 52649 12633 52683
rect 12633 52649 12667 52683
rect 12667 52649 12676 52683
rect 12624 52640 12676 52649
rect 13636 52640 13688 52692
rect 24768 52640 24820 52692
rect 4988 52572 5040 52624
rect 25780 52572 25832 52624
rect 6644 52504 6696 52556
rect 7748 52547 7800 52556
rect 7748 52513 7757 52547
rect 7757 52513 7791 52547
rect 7791 52513 7800 52547
rect 7748 52504 7800 52513
rect 10692 52504 10744 52556
rect 3424 52436 3476 52488
rect 6828 52436 6880 52488
rect 8852 52436 8904 52488
rect 9588 52436 9640 52488
rect 12808 52479 12860 52488
rect 12808 52445 12817 52479
rect 12817 52445 12851 52479
rect 12851 52445 12860 52479
rect 12808 52436 12860 52445
rect 16304 52436 16356 52488
rect 25320 52479 25372 52488
rect 25320 52445 25329 52479
rect 25329 52445 25363 52479
rect 25363 52445 25372 52479
rect 25320 52436 25372 52445
rect 9312 52411 9364 52420
rect 9312 52377 9321 52411
rect 9321 52377 9355 52411
rect 9355 52377 9364 52411
rect 9312 52368 9364 52377
rect 13360 52368 13412 52420
rect 4620 52343 4672 52352
rect 4620 52309 4629 52343
rect 4629 52309 4663 52343
rect 4663 52309 4672 52343
rect 4620 52300 4672 52309
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 3332 52028 3384 52080
rect 6552 52096 6604 52148
rect 7196 52139 7248 52148
rect 7196 52105 7205 52139
rect 7205 52105 7239 52139
rect 7239 52105 7248 52139
rect 7196 52096 7248 52105
rect 11888 52139 11940 52148
rect 11888 52105 11897 52139
rect 11897 52105 11931 52139
rect 11931 52105 11940 52139
rect 11888 52096 11940 52105
rect 12532 52139 12584 52148
rect 12532 52105 12541 52139
rect 12541 52105 12575 52139
rect 12575 52105 12584 52139
rect 12532 52096 12584 52105
rect 13360 52096 13412 52148
rect 25228 52139 25280 52148
rect 25228 52105 25237 52139
rect 25237 52105 25271 52139
rect 25271 52105 25280 52139
rect 25228 52096 25280 52105
rect 3884 52028 3936 52080
rect 4804 52071 4856 52080
rect 4804 52037 4813 52071
rect 4813 52037 4847 52071
rect 4847 52037 4856 52071
rect 4804 52028 4856 52037
rect 6460 51960 6512 52012
rect 9680 52028 9732 52080
rect 8760 51960 8812 52012
rect 10876 52003 10928 52012
rect 10876 51969 10885 52003
rect 10885 51969 10919 52003
rect 10919 51969 10928 52003
rect 10876 51960 10928 51969
rect 11704 52003 11756 52012
rect 11704 51969 11713 52003
rect 11713 51969 11747 52003
rect 11747 51969 11756 52003
rect 11704 51960 11756 51969
rect 12348 52003 12400 52012
rect 12348 51969 12357 52003
rect 12357 51969 12391 52003
rect 12391 51969 12400 52003
rect 12348 51960 12400 51969
rect 4804 51892 4856 51944
rect 8484 51935 8536 51944
rect 8484 51901 8493 51935
rect 8493 51901 8527 51935
rect 8527 51901 8536 51935
rect 8484 51892 8536 51901
rect 9128 51824 9180 51876
rect 25320 51756 25372 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 9956 51552 10008 51604
rect 2872 51459 2924 51468
rect 2872 51425 2881 51459
rect 2881 51425 2915 51459
rect 2915 51425 2924 51459
rect 2872 51416 2924 51425
rect 5540 51459 5592 51468
rect 5540 51425 5549 51459
rect 5549 51425 5583 51459
rect 5583 51425 5592 51459
rect 5540 51416 5592 51425
rect 7012 51416 7064 51468
rect 4620 51391 4672 51400
rect 4620 51357 4629 51391
rect 4629 51357 4663 51391
rect 4663 51357 4672 51391
rect 4620 51348 4672 51357
rect 6644 51391 6696 51400
rect 6644 51357 6653 51391
rect 6653 51357 6687 51391
rect 6687 51357 6696 51391
rect 6644 51348 6696 51357
rect 8484 51391 8536 51400
rect 8484 51357 8493 51391
rect 8493 51357 8527 51391
rect 8527 51357 8536 51391
rect 8484 51348 8536 51357
rect 9036 51348 9088 51400
rect 25320 51391 25372 51400
rect 25320 51357 25329 51391
rect 25329 51357 25363 51391
rect 25363 51357 25372 51391
rect 25320 51348 25372 51357
rect 5540 51280 5592 51332
rect 3976 51255 4028 51264
rect 3976 51221 3985 51255
rect 3985 51221 4019 51255
rect 4019 51221 4028 51255
rect 3976 51212 4028 51221
rect 24860 51212 24912 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 3424 51008 3476 51060
rect 5540 51008 5592 51060
rect 2780 50983 2832 50992
rect 2780 50949 2789 50983
rect 2789 50949 2823 50983
rect 2823 50949 2832 50983
rect 2780 50940 2832 50949
rect 4160 50940 4212 50992
rect 6736 50940 6788 50992
rect 7840 50940 7892 50992
rect 9588 50983 9640 50992
rect 9588 50949 9597 50983
rect 9597 50949 9631 50983
rect 9631 50949 9640 50983
rect 9588 50940 9640 50949
rect 1584 50915 1636 50924
rect 1584 50881 1593 50915
rect 1593 50881 1627 50915
rect 1627 50881 1636 50915
rect 1584 50872 1636 50881
rect 3700 50915 3752 50924
rect 3700 50881 3709 50915
rect 3709 50881 3743 50915
rect 3743 50881 3752 50915
rect 3700 50872 3752 50881
rect 5448 50915 5500 50924
rect 5448 50881 5457 50915
rect 5457 50881 5491 50915
rect 5491 50881 5500 50915
rect 5448 50872 5500 50881
rect 6092 50872 6144 50924
rect 9220 50872 9272 50924
rect 25320 50915 25372 50924
rect 25320 50881 25329 50915
rect 25329 50881 25363 50915
rect 25363 50881 25372 50915
rect 25320 50872 25372 50881
rect 25504 50668 25556 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 8576 50464 8628 50516
rect 2228 50371 2280 50380
rect 2228 50337 2237 50371
rect 2237 50337 2271 50371
rect 2271 50337 2280 50371
rect 2228 50328 2280 50337
rect 5632 50328 5684 50380
rect 25412 50328 25464 50380
rect 3884 50260 3936 50312
rect 3976 50303 4028 50312
rect 3976 50269 3985 50303
rect 3985 50269 4019 50303
rect 4019 50269 4028 50303
rect 3976 50260 4028 50269
rect 7472 50303 7524 50312
rect 7472 50269 7481 50303
rect 7481 50269 7515 50303
rect 7515 50269 7524 50303
rect 7472 50260 7524 50269
rect 9404 50303 9456 50312
rect 9404 50269 9413 50303
rect 9413 50269 9447 50303
rect 9447 50269 9456 50303
rect 9404 50260 9456 50269
rect 25320 50303 25372 50312
rect 25320 50269 25329 50303
rect 25329 50269 25363 50303
rect 25363 50269 25372 50303
rect 25320 50260 25372 50269
rect 4252 50124 4304 50176
rect 21548 50124 21600 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 1860 49852 1912 49904
rect 3424 49784 3476 49836
rect 10048 49920 10100 49972
rect 12348 49920 12400 49972
rect 4252 49895 4304 49904
rect 4252 49861 4261 49895
rect 4261 49861 4295 49895
rect 4295 49861 4304 49895
rect 4252 49852 4304 49861
rect 7748 49784 7800 49836
rect 9496 49895 9548 49904
rect 9496 49861 9505 49895
rect 9505 49861 9539 49895
rect 9539 49861 9548 49895
rect 9496 49852 9548 49861
rect 11060 49784 11112 49836
rect 11428 49784 11480 49836
rect 8576 49716 8628 49768
rect 19800 49716 19852 49768
rect 25412 49716 25464 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 12808 49419 12860 49428
rect 12808 49385 12817 49419
rect 12817 49385 12851 49419
rect 12851 49385 12860 49419
rect 12808 49376 12860 49385
rect 1492 49240 1544 49292
rect 13544 49172 13596 49224
rect 25320 49215 25372 49224
rect 25320 49181 25329 49215
rect 25329 49181 25363 49215
rect 25363 49181 25372 49215
rect 25320 49172 25372 49181
rect 3516 49036 3568 49088
rect 18972 49036 19024 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 25872 48696 25924 48748
rect 25228 48628 25280 48680
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 18328 48263 18380 48272
rect 17316 48195 17368 48204
rect 17316 48161 17325 48195
rect 17325 48161 17359 48195
rect 17359 48161 17368 48195
rect 17316 48152 17368 48161
rect 18328 48229 18337 48263
rect 18337 48229 18371 48263
rect 18371 48229 18380 48263
rect 18328 48220 18380 48229
rect 18696 48220 18748 48272
rect 17592 48127 17644 48136
rect 17592 48093 17601 48127
rect 17601 48093 17635 48127
rect 17635 48093 17644 48127
rect 17592 48084 17644 48093
rect 18788 48084 18840 48136
rect 17684 47948 17736 48000
rect 19524 47948 19576 48000
rect 25228 47991 25280 48000
rect 25228 47957 25237 47991
rect 25237 47957 25271 47991
rect 25271 47957 25280 47991
rect 25228 47948 25280 47957
rect 25320 47948 25372 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9312 47744 9364 47796
rect 11704 47744 11756 47796
rect 16120 47744 16172 47796
rect 18236 47744 18288 47796
rect 19064 47676 19116 47728
rect 19524 47719 19576 47728
rect 19524 47685 19533 47719
rect 19533 47685 19567 47719
rect 19567 47685 19576 47719
rect 19524 47676 19576 47685
rect 10968 47608 11020 47660
rect 11704 47651 11756 47660
rect 11704 47617 11713 47651
rect 11713 47617 11747 47651
rect 11747 47617 11756 47651
rect 11704 47608 11756 47617
rect 20168 47608 20220 47660
rect 17408 47583 17460 47592
rect 17408 47549 17417 47583
rect 17417 47549 17451 47583
rect 17451 47549 17460 47583
rect 17408 47540 17460 47549
rect 16948 47404 17000 47456
rect 17776 47404 17828 47456
rect 19524 47404 19576 47456
rect 25044 47583 25096 47592
rect 25044 47549 25053 47583
rect 25053 47549 25087 47583
rect 25087 47549 25096 47583
rect 25044 47540 25096 47549
rect 25320 47583 25372 47592
rect 25320 47549 25329 47583
rect 25329 47549 25363 47583
rect 25363 47549 25372 47583
rect 25320 47540 25372 47549
rect 20720 47404 20772 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 7472 47200 7524 47252
rect 18236 47200 18288 47252
rect 18512 47200 18564 47252
rect 19340 47243 19392 47252
rect 19340 47209 19349 47243
rect 19349 47209 19383 47243
rect 19383 47209 19392 47243
rect 19340 47200 19392 47209
rect 20536 47200 20588 47252
rect 17500 47132 17552 47184
rect 19892 47132 19944 47184
rect 10048 47107 10100 47116
rect 10048 47073 10057 47107
rect 10057 47073 10091 47107
rect 10091 47073 10100 47107
rect 10048 47064 10100 47073
rect 15476 47064 15528 47116
rect 16580 47064 16632 47116
rect 8944 46996 8996 47048
rect 18788 47107 18840 47116
rect 18788 47073 18797 47107
rect 18797 47073 18831 47107
rect 18831 47073 18840 47107
rect 18788 47064 18840 47073
rect 20076 47107 20128 47116
rect 20076 47073 20085 47107
rect 20085 47073 20119 47107
rect 20119 47073 20128 47107
rect 20076 47064 20128 47073
rect 20168 47107 20220 47116
rect 20168 47073 20177 47107
rect 20177 47073 20211 47107
rect 20211 47073 20220 47107
rect 20168 47064 20220 47073
rect 21548 47064 21600 47116
rect 10324 46971 10376 46980
rect 10324 46937 10333 46971
rect 10333 46937 10367 46971
rect 10367 46937 10376 46971
rect 10324 46928 10376 46937
rect 11060 46928 11112 46980
rect 18604 46996 18656 47048
rect 19616 46996 19668 47048
rect 22468 47132 22520 47184
rect 24124 47064 24176 47116
rect 11796 46903 11848 46912
rect 11796 46869 11805 46903
rect 11805 46869 11839 46903
rect 11839 46869 11848 46903
rect 11796 46860 11848 46869
rect 12808 46860 12860 46912
rect 14188 46903 14240 46912
rect 14188 46869 14197 46903
rect 14197 46869 14231 46903
rect 14231 46869 14240 46903
rect 14188 46860 14240 46869
rect 17132 46971 17184 46980
rect 17132 46937 17141 46971
rect 17141 46937 17175 46971
rect 17175 46937 17184 46971
rect 17132 46928 17184 46937
rect 18512 46971 18564 46980
rect 18512 46937 18521 46971
rect 18521 46937 18555 46971
rect 18555 46937 18564 46971
rect 18512 46928 18564 46937
rect 16856 46860 16908 46912
rect 17868 46860 17920 46912
rect 18880 46928 18932 46980
rect 21916 46928 21968 46980
rect 24492 46971 24544 46980
rect 24492 46937 24501 46971
rect 24501 46937 24535 46971
rect 24535 46937 24544 46971
rect 24492 46928 24544 46937
rect 25320 46860 25372 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 9036 46699 9088 46708
rect 9036 46665 9045 46699
rect 9045 46665 9079 46699
rect 9079 46665 9088 46699
rect 9036 46656 9088 46665
rect 9220 46656 9272 46708
rect 11060 46656 11112 46708
rect 6828 46588 6880 46640
rect 7380 46316 7432 46368
rect 9128 46520 9180 46572
rect 14096 46656 14148 46708
rect 14188 46588 14240 46640
rect 17408 46656 17460 46708
rect 18788 46656 18840 46708
rect 19156 46656 19208 46708
rect 15292 46588 15344 46640
rect 16120 46588 16172 46640
rect 16856 46588 16908 46640
rect 17868 46588 17920 46640
rect 23388 46656 23440 46708
rect 18604 46563 18656 46572
rect 18604 46529 18613 46563
rect 18613 46529 18647 46563
rect 18647 46529 18656 46563
rect 18604 46520 18656 46529
rect 22192 46588 22244 46640
rect 13820 46495 13872 46504
rect 13820 46461 13829 46495
rect 13829 46461 13863 46495
rect 13863 46461 13872 46495
rect 13820 46452 13872 46461
rect 12440 46316 12492 46368
rect 12532 46316 12584 46368
rect 16672 46452 16724 46504
rect 18328 46495 18380 46504
rect 18328 46461 18337 46495
rect 18337 46461 18371 46495
rect 18371 46461 18380 46495
rect 18328 46452 18380 46461
rect 21180 46452 21232 46504
rect 22560 46495 22612 46504
rect 22560 46461 22569 46495
rect 22569 46461 22603 46495
rect 22603 46461 22612 46495
rect 22560 46452 22612 46461
rect 22744 46563 22796 46572
rect 22744 46529 22753 46563
rect 22753 46529 22787 46563
rect 22787 46529 22796 46563
rect 22744 46520 22796 46529
rect 25964 46520 26016 46572
rect 23664 46452 23716 46504
rect 25320 46495 25372 46504
rect 25320 46461 25329 46495
rect 25329 46461 25363 46495
rect 25363 46461 25372 46495
rect 25320 46452 25372 46461
rect 17316 46316 17368 46368
rect 17592 46316 17644 46368
rect 19524 46316 19576 46368
rect 25044 46316 25096 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 11428 46155 11480 46164
rect 11428 46121 11437 46155
rect 11437 46121 11471 46155
rect 11471 46121 11480 46155
rect 11428 46112 11480 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 16212 46112 16264 46164
rect 16488 46112 16540 46164
rect 16672 46155 16724 46164
rect 16672 46121 16681 46155
rect 16681 46121 16715 46155
rect 16715 46121 16724 46155
rect 16672 46112 16724 46121
rect 17132 46112 17184 46164
rect 6184 46044 6236 46096
rect 8484 46044 8536 46096
rect 11796 45976 11848 46028
rect 12532 45976 12584 46028
rect 12716 45976 12768 46028
rect 16212 46019 16264 46028
rect 16212 45985 16221 46019
rect 16221 45985 16255 46019
rect 16255 45985 16264 46019
rect 16212 45976 16264 45985
rect 20628 45976 20680 46028
rect 21916 45976 21968 46028
rect 22376 45976 22428 46028
rect 17040 45908 17092 45960
rect 17592 45908 17644 45960
rect 24032 45951 24084 45960
rect 24032 45917 24041 45951
rect 24041 45917 24075 45951
rect 24075 45917 24084 45951
rect 24032 45908 24084 45917
rect 8760 45772 8812 45824
rect 11888 45840 11940 45892
rect 9680 45815 9732 45824
rect 9680 45781 9689 45815
rect 9689 45781 9723 45815
rect 9723 45781 9732 45815
rect 9680 45772 9732 45781
rect 11428 45772 11480 45824
rect 14188 45840 14240 45892
rect 14556 45840 14608 45892
rect 15384 45840 15436 45892
rect 16856 45840 16908 45892
rect 19248 45840 19300 45892
rect 20444 45840 20496 45892
rect 23664 45840 23716 45892
rect 24952 45840 25004 45892
rect 12808 45772 12860 45824
rect 13452 45772 13504 45824
rect 14924 45772 14976 45824
rect 16120 45772 16172 45824
rect 16580 45772 16632 45824
rect 20260 45815 20312 45824
rect 20260 45781 20269 45815
rect 20269 45781 20303 45815
rect 20303 45781 20312 45815
rect 20260 45772 20312 45781
rect 22376 45772 22428 45824
rect 23480 45772 23532 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 3976 45568 4028 45620
rect 9496 45568 9548 45620
rect 11060 45568 11112 45620
rect 13820 45568 13872 45620
rect 18328 45568 18380 45620
rect 8576 45500 8628 45552
rect 9312 45543 9364 45552
rect 9312 45509 9321 45543
rect 9321 45509 9355 45543
rect 9355 45509 9364 45543
rect 9312 45500 9364 45509
rect 11520 45500 11572 45552
rect 16856 45543 16908 45552
rect 16856 45509 16865 45543
rect 16865 45509 16899 45543
rect 16899 45509 16908 45543
rect 16856 45500 16908 45509
rect 20628 45500 20680 45552
rect 20720 45543 20772 45552
rect 20720 45509 20729 45543
rect 20729 45509 20763 45543
rect 20763 45509 20772 45543
rect 20720 45500 20772 45509
rect 23388 45500 23440 45552
rect 23480 45543 23532 45552
rect 23480 45509 23489 45543
rect 23489 45509 23523 45543
rect 23523 45509 23532 45543
rect 23480 45500 23532 45509
rect 12256 45432 12308 45484
rect 13728 45475 13780 45484
rect 13728 45441 13737 45475
rect 13737 45441 13771 45475
rect 13771 45441 13780 45475
rect 13728 45432 13780 45441
rect 14740 45432 14792 45484
rect 17408 45432 17460 45484
rect 18328 45432 18380 45484
rect 24032 45432 24084 45484
rect 6552 45228 6604 45280
rect 11244 45364 11296 45416
rect 13820 45407 13872 45416
rect 13820 45373 13829 45407
rect 13829 45373 13863 45407
rect 13863 45373 13872 45407
rect 13820 45364 13872 45373
rect 10324 45296 10376 45348
rect 12164 45296 12216 45348
rect 13544 45296 13596 45348
rect 13636 45296 13688 45348
rect 21180 45364 21232 45416
rect 24492 45407 24544 45416
rect 24492 45373 24501 45407
rect 24501 45373 24535 45407
rect 24535 45373 24544 45407
rect 24492 45364 24544 45373
rect 24768 45407 24820 45416
rect 24768 45373 24777 45407
rect 24777 45373 24811 45407
rect 24811 45373 24820 45407
rect 24768 45364 24820 45373
rect 10048 45228 10100 45280
rect 12256 45271 12308 45280
rect 12256 45237 12265 45271
rect 12265 45237 12299 45271
rect 12299 45237 12308 45271
rect 12256 45228 12308 45237
rect 15384 45228 15436 45280
rect 15568 45228 15620 45280
rect 19156 45228 19208 45280
rect 21916 45228 21968 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 6092 45067 6144 45076
rect 6092 45033 6101 45067
rect 6101 45033 6135 45067
rect 6135 45033 6144 45067
rect 6092 45024 6144 45033
rect 6644 45067 6696 45076
rect 6644 45033 6653 45067
rect 6653 45033 6687 45067
rect 6687 45033 6696 45067
rect 6644 45024 6696 45033
rect 7840 45024 7892 45076
rect 8668 45024 8720 45076
rect 12072 45067 12124 45076
rect 12072 45033 12081 45067
rect 12081 45033 12115 45067
rect 12115 45033 12124 45067
rect 12072 45024 12124 45033
rect 16580 45024 16632 45076
rect 7288 44999 7340 45008
rect 7288 44965 7297 44999
rect 7297 44965 7331 44999
rect 7331 44965 7340 44999
rect 7288 44956 7340 44965
rect 8852 44956 8904 45008
rect 10876 44956 10928 45008
rect 5908 44863 5960 44872
rect 5908 44829 5917 44863
rect 5917 44829 5951 44863
rect 5951 44829 5960 44863
rect 5908 44820 5960 44829
rect 7656 44820 7708 44872
rect 12532 44820 12584 44872
rect 13636 44820 13688 44872
rect 6644 44752 6696 44804
rect 7288 44752 7340 44804
rect 8484 44752 8536 44804
rect 10508 44795 10560 44804
rect 10508 44761 10517 44795
rect 10517 44761 10551 44795
rect 10551 44761 10560 44795
rect 10508 44752 10560 44761
rect 11244 44795 11296 44804
rect 11244 44761 11253 44795
rect 11253 44761 11287 44795
rect 11287 44761 11296 44795
rect 11244 44752 11296 44761
rect 14280 44752 14332 44804
rect 12808 44684 12860 44736
rect 15568 44795 15620 44804
rect 15568 44761 15577 44795
rect 15577 44761 15611 44795
rect 15611 44761 15620 44795
rect 15568 44752 15620 44761
rect 20168 45024 20220 45076
rect 24952 45024 25004 45076
rect 19524 44956 19576 45008
rect 18880 44863 18932 44872
rect 18880 44829 18889 44863
rect 18889 44829 18923 44863
rect 18923 44829 18932 44863
rect 18880 44820 18932 44829
rect 21180 44863 21232 44872
rect 21180 44829 21189 44863
rect 21189 44829 21223 44863
rect 21223 44829 21232 44863
rect 21180 44820 21232 44829
rect 22008 44820 22060 44872
rect 24032 44888 24084 44940
rect 17592 44752 17644 44804
rect 20628 44752 20680 44804
rect 21364 44752 21416 44804
rect 21548 44752 21600 44804
rect 23480 44752 23532 44804
rect 16212 44684 16264 44736
rect 16488 44684 16540 44736
rect 17040 44727 17092 44736
rect 17040 44693 17049 44727
rect 17049 44693 17083 44727
rect 17083 44693 17092 44727
rect 17040 44684 17092 44693
rect 21272 44684 21324 44736
rect 21824 44727 21876 44736
rect 21824 44693 21833 44727
rect 21833 44693 21867 44727
rect 21867 44693 21876 44727
rect 21824 44684 21876 44693
rect 22744 44684 22796 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 6000 44480 6052 44532
rect 9496 44480 9548 44532
rect 11888 44523 11940 44532
rect 11888 44489 11897 44523
rect 11897 44489 11931 44523
rect 11931 44489 11940 44523
rect 11888 44480 11940 44489
rect 14372 44480 14424 44532
rect 21364 44523 21416 44532
rect 21364 44489 21373 44523
rect 21373 44489 21407 44523
rect 21407 44489 21416 44523
rect 21364 44480 21416 44489
rect 21824 44480 21876 44532
rect 23296 44480 23348 44532
rect 6460 44412 6512 44464
rect 8392 44412 8444 44464
rect 17592 44412 17644 44464
rect 21916 44412 21968 44464
rect 6828 44344 6880 44396
rect 9220 44387 9272 44396
rect 9220 44353 9229 44387
rect 9229 44353 9263 44387
rect 9263 44353 9272 44387
rect 9220 44344 9272 44353
rect 14556 44344 14608 44396
rect 14924 44344 14976 44396
rect 16672 44344 16724 44396
rect 19156 44344 19208 44396
rect 20168 44344 20220 44396
rect 12348 44319 12400 44328
rect 12348 44285 12357 44319
rect 12357 44285 12391 44319
rect 12391 44285 12400 44319
rect 12348 44276 12400 44285
rect 11612 44251 11664 44260
rect 11612 44217 11621 44251
rect 11621 44217 11655 44251
rect 11655 44217 11664 44251
rect 11612 44208 11664 44217
rect 12256 44208 12308 44260
rect 12716 44276 12768 44328
rect 13452 44319 13504 44328
rect 13452 44285 13461 44319
rect 13461 44285 13495 44319
rect 13495 44285 13504 44319
rect 13452 44276 13504 44285
rect 16488 44276 16540 44328
rect 17132 44319 17184 44328
rect 17132 44285 17141 44319
rect 17141 44285 17175 44319
rect 17175 44285 17184 44319
rect 17132 44276 17184 44285
rect 17776 44276 17828 44328
rect 23572 44276 23624 44328
rect 24676 44276 24728 44328
rect 24768 44319 24820 44328
rect 24768 44285 24777 44319
rect 24777 44285 24811 44319
rect 24811 44285 24820 44319
rect 24768 44276 24820 44285
rect 7288 44140 7340 44192
rect 14740 44140 14792 44192
rect 15200 44140 15252 44192
rect 18328 44140 18380 44192
rect 19616 44140 19668 44192
rect 22100 44183 22152 44192
rect 22100 44149 22109 44183
rect 22109 44149 22143 44183
rect 22143 44149 22152 44183
rect 22100 44140 22152 44149
rect 22836 44140 22888 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 7564 43936 7616 43988
rect 9404 43936 9456 43988
rect 12348 43936 12400 43988
rect 13820 43936 13872 43988
rect 15568 43936 15620 43988
rect 9312 43843 9364 43852
rect 9312 43809 9321 43843
rect 9321 43809 9355 43843
rect 9355 43809 9364 43843
rect 9312 43800 9364 43809
rect 9496 43843 9548 43852
rect 9496 43809 9505 43843
rect 9505 43809 9539 43843
rect 9539 43809 9548 43843
rect 9496 43800 9548 43809
rect 10968 43868 11020 43920
rect 16120 43868 16172 43920
rect 12624 43843 12676 43852
rect 12624 43809 12633 43843
rect 12633 43809 12667 43843
rect 12667 43809 12676 43843
rect 12624 43800 12676 43809
rect 10232 43732 10284 43784
rect 14740 43800 14792 43852
rect 17684 43843 17736 43852
rect 17684 43809 17693 43843
rect 17693 43809 17727 43843
rect 17727 43809 17736 43843
rect 17684 43800 17736 43809
rect 22652 43936 22704 43988
rect 19340 43868 19392 43920
rect 10784 43664 10836 43716
rect 16856 43664 16908 43716
rect 21088 43800 21140 43852
rect 22836 43868 22888 43920
rect 23480 43979 23532 43988
rect 23480 43945 23489 43979
rect 23489 43945 23523 43979
rect 23523 43945 23532 43979
rect 23480 43936 23532 43945
rect 25688 43868 25740 43920
rect 22744 43800 22796 43852
rect 24676 43800 24728 43852
rect 22192 43732 22244 43784
rect 24032 43732 24084 43784
rect 12348 43639 12400 43648
rect 12348 43605 12357 43639
rect 12357 43605 12391 43639
rect 12391 43605 12400 43639
rect 12348 43596 12400 43605
rect 14924 43639 14976 43648
rect 14924 43605 14933 43639
rect 14933 43605 14967 43639
rect 14967 43605 14976 43639
rect 14924 43596 14976 43605
rect 15844 43639 15896 43648
rect 15844 43605 15853 43639
rect 15853 43605 15887 43639
rect 15887 43605 15896 43639
rect 15844 43596 15896 43605
rect 17224 43639 17276 43648
rect 17224 43605 17233 43639
rect 17233 43605 17267 43639
rect 17267 43605 17276 43639
rect 17224 43596 17276 43605
rect 17776 43596 17828 43648
rect 19708 43639 19760 43648
rect 19708 43605 19717 43639
rect 19717 43605 19751 43639
rect 19751 43605 19760 43639
rect 19708 43596 19760 43605
rect 20628 43664 20680 43716
rect 22008 43664 22060 43716
rect 23664 43664 23716 43716
rect 21272 43596 21324 43648
rect 22468 43596 22520 43648
rect 22652 43639 22704 43648
rect 22652 43605 22661 43639
rect 22661 43605 22695 43639
rect 22695 43605 22704 43639
rect 22652 43596 22704 43605
rect 23480 43596 23532 43648
rect 24584 43596 24636 43648
rect 24952 43596 25004 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 7748 43392 7800 43444
rect 12808 43392 12860 43444
rect 15476 43392 15528 43444
rect 9404 43324 9456 43376
rect 10048 43324 10100 43376
rect 1308 43256 1360 43308
rect 7840 43256 7892 43308
rect 10416 43299 10468 43308
rect 10416 43265 10425 43299
rect 10425 43265 10459 43299
rect 10459 43265 10468 43299
rect 10416 43256 10468 43265
rect 14832 43256 14884 43308
rect 11060 43188 11112 43240
rect 11152 43231 11204 43240
rect 11152 43197 11161 43231
rect 11161 43197 11195 43231
rect 11195 43197 11204 43231
rect 11152 43188 11204 43197
rect 12716 43231 12768 43240
rect 12716 43197 12725 43231
rect 12725 43197 12759 43231
rect 12759 43197 12768 43231
rect 12716 43188 12768 43197
rect 15476 43231 15528 43240
rect 15476 43197 15485 43231
rect 15485 43197 15519 43231
rect 15519 43197 15528 43231
rect 15476 43188 15528 43197
rect 15568 43231 15620 43240
rect 15568 43197 15577 43231
rect 15577 43197 15611 43231
rect 15611 43197 15620 43231
rect 15568 43188 15620 43197
rect 3792 43120 3844 43172
rect 15292 43120 15344 43172
rect 16580 43392 16632 43444
rect 17500 43392 17552 43444
rect 19432 43392 19484 43444
rect 19708 43392 19760 43444
rect 17776 43256 17828 43308
rect 22284 43435 22336 43444
rect 22284 43401 22293 43435
rect 22293 43401 22327 43435
rect 22327 43401 22336 43435
rect 22284 43392 22336 43401
rect 22376 43392 22428 43444
rect 17132 43231 17184 43240
rect 17132 43197 17141 43231
rect 17141 43197 17175 43231
rect 17175 43197 17184 43231
rect 17132 43188 17184 43197
rect 17868 43188 17920 43240
rect 21364 43256 21416 43308
rect 21732 43256 21784 43308
rect 23388 43392 23440 43444
rect 24952 43367 25004 43376
rect 24952 43333 24961 43367
rect 24961 43333 24995 43367
rect 24995 43333 25004 43367
rect 24952 43324 25004 43333
rect 23848 43256 23900 43308
rect 19524 43188 19576 43240
rect 19616 43231 19668 43240
rect 19616 43197 19625 43231
rect 19625 43197 19659 43231
rect 19659 43197 19668 43231
rect 19616 43188 19668 43197
rect 18420 43120 18472 43172
rect 22468 43188 22520 43240
rect 22376 43120 22428 43172
rect 3516 43052 3568 43104
rect 8668 43095 8720 43104
rect 8668 43061 8677 43095
rect 8677 43061 8711 43095
rect 8711 43061 8720 43095
rect 8668 43052 8720 43061
rect 12808 43052 12860 43104
rect 13452 43052 13504 43104
rect 15108 43052 15160 43104
rect 18880 43052 18932 43104
rect 19524 43052 19576 43104
rect 20628 43052 20680 43104
rect 20996 43095 21048 43104
rect 20996 43061 21005 43095
rect 21005 43061 21039 43095
rect 21039 43061 21048 43095
rect 20996 43052 21048 43061
rect 21364 43095 21416 43104
rect 21364 43061 21373 43095
rect 21373 43061 21407 43095
rect 21407 43061 21416 43095
rect 21364 43052 21416 43061
rect 21456 43052 21508 43104
rect 23388 43120 23440 43172
rect 25320 43188 25372 43240
rect 26056 43120 26108 43172
rect 23296 43052 23348 43104
rect 23572 43052 23624 43104
rect 24308 43052 24360 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 14924 42848 14976 42900
rect 17500 42848 17552 42900
rect 19708 42848 19760 42900
rect 13452 42780 13504 42832
rect 4804 42712 4856 42764
rect 5448 42712 5500 42764
rect 10416 42712 10468 42764
rect 12624 42712 12676 42764
rect 17316 42712 17368 42764
rect 19616 42780 19668 42832
rect 20260 42712 20312 42764
rect 21548 42780 21600 42832
rect 21732 42780 21784 42832
rect 23572 42780 23624 42832
rect 25780 42780 25832 42832
rect 21272 42755 21324 42764
rect 21272 42721 21281 42755
rect 21281 42721 21315 42755
rect 21315 42721 21324 42755
rect 21272 42712 21324 42721
rect 22008 42712 22060 42764
rect 25320 42712 25372 42764
rect 8576 42687 8628 42696
rect 8576 42653 8585 42687
rect 8585 42653 8619 42687
rect 8619 42653 8628 42687
rect 8576 42644 8628 42653
rect 14188 42644 14240 42696
rect 16764 42644 16816 42696
rect 21456 42644 21508 42696
rect 24032 42644 24084 42696
rect 25228 42687 25280 42696
rect 25228 42653 25237 42687
rect 25237 42653 25271 42687
rect 25271 42653 25280 42687
rect 25228 42644 25280 42653
rect 5264 42551 5316 42560
rect 5264 42517 5273 42551
rect 5273 42517 5307 42551
rect 5307 42517 5316 42551
rect 5264 42508 5316 42517
rect 11244 42576 11296 42628
rect 11336 42619 11388 42628
rect 11336 42585 11345 42619
rect 11345 42585 11379 42619
rect 11379 42585 11388 42619
rect 11336 42576 11388 42585
rect 12624 42576 12676 42628
rect 6368 42551 6420 42560
rect 6368 42517 6377 42551
rect 6377 42517 6411 42551
rect 6411 42517 6420 42551
rect 6368 42508 6420 42517
rect 7748 42508 7800 42560
rect 8944 42508 8996 42560
rect 9404 42508 9456 42560
rect 9588 42551 9640 42560
rect 9588 42517 9597 42551
rect 9597 42517 9631 42551
rect 9631 42517 9640 42551
rect 9588 42508 9640 42517
rect 13360 42551 13412 42560
rect 13360 42517 13369 42551
rect 13369 42517 13403 42551
rect 13403 42517 13412 42551
rect 13360 42508 13412 42517
rect 15660 42576 15712 42628
rect 14832 42508 14884 42560
rect 15844 42508 15896 42560
rect 19800 42576 19852 42628
rect 20536 42576 20588 42628
rect 20628 42576 20680 42628
rect 19984 42551 20036 42560
rect 19984 42517 19993 42551
rect 19993 42517 20027 42551
rect 20027 42517 20036 42551
rect 19984 42508 20036 42517
rect 20352 42551 20404 42560
rect 20352 42517 20361 42551
rect 20361 42517 20395 42551
rect 20395 42517 20404 42551
rect 20352 42508 20404 42517
rect 22192 42508 22244 42560
rect 23848 42576 23900 42628
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 4988 42347 5040 42356
rect 4988 42313 4997 42347
rect 4997 42313 5031 42347
rect 5031 42313 5040 42347
rect 4988 42304 5040 42313
rect 11336 42304 11388 42356
rect 11704 42347 11756 42356
rect 11704 42313 11713 42347
rect 11713 42313 11747 42347
rect 11747 42313 11756 42347
rect 11704 42304 11756 42313
rect 13360 42347 13412 42356
rect 13360 42313 13369 42347
rect 13369 42313 13403 42347
rect 13403 42313 13412 42347
rect 13360 42304 13412 42313
rect 13728 42347 13780 42356
rect 13728 42313 13737 42347
rect 13737 42313 13771 42347
rect 13771 42313 13780 42347
rect 13728 42304 13780 42313
rect 14372 42304 14424 42356
rect 18788 42304 18840 42356
rect 3424 42279 3476 42288
rect 3424 42245 3433 42279
rect 3433 42245 3467 42279
rect 3467 42245 3476 42279
rect 3424 42236 3476 42245
rect 3884 42236 3936 42288
rect 4344 42211 4396 42220
rect 4344 42177 4353 42211
rect 4353 42177 4387 42211
rect 4387 42177 4396 42211
rect 4344 42168 4396 42177
rect 8392 42236 8444 42288
rect 4896 42100 4948 42152
rect 9220 42168 9272 42220
rect 9496 42168 9548 42220
rect 11796 42168 11848 42220
rect 7748 42100 7800 42152
rect 14740 42236 14792 42288
rect 14924 42236 14976 42288
rect 16212 42236 16264 42288
rect 19800 42304 19852 42356
rect 13728 42168 13780 42220
rect 15568 42168 15620 42220
rect 16580 42168 16632 42220
rect 13360 42100 13412 42152
rect 20628 42236 20680 42288
rect 21272 42304 21324 42356
rect 22560 42304 22612 42356
rect 23848 42236 23900 42288
rect 24400 42279 24452 42288
rect 24400 42245 24409 42279
rect 24409 42245 24443 42279
rect 24443 42245 24452 42279
rect 24400 42236 24452 42245
rect 21824 42168 21876 42220
rect 22560 42211 22612 42220
rect 22560 42177 22569 42211
rect 22569 42177 22603 42211
rect 22603 42177 22612 42211
rect 22560 42168 22612 42177
rect 14740 42032 14792 42084
rect 6184 41964 6236 42016
rect 10508 41964 10560 42016
rect 13912 41964 13964 42016
rect 15476 42007 15528 42016
rect 15476 41973 15485 42007
rect 15485 41973 15519 42007
rect 15519 41973 15528 42007
rect 15476 41964 15528 41973
rect 15844 41964 15896 42016
rect 20996 42100 21048 42152
rect 22836 42100 22888 42152
rect 20076 42032 20128 42084
rect 24860 42032 24912 42084
rect 25320 42032 25372 42084
rect 18972 41964 19024 42016
rect 19432 41964 19484 42016
rect 20168 41964 20220 42016
rect 20904 42007 20956 42016
rect 20904 41973 20913 42007
rect 20913 41973 20947 42007
rect 20947 41973 20956 42007
rect 20904 41964 20956 41973
rect 22560 41964 22612 42016
rect 23204 41964 23256 42016
rect 25412 41964 25464 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 4344 41760 4396 41812
rect 8576 41760 8628 41812
rect 9496 41760 9548 41812
rect 3700 41692 3752 41744
rect 8392 41624 8444 41676
rect 7564 41556 7616 41608
rect 9220 41624 9272 41676
rect 12624 41760 12676 41812
rect 14372 41760 14424 41812
rect 16672 41760 16724 41812
rect 17592 41760 17644 41812
rect 22560 41760 22612 41812
rect 15200 41624 15252 41676
rect 16580 41624 16632 41676
rect 16948 41667 17000 41676
rect 16948 41633 16957 41667
rect 16957 41633 16991 41667
rect 16991 41633 17000 41667
rect 16948 41624 17000 41633
rect 11704 41556 11756 41608
rect 12716 41556 12768 41608
rect 14188 41556 14240 41608
rect 15660 41556 15712 41608
rect 17868 41624 17920 41676
rect 19432 41624 19484 41676
rect 22008 41624 22060 41676
rect 22744 41624 22796 41676
rect 17316 41556 17368 41608
rect 20720 41556 20772 41608
rect 20812 41599 20864 41608
rect 20812 41565 20821 41599
rect 20821 41565 20855 41599
rect 20855 41565 20864 41599
rect 20812 41556 20864 41565
rect 22836 41556 22888 41608
rect 24492 41692 24544 41744
rect 25228 41760 25280 41812
rect 23848 41624 23900 41676
rect 24768 41624 24820 41676
rect 25044 41667 25096 41676
rect 25044 41633 25053 41667
rect 25053 41633 25087 41667
rect 25087 41633 25096 41667
rect 25044 41624 25096 41633
rect 5080 41531 5132 41540
rect 5080 41497 5089 41531
rect 5089 41497 5123 41531
rect 5123 41497 5132 41531
rect 5080 41488 5132 41497
rect 6552 41531 6604 41540
rect 6552 41497 6561 41531
rect 6561 41497 6595 41531
rect 6595 41497 6604 41531
rect 6552 41488 6604 41497
rect 11244 41488 11296 41540
rect 12072 41531 12124 41540
rect 12072 41497 12081 41531
rect 12081 41497 12115 41531
rect 12115 41497 12124 41531
rect 12072 41488 12124 41497
rect 20904 41488 20956 41540
rect 21272 41488 21324 41540
rect 21548 41488 21600 41540
rect 25044 41488 25096 41540
rect 25596 41488 25648 41540
rect 16396 41420 16448 41472
rect 17592 41420 17644 41472
rect 18512 41420 18564 41472
rect 20996 41463 21048 41472
rect 20996 41429 21005 41463
rect 21005 41429 21039 41463
rect 21039 41429 21048 41463
rect 20996 41420 21048 41429
rect 22468 41420 22520 41472
rect 22744 41420 22796 41472
rect 22836 41463 22888 41472
rect 22836 41429 22845 41463
rect 22845 41429 22879 41463
rect 22879 41429 22888 41463
rect 22836 41420 22888 41429
rect 24216 41463 24268 41472
rect 24216 41429 24225 41463
rect 24225 41429 24259 41463
rect 24259 41429 24268 41463
rect 24216 41420 24268 41429
rect 24584 41463 24636 41472
rect 24584 41429 24593 41463
rect 24593 41429 24627 41463
rect 24627 41429 24636 41463
rect 24584 41420 24636 41429
rect 24952 41463 25004 41472
rect 24952 41429 24961 41463
rect 24961 41429 24995 41463
rect 24995 41429 25004 41463
rect 24952 41420 25004 41429
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 4068 41216 4120 41268
rect 10968 41216 11020 41268
rect 7564 41148 7616 41200
rect 10416 41191 10468 41200
rect 1308 41080 1360 41132
rect 8116 41055 8168 41064
rect 8116 41021 8125 41055
rect 8125 41021 8159 41055
rect 8159 41021 8168 41055
rect 8116 41012 8168 41021
rect 8392 41055 8444 41064
rect 8392 41021 8401 41055
rect 8401 41021 8435 41055
rect 8435 41021 8444 41055
rect 10416 41157 10425 41191
rect 10425 41157 10459 41191
rect 10459 41157 10468 41191
rect 10416 41148 10468 41157
rect 10600 41080 10652 41132
rect 12072 41216 12124 41268
rect 13728 41216 13780 41268
rect 13820 41216 13872 41268
rect 14832 41216 14884 41268
rect 15844 41216 15896 41268
rect 17224 41216 17276 41268
rect 18420 41216 18472 41268
rect 18696 41216 18748 41268
rect 19064 41216 19116 41268
rect 19892 41259 19944 41268
rect 19892 41225 19901 41259
rect 19901 41225 19935 41259
rect 19935 41225 19944 41259
rect 19892 41216 19944 41225
rect 19984 41216 20036 41268
rect 20812 41216 20864 41268
rect 22008 41216 22060 41268
rect 22652 41259 22704 41268
rect 22652 41225 22661 41259
rect 22661 41225 22695 41259
rect 22695 41225 22704 41259
rect 22652 41216 22704 41225
rect 22836 41216 22888 41268
rect 23940 41216 23992 41268
rect 11428 41148 11480 41200
rect 8392 41012 8444 41021
rect 9312 41012 9364 41064
rect 10692 41012 10744 41064
rect 3424 40944 3476 40996
rect 8852 40987 8904 40996
rect 3700 40876 3752 40928
rect 6644 40919 6696 40928
rect 6644 40885 6653 40919
rect 6653 40885 6687 40919
rect 6687 40885 6696 40919
rect 6644 40876 6696 40885
rect 8852 40953 8861 40987
rect 8861 40953 8895 40987
rect 8895 40953 8904 40987
rect 8852 40944 8904 40953
rect 10140 40944 10192 40996
rect 11612 40944 11664 40996
rect 12256 41055 12308 41064
rect 12256 41021 12265 41055
rect 12265 41021 12299 41055
rect 12299 41021 12308 41055
rect 12256 41012 12308 41021
rect 13452 41080 13504 41132
rect 13636 41080 13688 41132
rect 16488 41148 16540 41200
rect 18972 41148 19024 41200
rect 15292 41080 15344 41132
rect 13544 40944 13596 40996
rect 9220 40876 9272 40928
rect 10416 40876 10468 40928
rect 11428 40876 11480 40928
rect 11980 40876 12032 40928
rect 13452 40876 13504 40928
rect 15476 41012 15528 41064
rect 15568 41055 15620 41064
rect 15568 41021 15577 41055
rect 15577 41021 15611 41055
rect 15611 41021 15620 41055
rect 15568 41012 15620 41021
rect 15936 41080 15988 41132
rect 18604 41123 18656 41132
rect 18604 41089 18613 41123
rect 18613 41089 18647 41123
rect 18647 41089 18656 41123
rect 18604 41080 18656 41089
rect 17040 41055 17092 41064
rect 17040 41021 17049 41055
rect 17049 41021 17083 41055
rect 17083 41021 17092 41055
rect 17040 41012 17092 41021
rect 18328 41055 18380 41064
rect 18328 41021 18337 41055
rect 18337 41021 18371 41055
rect 18371 41021 18380 41055
rect 18328 41012 18380 41021
rect 19892 41080 19944 41132
rect 21180 41148 21232 41200
rect 19156 41012 19208 41064
rect 22468 41080 22520 41132
rect 24492 41123 24544 41132
rect 24492 41089 24501 41123
rect 24501 41089 24535 41123
rect 24535 41089 24544 41123
rect 24492 41080 24544 41089
rect 21088 41055 21140 41064
rect 21088 41021 21097 41055
rect 21097 41021 21131 41055
rect 21131 41021 21140 41055
rect 21088 41012 21140 41021
rect 21916 41012 21968 41064
rect 22744 41012 22796 41064
rect 23756 41055 23808 41064
rect 23756 41021 23765 41055
rect 23765 41021 23799 41055
rect 23799 41021 23808 41055
rect 23756 41012 23808 41021
rect 15292 40876 15344 40928
rect 16304 40876 16356 40928
rect 17592 40919 17644 40928
rect 17592 40885 17601 40919
rect 17601 40885 17635 40919
rect 17635 40885 17644 40919
rect 17592 40876 17644 40885
rect 18696 40876 18748 40928
rect 19432 40919 19484 40928
rect 19432 40885 19441 40919
rect 19441 40885 19475 40919
rect 19475 40885 19484 40919
rect 19432 40876 19484 40885
rect 21088 40876 21140 40928
rect 21456 40876 21508 40928
rect 22008 40944 22060 40996
rect 22468 40876 22520 40928
rect 24860 40876 24912 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 8116 40672 8168 40724
rect 10968 40672 11020 40724
rect 7104 40604 7156 40656
rect 10416 40604 10468 40656
rect 13544 40672 13596 40724
rect 13728 40672 13780 40724
rect 14004 40672 14056 40724
rect 14740 40672 14792 40724
rect 17316 40672 17368 40724
rect 22468 40672 22520 40724
rect 25136 40672 25188 40724
rect 9036 40536 9088 40588
rect 14464 40604 14516 40656
rect 16764 40604 16816 40656
rect 21732 40604 21784 40656
rect 22008 40604 22060 40656
rect 7196 40468 7248 40520
rect 12072 40536 12124 40588
rect 14004 40536 14056 40588
rect 14832 40536 14884 40588
rect 16304 40579 16356 40588
rect 16304 40545 16313 40579
rect 16313 40545 16347 40579
rect 16347 40545 16356 40579
rect 16304 40536 16356 40545
rect 11980 40511 12032 40520
rect 11980 40477 11989 40511
rect 11989 40477 12023 40511
rect 12023 40477 12032 40511
rect 11980 40468 12032 40477
rect 12532 40468 12584 40520
rect 13452 40468 13504 40520
rect 17408 40536 17460 40588
rect 18512 40536 18564 40588
rect 18972 40536 19024 40588
rect 20720 40536 20772 40588
rect 21916 40536 21968 40588
rect 22560 40536 22612 40588
rect 8852 40400 8904 40452
rect 10784 40443 10836 40452
rect 10784 40409 10793 40443
rect 10793 40409 10827 40443
rect 10827 40409 10836 40443
rect 10784 40400 10836 40409
rect 11244 40400 11296 40452
rect 14556 40400 14608 40452
rect 14924 40400 14976 40452
rect 9036 40332 9088 40384
rect 9312 40332 9364 40384
rect 10324 40332 10376 40384
rect 10416 40375 10468 40384
rect 10416 40341 10425 40375
rect 10425 40341 10459 40375
rect 10459 40341 10468 40375
rect 10416 40332 10468 40341
rect 10968 40332 11020 40384
rect 11060 40332 11112 40384
rect 11428 40332 11480 40384
rect 12716 40332 12768 40384
rect 13544 40375 13596 40384
rect 13544 40341 13553 40375
rect 13553 40341 13587 40375
rect 13587 40341 13596 40375
rect 13544 40332 13596 40341
rect 17868 40400 17920 40452
rect 18512 40400 18564 40452
rect 20444 40468 20496 40520
rect 21180 40511 21232 40520
rect 21180 40477 21189 40511
rect 21189 40477 21223 40511
rect 21223 40477 21232 40511
rect 21180 40468 21232 40477
rect 21640 40468 21692 40520
rect 22192 40468 22244 40520
rect 23756 40468 23808 40520
rect 19892 40400 19944 40452
rect 18972 40332 19024 40384
rect 19524 40332 19576 40384
rect 21088 40375 21140 40384
rect 21088 40341 21097 40375
rect 21097 40341 21131 40375
rect 21131 40341 21140 40375
rect 21088 40332 21140 40341
rect 21732 40400 21784 40452
rect 25504 40536 25556 40588
rect 24216 40468 24268 40520
rect 24492 40468 24544 40520
rect 22468 40332 22520 40384
rect 24308 40400 24360 40452
rect 23296 40375 23348 40384
rect 23296 40341 23305 40375
rect 23305 40341 23339 40375
rect 23339 40341 23348 40375
rect 23296 40332 23348 40341
rect 25228 40375 25280 40384
rect 25228 40341 25237 40375
rect 25237 40341 25271 40375
rect 25271 40341 25280 40375
rect 25228 40332 25280 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 11060 40128 11112 40180
rect 11336 40128 11388 40180
rect 13452 40171 13504 40180
rect 13452 40137 13461 40171
rect 13461 40137 13495 40171
rect 13495 40137 13504 40171
rect 13452 40128 13504 40137
rect 15936 40128 15988 40180
rect 16856 40171 16908 40180
rect 16856 40137 16865 40171
rect 16865 40137 16899 40171
rect 16899 40137 16908 40171
rect 16856 40128 16908 40137
rect 19432 40128 19484 40180
rect 19984 40171 20036 40180
rect 19984 40137 19993 40171
rect 19993 40137 20027 40171
rect 20027 40137 20036 40171
rect 19984 40128 20036 40137
rect 9036 40060 9088 40112
rect 9220 40060 9272 40112
rect 11980 40103 12032 40112
rect 11980 40069 11989 40103
rect 11989 40069 12023 40103
rect 12023 40069 12032 40103
rect 11980 40060 12032 40069
rect 13636 40060 13688 40112
rect 16764 40060 16816 40112
rect 17776 40060 17828 40112
rect 18328 40060 18380 40112
rect 11704 40035 11756 40044
rect 11704 40001 11713 40035
rect 11713 40001 11747 40035
rect 11747 40001 11756 40035
rect 11704 39992 11756 40001
rect 10508 39924 10560 39976
rect 15384 39992 15436 40044
rect 17316 40035 17368 40044
rect 17316 40001 17325 40035
rect 17325 40001 17359 40035
rect 17359 40001 17368 40035
rect 17316 39992 17368 40001
rect 21364 40128 21416 40180
rect 24952 40128 25004 40180
rect 20996 40060 21048 40112
rect 21916 40060 21968 40112
rect 14832 39967 14884 39976
rect 14832 39933 14841 39967
rect 14841 39933 14875 39967
rect 14875 39933 14884 39967
rect 14832 39924 14884 39933
rect 15936 39924 15988 39976
rect 22192 39992 22244 40044
rect 18880 39924 18932 39976
rect 21640 39924 21692 39976
rect 22008 39924 22060 39976
rect 24768 40060 24820 40112
rect 25320 40035 25372 40044
rect 25320 40001 25329 40035
rect 25329 40001 25363 40035
rect 25363 40001 25372 40035
rect 25320 39992 25372 40001
rect 6644 39788 6696 39840
rect 8576 39788 8628 39840
rect 10968 39788 11020 39840
rect 11244 39831 11296 39840
rect 11244 39797 11253 39831
rect 11253 39797 11287 39831
rect 11287 39797 11296 39831
rect 11244 39788 11296 39797
rect 11520 39788 11572 39840
rect 17684 39856 17736 39908
rect 13452 39788 13504 39840
rect 14832 39788 14884 39840
rect 14924 39788 14976 39840
rect 16948 39788 17000 39840
rect 20260 39831 20312 39840
rect 20260 39797 20269 39831
rect 20269 39797 20303 39831
rect 20303 39797 20312 39831
rect 20260 39788 20312 39797
rect 22192 39856 22244 39908
rect 25044 39967 25096 39976
rect 25044 39933 25053 39967
rect 25053 39933 25087 39967
rect 25087 39933 25096 39967
rect 25044 39924 25096 39933
rect 22560 39788 22612 39840
rect 23572 39788 23624 39840
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 7196 39627 7248 39636
rect 7196 39593 7205 39627
rect 7205 39593 7239 39627
rect 7239 39593 7248 39627
rect 7196 39584 7248 39593
rect 7564 39627 7616 39636
rect 7564 39593 7573 39627
rect 7573 39593 7607 39627
rect 7607 39593 7616 39627
rect 7564 39584 7616 39593
rect 9128 39627 9180 39636
rect 9128 39593 9137 39627
rect 9137 39593 9171 39627
rect 9171 39593 9180 39627
rect 9128 39584 9180 39593
rect 11244 39584 11296 39636
rect 12348 39584 12400 39636
rect 12440 39516 12492 39568
rect 15568 39584 15620 39636
rect 18604 39584 18656 39636
rect 20260 39584 20312 39636
rect 25044 39584 25096 39636
rect 8300 39448 8352 39500
rect 11520 39448 11572 39500
rect 11980 39448 12032 39500
rect 12716 39516 12768 39568
rect 14096 39516 14148 39568
rect 16672 39516 16724 39568
rect 17868 39516 17920 39568
rect 5448 39423 5500 39432
rect 5448 39389 5457 39423
rect 5457 39389 5491 39423
rect 5491 39389 5500 39423
rect 5448 39380 5500 39389
rect 9588 39380 9640 39432
rect 11152 39423 11204 39432
rect 11152 39389 11161 39423
rect 11161 39389 11195 39423
rect 11195 39389 11204 39423
rect 11152 39380 11204 39389
rect 12992 39448 13044 39500
rect 16488 39448 16540 39500
rect 17132 39448 17184 39500
rect 15568 39380 15620 39432
rect 19432 39448 19484 39500
rect 20260 39491 20312 39500
rect 20260 39457 20269 39491
rect 20269 39457 20303 39491
rect 20303 39457 20312 39491
rect 20260 39448 20312 39457
rect 22284 39516 22336 39568
rect 22652 39516 22704 39568
rect 23756 39448 23808 39500
rect 17408 39380 17460 39432
rect 21180 39380 21232 39432
rect 21640 39380 21692 39432
rect 24676 39423 24728 39432
rect 24676 39389 24685 39423
rect 24685 39389 24719 39423
rect 24719 39389 24728 39423
rect 24676 39380 24728 39389
rect 5356 39312 5408 39364
rect 7564 39312 7616 39364
rect 8760 39244 8812 39296
rect 9496 39287 9548 39296
rect 9496 39253 9505 39287
rect 9505 39253 9539 39287
rect 9539 39253 9548 39287
rect 9496 39244 9548 39253
rect 9588 39287 9640 39296
rect 9588 39253 9597 39287
rect 9597 39253 9631 39287
rect 9631 39253 9640 39287
rect 9588 39244 9640 39253
rect 11336 39244 11388 39296
rect 13268 39287 13320 39296
rect 13268 39253 13277 39287
rect 13277 39253 13311 39287
rect 13311 39253 13320 39287
rect 13268 39244 13320 39253
rect 15476 39287 15528 39296
rect 15476 39253 15485 39287
rect 15485 39253 15519 39287
rect 15519 39253 15528 39287
rect 15476 39244 15528 39253
rect 15568 39287 15620 39296
rect 15568 39253 15577 39287
rect 15577 39253 15611 39287
rect 15611 39253 15620 39287
rect 15568 39244 15620 39253
rect 16304 39244 16356 39296
rect 18420 39287 18472 39296
rect 18420 39253 18429 39287
rect 18429 39253 18463 39287
rect 18463 39253 18472 39287
rect 18420 39244 18472 39253
rect 18604 39244 18656 39296
rect 20904 39287 20956 39296
rect 20904 39253 20913 39287
rect 20913 39253 20947 39287
rect 20947 39253 20956 39287
rect 20904 39244 20956 39253
rect 22192 39244 22244 39296
rect 22284 39287 22336 39296
rect 22284 39253 22293 39287
rect 22293 39253 22327 39287
rect 22327 39253 22336 39287
rect 22284 39244 22336 39253
rect 25228 39312 25280 39364
rect 24768 39244 24820 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 5356 39083 5408 39092
rect 5356 39049 5365 39083
rect 5365 39049 5399 39083
rect 5399 39049 5408 39083
rect 5356 39040 5408 39049
rect 5908 39040 5960 39092
rect 7380 39040 7432 39092
rect 8760 39083 8812 39092
rect 8760 39049 8769 39083
rect 8769 39049 8803 39083
rect 8803 39049 8812 39083
rect 8760 39040 8812 39049
rect 9404 39040 9456 39092
rect 9588 39040 9640 39092
rect 12440 39040 12492 39092
rect 6000 38947 6052 38956
rect 6000 38913 6009 38947
rect 6009 38913 6043 38947
rect 6043 38913 6052 38947
rect 6000 38904 6052 38913
rect 6092 38904 6144 38956
rect 7012 38879 7064 38888
rect 7012 38845 7021 38879
rect 7021 38845 7055 38879
rect 7055 38845 7064 38879
rect 7012 38836 7064 38845
rect 17868 39040 17920 39092
rect 20352 39083 20404 39092
rect 20352 39049 20361 39083
rect 20361 39049 20395 39083
rect 20395 39049 20404 39083
rect 20352 39040 20404 39049
rect 23296 39040 23348 39092
rect 23664 39040 23716 39092
rect 13820 38972 13872 39024
rect 13912 39015 13964 39024
rect 13912 38981 13921 39015
rect 13921 38981 13955 39015
rect 13955 38981 13964 39015
rect 13912 38972 13964 38981
rect 17316 38972 17368 39024
rect 18604 38972 18656 39024
rect 10324 38904 10376 38956
rect 14188 38947 14240 38956
rect 14188 38913 14197 38947
rect 14197 38913 14231 38947
rect 14231 38913 14240 38947
rect 14188 38904 14240 38913
rect 15660 38904 15712 38956
rect 8576 38879 8628 38888
rect 8576 38845 8585 38879
rect 8585 38845 8619 38879
rect 8619 38845 8628 38879
rect 8576 38836 8628 38845
rect 9956 38879 10008 38888
rect 9956 38845 9965 38879
rect 9965 38845 9999 38879
rect 9999 38845 10008 38879
rect 9956 38836 10008 38845
rect 10048 38836 10100 38888
rect 11704 38879 11756 38888
rect 11704 38845 11713 38879
rect 11713 38845 11747 38879
rect 11747 38845 11756 38879
rect 11704 38836 11756 38845
rect 9036 38768 9088 38820
rect 12348 38768 12400 38820
rect 12624 38768 12676 38820
rect 9680 38700 9732 38752
rect 15844 38836 15896 38888
rect 14188 38768 14240 38820
rect 13268 38700 13320 38752
rect 13452 38700 13504 38752
rect 13820 38700 13872 38752
rect 14556 38700 14608 38752
rect 15384 38768 15436 38820
rect 16304 38700 16356 38752
rect 16672 38700 16724 38752
rect 17684 38700 17736 38752
rect 20996 38972 21048 39024
rect 22468 38972 22520 39024
rect 24584 38972 24636 39024
rect 19708 38904 19760 38956
rect 22192 38904 22244 38956
rect 18880 38768 18932 38820
rect 20168 38879 20220 38888
rect 20168 38845 20177 38879
rect 20177 38845 20211 38879
rect 20211 38845 20220 38879
rect 20168 38836 20220 38845
rect 20720 38836 20772 38888
rect 21824 38836 21876 38888
rect 21548 38768 21600 38820
rect 22560 38836 22612 38888
rect 24308 38904 24360 38956
rect 24032 38836 24084 38888
rect 24768 38836 24820 38888
rect 25872 38768 25924 38820
rect 20720 38700 20772 38752
rect 20812 38743 20864 38752
rect 20812 38709 20821 38743
rect 20821 38709 20855 38743
rect 20855 38709 20864 38743
rect 20812 38700 20864 38709
rect 20996 38700 21048 38752
rect 22008 38743 22060 38752
rect 22008 38709 22017 38743
rect 22017 38709 22051 38743
rect 22051 38709 22060 38743
rect 22008 38700 22060 38709
rect 22468 38700 22520 38752
rect 23572 38700 23624 38752
rect 24308 38700 24360 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 10692 38496 10744 38548
rect 11796 38496 11848 38548
rect 8484 38428 8536 38480
rect 5448 38360 5500 38412
rect 6552 38360 6604 38412
rect 6644 38360 6696 38412
rect 1308 38292 1360 38344
rect 4068 38156 4120 38208
rect 6368 38224 6420 38276
rect 8300 38292 8352 38344
rect 9956 38292 10008 38344
rect 11060 38403 11112 38412
rect 11060 38369 11069 38403
rect 11069 38369 11103 38403
rect 11103 38369 11112 38403
rect 11060 38360 11112 38369
rect 11980 38428 12032 38480
rect 12440 38360 12492 38412
rect 11704 38292 11756 38344
rect 16120 38428 16172 38480
rect 7472 38156 7524 38208
rect 8300 38156 8352 38208
rect 12808 38224 12860 38276
rect 9864 38156 9916 38208
rect 11244 38199 11296 38208
rect 11244 38165 11253 38199
rect 11253 38165 11287 38199
rect 11287 38165 11296 38199
rect 11244 38156 11296 38165
rect 15384 38360 15436 38412
rect 15660 38403 15712 38412
rect 15660 38369 15669 38403
rect 15669 38369 15703 38403
rect 15703 38369 15712 38403
rect 15660 38360 15712 38369
rect 15844 38360 15896 38412
rect 16580 38428 16632 38480
rect 16396 38360 16448 38412
rect 18328 38496 18380 38548
rect 19340 38496 19392 38548
rect 23572 38496 23624 38548
rect 24400 38496 24452 38548
rect 18604 38428 18656 38480
rect 21548 38428 21600 38480
rect 22652 38428 22704 38480
rect 14924 38292 14976 38344
rect 17408 38292 17460 38344
rect 13820 38224 13872 38276
rect 19616 38360 19668 38412
rect 20076 38360 20128 38412
rect 17776 38335 17828 38344
rect 17776 38301 17785 38335
rect 17785 38301 17819 38335
rect 17819 38301 17828 38335
rect 17776 38292 17828 38301
rect 18328 38292 18380 38344
rect 18880 38292 18932 38344
rect 21364 38335 21416 38344
rect 21364 38301 21373 38335
rect 21373 38301 21407 38335
rect 21407 38301 21416 38335
rect 21364 38292 21416 38301
rect 19156 38224 19208 38276
rect 20076 38224 20128 38276
rect 22100 38403 22152 38412
rect 22100 38369 22109 38403
rect 22109 38369 22143 38403
rect 22143 38369 22152 38403
rect 22100 38360 22152 38369
rect 22008 38292 22060 38344
rect 23388 38360 23440 38412
rect 24400 38292 24452 38344
rect 25228 38335 25280 38344
rect 25228 38301 25237 38335
rect 25237 38301 25271 38335
rect 25271 38301 25280 38335
rect 25228 38292 25280 38301
rect 14740 38156 14792 38208
rect 15384 38199 15436 38208
rect 15384 38165 15393 38199
rect 15393 38165 15427 38199
rect 15427 38165 15436 38199
rect 15384 38156 15436 38165
rect 16764 38156 16816 38208
rect 17224 38156 17276 38208
rect 17960 38156 18012 38208
rect 20628 38156 20680 38208
rect 22100 38224 22152 38276
rect 22284 38224 22336 38276
rect 22376 38156 22428 38208
rect 22560 38199 22612 38208
rect 22560 38165 22569 38199
rect 22569 38165 22603 38199
rect 22603 38165 22612 38199
rect 22560 38156 22612 38165
rect 23388 38199 23440 38208
rect 23388 38165 23397 38199
rect 23397 38165 23431 38199
rect 23431 38165 23440 38199
rect 23388 38156 23440 38165
rect 23848 38156 23900 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 5448 37952 5500 38004
rect 6000 37995 6052 38004
rect 6000 37961 6009 37995
rect 6009 37961 6043 37995
rect 6043 37961 6052 37995
rect 6000 37952 6052 37961
rect 8852 37995 8904 38004
rect 6368 37884 6420 37936
rect 8852 37961 8861 37995
rect 8861 37961 8895 37995
rect 8895 37961 8904 37995
rect 8852 37952 8904 37961
rect 10416 37952 10468 38004
rect 10600 37995 10652 38004
rect 10600 37961 10609 37995
rect 10609 37961 10643 37995
rect 10643 37961 10652 37995
rect 10600 37952 10652 37961
rect 8300 37927 8352 37936
rect 8300 37893 8309 37927
rect 8309 37893 8343 37927
rect 8343 37893 8352 37927
rect 8300 37884 8352 37893
rect 8668 37816 8720 37868
rect 14740 37952 14792 38004
rect 15384 37952 15436 38004
rect 16488 37952 16540 38004
rect 16856 37995 16908 38004
rect 16856 37961 16865 37995
rect 16865 37961 16899 37995
rect 16899 37961 16908 37995
rect 16856 37952 16908 37961
rect 14556 37884 14608 37936
rect 5540 37748 5592 37800
rect 7104 37748 7156 37800
rect 8576 37791 8628 37800
rect 8576 37757 8585 37791
rect 8585 37757 8619 37791
rect 8619 37757 8628 37791
rect 8576 37748 8628 37757
rect 9588 37748 9640 37800
rect 15200 37816 15252 37868
rect 15568 37884 15620 37936
rect 19524 37995 19576 38004
rect 19524 37961 19533 37995
rect 19533 37961 19567 37995
rect 19567 37961 19576 37995
rect 19524 37952 19576 37961
rect 20628 37995 20680 38004
rect 20628 37961 20637 37995
rect 20637 37961 20671 37995
rect 20671 37961 20680 37995
rect 20628 37952 20680 37961
rect 18420 37884 18472 37936
rect 18880 37884 18932 37936
rect 21272 37995 21324 38004
rect 21272 37961 21281 37995
rect 21281 37961 21315 37995
rect 21315 37961 21324 37995
rect 21272 37952 21324 37961
rect 15660 37816 15712 37868
rect 16120 37816 16172 37868
rect 16948 37816 17000 37868
rect 11428 37680 11480 37732
rect 14004 37791 14056 37800
rect 14004 37757 14013 37791
rect 14013 37757 14047 37791
rect 14047 37757 14056 37791
rect 14004 37748 14056 37757
rect 14280 37748 14332 37800
rect 15384 37791 15436 37800
rect 15384 37757 15393 37791
rect 15393 37757 15427 37791
rect 15427 37757 15436 37791
rect 15384 37748 15436 37757
rect 20352 37816 20404 37868
rect 21732 37884 21784 37936
rect 22192 37952 22244 38004
rect 22376 37816 22428 37868
rect 17776 37748 17828 37800
rect 16120 37680 16172 37732
rect 19432 37680 19484 37732
rect 8944 37612 8996 37664
rect 11612 37612 11664 37664
rect 13728 37612 13780 37664
rect 17316 37612 17368 37664
rect 21548 37748 21600 37800
rect 22284 37748 22336 37800
rect 23756 37952 23808 38004
rect 24400 37995 24452 38004
rect 24400 37961 24409 37995
rect 24409 37961 24443 37995
rect 24443 37961 24452 37995
rect 24400 37952 24452 37961
rect 23664 37884 23716 37936
rect 24216 37816 24268 37868
rect 24768 37816 24820 37868
rect 22468 37680 22520 37732
rect 23664 37748 23716 37800
rect 21548 37612 21600 37664
rect 25504 37612 25556 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 7656 37408 7708 37460
rect 11060 37408 11112 37460
rect 11980 37408 12032 37460
rect 14464 37451 14516 37460
rect 14464 37417 14473 37451
rect 14473 37417 14507 37451
rect 14507 37417 14516 37451
rect 14464 37408 14516 37417
rect 16120 37451 16172 37460
rect 16120 37417 16129 37451
rect 16129 37417 16163 37451
rect 16163 37417 16172 37451
rect 16120 37408 16172 37417
rect 18880 37408 18932 37460
rect 19064 37408 19116 37460
rect 21272 37408 21324 37460
rect 23664 37408 23716 37460
rect 24124 37408 24176 37460
rect 24216 37451 24268 37460
rect 24216 37417 24225 37451
rect 24225 37417 24259 37451
rect 24259 37417 24268 37451
rect 24216 37408 24268 37417
rect 6552 37340 6604 37392
rect 8576 37340 8628 37392
rect 6000 37272 6052 37324
rect 9220 37315 9272 37324
rect 9220 37281 9229 37315
rect 9229 37281 9263 37315
rect 9263 37281 9272 37315
rect 9220 37272 9272 37281
rect 9312 37272 9364 37324
rect 8944 37204 8996 37256
rect 10600 37204 10652 37256
rect 11336 37272 11388 37324
rect 14372 37340 14424 37392
rect 8668 37136 8720 37188
rect 12624 37204 12676 37256
rect 14004 37204 14056 37256
rect 13636 37136 13688 37188
rect 14832 37272 14884 37324
rect 23296 37340 23348 37392
rect 15936 37272 15988 37324
rect 17224 37272 17276 37324
rect 17868 37272 17920 37324
rect 17316 37204 17368 37256
rect 18788 37204 18840 37256
rect 21272 37204 21324 37256
rect 22100 37204 22152 37256
rect 24032 37204 24084 37256
rect 24124 37204 24176 37256
rect 24400 37204 24452 37256
rect 18604 37136 18656 37188
rect 19340 37136 19392 37188
rect 22284 37179 22336 37188
rect 22284 37145 22293 37179
rect 22293 37145 22327 37179
rect 22327 37145 22336 37179
rect 22284 37136 22336 37145
rect 9128 37068 9180 37120
rect 10232 37068 10284 37120
rect 10876 37111 10928 37120
rect 10876 37077 10885 37111
rect 10885 37077 10919 37111
rect 10919 37077 10928 37111
rect 10876 37068 10928 37077
rect 11980 37068 12032 37120
rect 13820 37068 13872 37120
rect 14740 37111 14792 37120
rect 14740 37077 14749 37111
rect 14749 37077 14783 37111
rect 14783 37077 14792 37111
rect 14740 37068 14792 37077
rect 15292 37068 15344 37120
rect 15936 37068 15988 37120
rect 16580 37111 16632 37120
rect 16580 37077 16589 37111
rect 16589 37077 16623 37111
rect 16623 37077 16632 37111
rect 16580 37068 16632 37077
rect 17224 37068 17276 37120
rect 17408 37068 17460 37120
rect 18880 37068 18932 37120
rect 19616 37068 19668 37120
rect 20628 37068 20680 37120
rect 25964 37136 26016 37188
rect 22652 37068 22704 37120
rect 25044 37068 25096 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 7472 36907 7524 36916
rect 7472 36873 7481 36907
rect 7481 36873 7515 36907
rect 7515 36873 7524 36907
rect 7472 36864 7524 36873
rect 10048 36864 10100 36916
rect 10600 36864 10652 36916
rect 6368 36796 6420 36848
rect 7656 36796 7708 36848
rect 9036 36796 9088 36848
rect 15292 36864 15344 36916
rect 15936 36907 15988 36916
rect 15936 36873 15945 36907
rect 15945 36873 15979 36907
rect 15979 36873 15988 36907
rect 15936 36864 15988 36873
rect 16396 36907 16448 36916
rect 16396 36873 16405 36907
rect 16405 36873 16439 36907
rect 16439 36873 16448 36907
rect 16396 36864 16448 36873
rect 17224 36907 17276 36916
rect 17224 36873 17233 36907
rect 17233 36873 17267 36907
rect 17267 36873 17276 36907
rect 17224 36864 17276 36873
rect 19708 36864 19760 36916
rect 20168 36864 20220 36916
rect 21364 36864 21416 36916
rect 21640 36864 21692 36916
rect 22192 36864 22244 36916
rect 12624 36796 12676 36848
rect 13728 36796 13780 36848
rect 15108 36839 15160 36848
rect 15108 36805 15117 36839
rect 15117 36805 15151 36839
rect 15151 36805 15160 36839
rect 15108 36796 15160 36805
rect 9220 36771 9272 36780
rect 9220 36737 9229 36771
rect 9229 36737 9263 36771
rect 9263 36737 9272 36771
rect 9220 36728 9272 36737
rect 9404 36728 9456 36780
rect 10324 36703 10376 36712
rect 10324 36669 10333 36703
rect 10333 36669 10367 36703
rect 10367 36669 10376 36703
rect 10324 36660 10376 36669
rect 12716 36592 12768 36644
rect 15936 36728 15988 36780
rect 13728 36660 13780 36712
rect 17500 36660 17552 36712
rect 19616 36796 19668 36848
rect 20536 36796 20588 36848
rect 19984 36728 20036 36780
rect 18972 36635 19024 36644
rect 18972 36601 18981 36635
rect 18981 36601 19015 36635
rect 19015 36601 19024 36635
rect 18972 36592 19024 36601
rect 19524 36703 19576 36712
rect 19524 36669 19533 36703
rect 19533 36669 19567 36703
rect 19567 36669 19576 36703
rect 19524 36660 19576 36669
rect 20444 36660 20496 36712
rect 22468 36796 22520 36848
rect 23388 36864 23440 36916
rect 24676 36864 24728 36916
rect 23664 36796 23716 36848
rect 20996 36592 21048 36644
rect 21364 36592 21416 36644
rect 22192 36592 22244 36644
rect 6828 36524 6880 36576
rect 12164 36567 12216 36576
rect 12164 36533 12173 36567
rect 12173 36533 12207 36567
rect 12207 36533 12216 36567
rect 12164 36524 12216 36533
rect 12256 36567 12308 36576
rect 12256 36533 12265 36567
rect 12265 36533 12299 36567
rect 12299 36533 12308 36567
rect 12256 36524 12308 36533
rect 12348 36524 12400 36576
rect 14372 36524 14424 36576
rect 15936 36524 15988 36576
rect 19524 36524 19576 36576
rect 25044 36839 25096 36848
rect 25044 36805 25053 36839
rect 25053 36805 25087 36839
rect 25087 36805 25096 36839
rect 25044 36796 25096 36805
rect 25044 36660 25096 36712
rect 23388 36524 23440 36576
rect 24860 36524 24912 36576
rect 24952 36524 25004 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 7012 36320 7064 36372
rect 13360 36320 13412 36372
rect 15476 36320 15528 36372
rect 16580 36320 16632 36372
rect 17776 36320 17828 36372
rect 17316 36252 17368 36304
rect 5540 36184 5592 36236
rect 12532 36227 12584 36236
rect 12532 36193 12541 36227
rect 12541 36193 12575 36227
rect 12575 36193 12584 36227
rect 12532 36184 12584 36193
rect 14924 36184 14976 36236
rect 19800 36184 19852 36236
rect 21180 36252 21232 36304
rect 20904 36184 20956 36236
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 6552 36116 6604 36168
rect 11060 36116 11112 36168
rect 11704 36116 11756 36168
rect 12072 36116 12124 36168
rect 12164 36116 12216 36168
rect 15384 36116 15436 36168
rect 6920 36091 6972 36100
rect 6920 36057 6929 36091
rect 6929 36057 6963 36091
rect 6963 36057 6972 36091
rect 6920 36048 6972 36057
rect 7656 36048 7708 36100
rect 14280 36048 14332 36100
rect 16856 36116 16908 36168
rect 21088 36116 21140 36168
rect 25044 36320 25096 36372
rect 24676 36252 24728 36304
rect 22284 36227 22336 36236
rect 22284 36193 22293 36227
rect 22293 36193 22327 36227
rect 22327 36193 22336 36227
rect 22284 36184 22336 36193
rect 24952 36184 25004 36236
rect 23848 36116 23900 36168
rect 22652 36048 22704 36100
rect 23572 36048 23624 36100
rect 23940 36048 23992 36100
rect 4160 35980 4212 36032
rect 11796 35980 11848 36032
rect 12256 35980 12308 36032
rect 12716 36023 12768 36032
rect 12716 35989 12725 36023
rect 12725 35989 12759 36023
rect 12759 35989 12768 36023
rect 12716 35980 12768 35989
rect 12900 35980 12952 36032
rect 15200 35980 15252 36032
rect 15384 35980 15436 36032
rect 18420 35980 18472 36032
rect 19616 35980 19668 36032
rect 20904 35980 20956 36032
rect 24492 35980 24544 36032
rect 24584 36023 24636 36032
rect 24584 35989 24593 36023
rect 24593 35989 24627 36023
rect 24627 35989 24636 36023
rect 24584 35980 24636 35989
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 6552 35776 6604 35828
rect 6920 35776 6972 35828
rect 5908 35708 5960 35760
rect 8300 35708 8352 35760
rect 10324 35776 10376 35828
rect 11704 35819 11756 35828
rect 11704 35785 11713 35819
rect 11713 35785 11747 35819
rect 11747 35785 11756 35819
rect 11704 35776 11756 35785
rect 9772 35708 9824 35760
rect 13912 35776 13964 35828
rect 13452 35708 13504 35760
rect 17500 35708 17552 35760
rect 4528 35615 4580 35624
rect 4528 35581 4537 35615
rect 4537 35581 4571 35615
rect 4571 35581 4580 35615
rect 4528 35572 4580 35581
rect 6000 35615 6052 35624
rect 6000 35581 6009 35615
rect 6009 35581 6043 35615
rect 6043 35581 6052 35615
rect 6000 35572 6052 35581
rect 7012 35479 7064 35488
rect 7012 35445 7021 35479
rect 7021 35445 7055 35479
rect 7055 35445 7064 35479
rect 7012 35436 7064 35445
rect 10692 35640 10744 35692
rect 12072 35640 12124 35692
rect 17224 35640 17276 35692
rect 19432 35776 19484 35828
rect 23664 35776 23716 35828
rect 18420 35708 18472 35760
rect 24400 35708 24452 35760
rect 19248 35640 19300 35692
rect 8760 35615 8812 35624
rect 8760 35581 8769 35615
rect 8769 35581 8803 35615
rect 8803 35581 8812 35615
rect 8760 35572 8812 35581
rect 8852 35572 8904 35624
rect 12532 35572 12584 35624
rect 13452 35615 13504 35624
rect 13452 35581 13461 35615
rect 13461 35581 13495 35615
rect 13495 35581 13504 35615
rect 13452 35572 13504 35581
rect 17776 35572 17828 35624
rect 22652 35615 22704 35624
rect 22652 35581 22661 35615
rect 22661 35581 22695 35615
rect 22695 35581 22704 35615
rect 22652 35572 22704 35581
rect 24032 35572 24084 35624
rect 24676 35615 24728 35624
rect 24676 35581 24685 35615
rect 24685 35581 24719 35615
rect 24719 35581 24728 35615
rect 24676 35572 24728 35581
rect 24952 35615 25004 35624
rect 24952 35581 24961 35615
rect 24961 35581 24995 35615
rect 24995 35581 25004 35615
rect 24952 35572 25004 35581
rect 25136 35572 25188 35624
rect 25596 35572 25648 35624
rect 12440 35436 12492 35488
rect 13360 35436 13412 35488
rect 16304 35436 16356 35488
rect 18328 35436 18380 35488
rect 22008 35436 22060 35488
rect 22468 35436 22520 35488
rect 25320 35436 25372 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 4528 35232 4580 35284
rect 7748 35232 7800 35284
rect 8300 35232 8352 35284
rect 8944 35275 8996 35284
rect 8944 35241 8953 35275
rect 8953 35241 8987 35275
rect 8987 35241 8996 35275
rect 8944 35232 8996 35241
rect 9496 35232 9548 35284
rect 9588 35164 9640 35216
rect 6552 35096 6604 35148
rect 7564 35096 7616 35148
rect 12624 35232 12676 35284
rect 13360 35232 13412 35284
rect 15660 35232 15712 35284
rect 17500 35232 17552 35284
rect 19156 35232 19208 35284
rect 19248 35232 19300 35284
rect 23940 35275 23992 35284
rect 23940 35241 23949 35275
rect 23949 35241 23983 35275
rect 23983 35241 23992 35275
rect 23940 35232 23992 35241
rect 24676 35232 24728 35284
rect 10048 35096 10100 35148
rect 10324 35096 10376 35148
rect 13452 35096 13504 35148
rect 15660 35096 15712 35148
rect 17224 35139 17276 35148
rect 17224 35105 17233 35139
rect 17233 35105 17267 35139
rect 17267 35105 17276 35139
rect 17224 35096 17276 35105
rect 5908 35028 5960 35080
rect 10784 35028 10836 35080
rect 18420 35096 18472 35148
rect 20260 35096 20312 35148
rect 7012 35003 7064 35012
rect 7012 34969 7021 35003
rect 7021 34969 7055 35003
rect 7055 34969 7064 35003
rect 7012 34960 7064 34969
rect 8944 34960 8996 35012
rect 10692 34960 10744 35012
rect 11796 34960 11848 35012
rect 13452 34960 13504 35012
rect 19340 35028 19392 35080
rect 23572 35164 23624 35216
rect 22192 35139 22244 35148
rect 22192 35105 22201 35139
rect 22201 35105 22235 35139
rect 22235 35105 22244 35139
rect 22192 35096 22244 35105
rect 24124 35096 24176 35148
rect 20996 35028 21048 35080
rect 22652 35028 22704 35080
rect 24032 35028 24084 35080
rect 24492 35028 24544 35080
rect 8300 34892 8352 34944
rect 9680 34935 9732 34944
rect 9680 34901 9689 34935
rect 9689 34901 9723 34935
rect 9723 34901 9732 34935
rect 9680 34892 9732 34901
rect 11704 34892 11756 34944
rect 12716 34935 12768 34944
rect 12716 34901 12725 34935
rect 12725 34901 12759 34935
rect 12759 34901 12768 34935
rect 12716 34892 12768 34901
rect 17224 34960 17276 35012
rect 21088 34960 21140 35012
rect 19248 34892 19300 34944
rect 21180 34935 21232 34944
rect 21180 34901 21189 34935
rect 21189 34901 21223 34935
rect 21223 34901 21232 34935
rect 21180 34892 21232 34901
rect 22652 34892 22704 34944
rect 22744 34935 22796 34944
rect 22744 34901 22753 34935
rect 22753 34901 22787 34935
rect 22787 34901 22796 34935
rect 22744 34892 22796 34901
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 4896 34731 4948 34740
rect 4896 34697 4905 34731
rect 4905 34697 4939 34731
rect 4939 34697 4948 34731
rect 4896 34688 4948 34697
rect 6092 34688 6144 34740
rect 7656 34688 7708 34740
rect 6736 34620 6788 34672
rect 5632 34595 5684 34604
rect 5632 34561 5641 34595
rect 5641 34561 5675 34595
rect 5675 34561 5684 34595
rect 5632 34552 5684 34561
rect 8576 34688 8628 34740
rect 9312 34688 9364 34740
rect 11060 34688 11112 34740
rect 11152 34688 11204 34740
rect 11428 34688 11480 34740
rect 12072 34688 12124 34740
rect 10324 34620 10376 34672
rect 11520 34620 11572 34672
rect 11980 34663 12032 34672
rect 11980 34629 11989 34663
rect 11989 34629 12023 34663
rect 12023 34629 12032 34663
rect 11980 34620 12032 34629
rect 12716 34688 12768 34740
rect 13636 34688 13688 34740
rect 14740 34688 14792 34740
rect 17224 34731 17276 34740
rect 17224 34697 17233 34731
rect 17233 34697 17267 34731
rect 17267 34697 17276 34731
rect 17224 34688 17276 34697
rect 17040 34620 17092 34672
rect 18604 34688 18656 34740
rect 21824 34663 21876 34672
rect 21824 34629 21833 34663
rect 21833 34629 21867 34663
rect 21867 34629 21876 34663
rect 21824 34620 21876 34629
rect 22560 34688 22612 34740
rect 22652 34688 22704 34740
rect 22836 34688 22888 34740
rect 24400 34688 24452 34740
rect 24768 34688 24820 34740
rect 5816 34484 5868 34536
rect 6552 34527 6604 34536
rect 6552 34493 6561 34527
rect 6561 34493 6595 34527
rect 6595 34493 6604 34527
rect 6552 34484 6604 34493
rect 6828 34527 6880 34536
rect 6828 34493 6837 34527
rect 6837 34493 6871 34527
rect 6871 34493 6880 34527
rect 6828 34484 6880 34493
rect 8852 34484 8904 34536
rect 9772 34484 9824 34536
rect 5540 34416 5592 34468
rect 11152 34527 11204 34536
rect 11152 34493 11161 34527
rect 11161 34493 11195 34527
rect 11195 34493 11204 34527
rect 11152 34484 11204 34493
rect 12348 34484 12400 34536
rect 12532 34484 12584 34536
rect 13636 34552 13688 34604
rect 13452 34527 13504 34536
rect 13452 34493 13461 34527
rect 13461 34493 13495 34527
rect 13495 34493 13504 34527
rect 13452 34484 13504 34493
rect 11060 34416 11112 34468
rect 18328 34552 18380 34604
rect 17776 34484 17828 34536
rect 19432 34552 19484 34604
rect 20260 34595 20312 34604
rect 20260 34561 20269 34595
rect 20269 34561 20303 34595
rect 20303 34561 20312 34595
rect 20260 34552 20312 34561
rect 20812 34552 20864 34604
rect 22376 34552 22428 34604
rect 24216 34552 24268 34604
rect 24308 34552 24360 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 18604 34416 18656 34468
rect 18696 34416 18748 34468
rect 20720 34484 20772 34536
rect 22100 34416 22152 34468
rect 23664 34484 23716 34536
rect 24032 34348 24084 34400
rect 25136 34391 25188 34400
rect 25136 34357 25145 34391
rect 25145 34357 25179 34391
rect 25179 34357 25188 34391
rect 25136 34348 25188 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 6828 34144 6880 34196
rect 8760 34144 8812 34196
rect 9128 34187 9180 34196
rect 9128 34153 9137 34187
rect 9137 34153 9171 34187
rect 9171 34153 9180 34187
rect 9128 34144 9180 34153
rect 9772 34144 9824 34196
rect 11244 34144 11296 34196
rect 11520 34144 11572 34196
rect 14188 34144 14240 34196
rect 14280 34187 14332 34196
rect 14280 34153 14289 34187
rect 14289 34153 14323 34187
rect 14323 34153 14332 34187
rect 14280 34144 14332 34153
rect 18420 34144 18472 34196
rect 21088 34144 21140 34196
rect 21364 34144 21416 34196
rect 5632 34008 5684 34060
rect 9588 34008 9640 34060
rect 11520 34051 11572 34060
rect 11520 34017 11529 34051
rect 11529 34017 11563 34051
rect 11563 34017 11572 34051
rect 11520 34008 11572 34017
rect 11888 34076 11940 34128
rect 12440 34076 12492 34128
rect 11704 34008 11756 34060
rect 16856 34076 16908 34128
rect 19708 34076 19760 34128
rect 6000 33940 6052 33992
rect 8576 33983 8628 33992
rect 8576 33949 8585 33983
rect 8585 33949 8619 33983
rect 8619 33949 8628 33983
rect 8576 33940 8628 33949
rect 11152 33940 11204 33992
rect 11244 33940 11296 33992
rect 15568 33983 15620 33992
rect 15568 33949 15577 33983
rect 15577 33949 15611 33983
rect 15611 33949 15620 33983
rect 15568 33940 15620 33949
rect 16856 33940 16908 33992
rect 19248 34008 19300 34060
rect 22468 34076 22520 34128
rect 12164 33872 12216 33924
rect 13544 33872 13596 33924
rect 15108 33872 15160 33924
rect 7840 33804 7892 33856
rect 11428 33847 11480 33856
rect 11428 33813 11437 33847
rect 11437 33813 11471 33847
rect 11471 33813 11480 33847
rect 11428 33804 11480 33813
rect 12716 33804 12768 33856
rect 13360 33847 13412 33856
rect 13360 33813 13369 33847
rect 13369 33813 13403 33847
rect 13403 33813 13412 33847
rect 13360 33804 13412 33813
rect 14096 33804 14148 33856
rect 20996 33940 21048 33992
rect 21364 34008 21416 34060
rect 21456 34051 21508 34060
rect 21456 34017 21465 34051
rect 21465 34017 21499 34051
rect 21499 34017 21508 34051
rect 21456 34008 21508 34017
rect 21824 33940 21876 33992
rect 22008 33983 22060 33992
rect 22008 33949 22017 33983
rect 22017 33949 22051 33983
rect 22051 33949 22060 33983
rect 22008 33940 22060 33949
rect 24860 34144 24912 34196
rect 25412 33940 25464 33992
rect 17776 33804 17828 33856
rect 21732 33872 21784 33924
rect 22468 33872 22520 33924
rect 19892 33847 19944 33856
rect 19892 33813 19901 33847
rect 19901 33813 19935 33847
rect 19935 33813 19944 33847
rect 19892 33804 19944 33813
rect 20720 33804 20772 33856
rect 20812 33847 20864 33856
rect 20812 33813 20821 33847
rect 20821 33813 20855 33847
rect 20855 33813 20864 33847
rect 20812 33804 20864 33813
rect 22652 33847 22704 33856
rect 22652 33813 22661 33847
rect 22661 33813 22695 33847
rect 22695 33813 22704 33847
rect 22652 33804 22704 33813
rect 23112 33847 23164 33856
rect 23112 33813 23121 33847
rect 23121 33813 23155 33847
rect 23155 33813 23164 33847
rect 23112 33804 23164 33813
rect 23204 33804 23256 33856
rect 23480 33804 23532 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 6184 33600 6236 33652
rect 7656 33643 7708 33652
rect 7656 33609 7665 33643
rect 7665 33609 7699 33643
rect 7699 33609 7708 33643
rect 7656 33600 7708 33609
rect 9680 33600 9732 33652
rect 10876 33600 10928 33652
rect 10784 33532 10836 33584
rect 12256 33600 12308 33652
rect 15108 33643 15160 33652
rect 15108 33609 15117 33643
rect 15117 33609 15151 33643
rect 15151 33609 15160 33643
rect 15108 33600 15160 33609
rect 17408 33600 17460 33652
rect 19616 33600 19668 33652
rect 19708 33600 19760 33652
rect 19248 33532 19300 33584
rect 23112 33600 23164 33652
rect 25228 33643 25280 33652
rect 25228 33609 25237 33643
rect 25237 33609 25271 33643
rect 25271 33609 25280 33643
rect 25228 33600 25280 33609
rect 23848 33532 23900 33584
rect 24492 33532 24544 33584
rect 1216 33464 1268 33516
rect 8392 33507 8444 33516
rect 8392 33473 8401 33507
rect 8401 33473 8435 33507
rect 8435 33473 8444 33507
rect 8392 33464 8444 33473
rect 11428 33464 11480 33516
rect 11796 33464 11848 33516
rect 14280 33464 14332 33516
rect 14464 33507 14516 33516
rect 14464 33473 14473 33507
rect 14473 33473 14507 33507
rect 14507 33473 14516 33507
rect 14464 33464 14516 33473
rect 16948 33464 17000 33516
rect 21180 33464 21232 33516
rect 9036 33396 9088 33448
rect 7104 33328 7156 33380
rect 9956 33396 10008 33448
rect 3884 33260 3936 33312
rect 9036 33303 9088 33312
rect 9036 33269 9045 33303
rect 9045 33269 9079 33303
rect 9079 33269 9088 33303
rect 9036 33260 9088 33269
rect 11060 33328 11112 33380
rect 12348 33396 12400 33448
rect 15200 33396 15252 33448
rect 16120 33439 16172 33448
rect 16120 33405 16129 33439
rect 16129 33405 16163 33439
rect 16163 33405 16172 33439
rect 16120 33396 16172 33405
rect 19432 33396 19484 33448
rect 20352 33396 20404 33448
rect 22468 33439 22520 33448
rect 22468 33405 22477 33439
rect 22477 33405 22511 33439
rect 22511 33405 22520 33439
rect 22468 33396 22520 33405
rect 23296 33396 23348 33448
rect 13360 33328 13412 33380
rect 17684 33328 17736 33380
rect 21824 33328 21876 33380
rect 23204 33328 23256 33380
rect 14096 33303 14148 33312
rect 14096 33269 14105 33303
rect 14105 33269 14139 33303
rect 14139 33269 14148 33303
rect 14096 33260 14148 33269
rect 15568 33303 15620 33312
rect 15568 33269 15577 33303
rect 15577 33269 15611 33303
rect 15611 33269 15620 33303
rect 15568 33260 15620 33269
rect 15936 33260 15988 33312
rect 16396 33260 16448 33312
rect 18328 33260 18380 33312
rect 18972 33260 19024 33312
rect 20720 33260 20772 33312
rect 22284 33260 22336 33312
rect 22560 33260 22612 33312
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 23756 33396 23808 33405
rect 24952 33260 25004 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 7564 33099 7616 33108
rect 7564 33065 7573 33099
rect 7573 33065 7607 33099
rect 7607 33065 7616 33099
rect 7564 33056 7616 33065
rect 7104 32920 7156 32972
rect 8944 33056 8996 33108
rect 9680 33056 9732 33108
rect 16212 33056 16264 33108
rect 5816 32895 5868 32904
rect 5816 32861 5825 32895
rect 5825 32861 5859 32895
rect 5859 32861 5868 32895
rect 5816 32852 5868 32861
rect 8392 32963 8444 32972
rect 8392 32929 8401 32963
rect 8401 32929 8435 32963
rect 8435 32929 8444 32963
rect 8392 32920 8444 32929
rect 15660 32920 15712 32972
rect 7564 32852 7616 32904
rect 16672 32852 16724 32904
rect 10968 32784 11020 32836
rect 12808 32784 12860 32836
rect 8300 32716 8352 32768
rect 14188 32716 14240 32768
rect 14832 32716 14884 32768
rect 15108 32716 15160 32768
rect 15660 32784 15712 32836
rect 17224 33056 17276 33108
rect 17684 33056 17736 33108
rect 18512 33056 18564 33108
rect 18880 33056 18932 33108
rect 23480 33099 23532 33108
rect 23480 33065 23489 33099
rect 23489 33065 23523 33099
rect 23523 33065 23532 33099
rect 23480 33056 23532 33065
rect 23848 33099 23900 33108
rect 23848 33065 23857 33099
rect 23857 33065 23891 33099
rect 23891 33065 23900 33099
rect 23848 33056 23900 33065
rect 25044 33056 25096 33108
rect 17408 32988 17460 33040
rect 19892 32988 19944 33040
rect 17500 32920 17552 32972
rect 19616 32920 19668 32972
rect 20260 32920 20312 32972
rect 17592 32852 17644 32904
rect 20352 32784 20404 32836
rect 22100 32988 22152 33040
rect 22284 32988 22336 33040
rect 21088 32920 21140 32972
rect 22008 32920 22060 32972
rect 21732 32852 21784 32904
rect 22376 32895 22428 32904
rect 22376 32861 22385 32895
rect 22385 32861 22419 32895
rect 22419 32861 22428 32895
rect 22376 32852 22428 32861
rect 22836 32852 22888 32904
rect 21824 32784 21876 32836
rect 16580 32716 16632 32768
rect 17224 32716 17276 32768
rect 17500 32759 17552 32768
rect 17500 32725 17509 32759
rect 17509 32725 17543 32759
rect 17543 32725 17552 32759
rect 17500 32716 17552 32725
rect 19340 32716 19392 32768
rect 19800 32716 19852 32768
rect 22376 32716 22428 32768
rect 24124 32784 24176 32836
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 24952 32784 25004 32836
rect 24676 32759 24728 32768
rect 24676 32725 24685 32759
rect 24685 32725 24719 32759
rect 24719 32725 24728 32759
rect 24676 32716 24728 32725
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 12808 32512 12860 32564
rect 15660 32512 15712 32564
rect 17316 32512 17368 32564
rect 17500 32512 17552 32564
rect 18788 32512 18840 32564
rect 8300 32487 8352 32496
rect 8300 32453 8309 32487
rect 8309 32453 8343 32487
rect 8343 32453 8352 32487
rect 8300 32444 8352 32453
rect 9680 32444 9732 32496
rect 10600 32444 10652 32496
rect 14188 32444 14240 32496
rect 14372 32487 14424 32496
rect 14372 32453 14381 32487
rect 14381 32453 14415 32487
rect 14415 32453 14424 32487
rect 14372 32444 14424 32453
rect 14648 32444 14700 32496
rect 17776 32444 17828 32496
rect 19524 32444 19576 32496
rect 5816 32376 5868 32428
rect 12808 32376 12860 32428
rect 7748 32308 7800 32360
rect 8024 32351 8076 32360
rect 8024 32317 8033 32351
rect 8033 32317 8067 32351
rect 8067 32317 8076 32351
rect 8024 32308 8076 32317
rect 9036 32308 9088 32360
rect 11704 32308 11756 32360
rect 13728 32376 13780 32428
rect 16120 32376 16172 32428
rect 16948 32376 17000 32428
rect 17408 32376 17460 32428
rect 19156 32419 19208 32428
rect 19156 32385 19165 32419
rect 19165 32385 19199 32419
rect 19199 32385 19208 32419
rect 19156 32376 19208 32385
rect 19800 32376 19852 32428
rect 20628 32512 20680 32564
rect 20352 32487 20404 32496
rect 20352 32453 20361 32487
rect 20361 32453 20395 32487
rect 20395 32453 20404 32487
rect 20352 32444 20404 32453
rect 21548 32444 21600 32496
rect 22192 32512 22244 32564
rect 22376 32512 22428 32564
rect 22468 32555 22520 32564
rect 22468 32521 22477 32555
rect 22477 32521 22511 32555
rect 22511 32521 22520 32555
rect 22468 32512 22520 32521
rect 23756 32512 23808 32564
rect 23572 32444 23624 32496
rect 13452 32308 13504 32360
rect 17132 32308 17184 32360
rect 19340 32308 19392 32360
rect 9588 32240 9640 32292
rect 15108 32240 15160 32292
rect 16856 32240 16908 32292
rect 17500 32240 17552 32292
rect 18880 32240 18932 32292
rect 20536 32351 20588 32360
rect 20536 32317 20545 32351
rect 20545 32317 20579 32351
rect 20579 32317 20588 32351
rect 20536 32308 20588 32317
rect 21548 32308 21600 32360
rect 21916 32308 21968 32360
rect 19800 32240 19852 32292
rect 6920 32172 6972 32224
rect 7104 32172 7156 32224
rect 7288 32172 7340 32224
rect 10968 32172 11020 32224
rect 14832 32215 14884 32224
rect 14832 32181 14841 32215
rect 14841 32181 14875 32215
rect 14875 32181 14884 32215
rect 14832 32172 14884 32181
rect 14924 32172 14976 32224
rect 17592 32215 17644 32224
rect 17592 32181 17601 32215
rect 17601 32181 17635 32215
rect 17635 32181 17644 32215
rect 17592 32172 17644 32181
rect 19156 32172 19208 32224
rect 19340 32172 19392 32224
rect 22192 32351 22244 32360
rect 22192 32317 22201 32351
rect 22201 32317 22235 32351
rect 22235 32317 22244 32351
rect 22192 32308 22244 32317
rect 22376 32351 22428 32360
rect 22376 32317 22385 32351
rect 22385 32317 22419 32351
rect 22419 32317 22428 32351
rect 22376 32308 22428 32317
rect 23480 32419 23532 32428
rect 23480 32385 23489 32419
rect 23489 32385 23523 32419
rect 23523 32385 23532 32419
rect 23480 32376 23532 32385
rect 24216 32376 24268 32428
rect 24676 32419 24728 32428
rect 24676 32385 24685 32419
rect 24685 32385 24719 32419
rect 24719 32385 24728 32419
rect 24676 32376 24728 32385
rect 25136 32308 25188 32360
rect 25228 32351 25280 32360
rect 25228 32317 25237 32351
rect 25237 32317 25271 32351
rect 25271 32317 25280 32351
rect 25228 32308 25280 32317
rect 25596 32308 25648 32360
rect 24032 32240 24084 32292
rect 22836 32215 22888 32224
rect 22836 32181 22845 32215
rect 22845 32181 22879 32215
rect 22879 32181 22888 32215
rect 22836 32172 22888 32181
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 6920 31968 6972 32020
rect 9680 31968 9732 32020
rect 11152 31968 11204 32020
rect 11704 31968 11756 32020
rect 12624 31968 12676 32020
rect 15660 31968 15712 32020
rect 8024 31832 8076 31884
rect 8852 31832 8904 31884
rect 10232 31832 10284 31884
rect 11428 31832 11480 31884
rect 11704 31832 11756 31884
rect 12072 31832 12124 31884
rect 12348 31832 12400 31884
rect 12808 31875 12860 31884
rect 12808 31841 12817 31875
rect 12817 31841 12851 31875
rect 12851 31841 12860 31875
rect 12808 31832 12860 31841
rect 9588 31764 9640 31816
rect 13360 31764 13412 31816
rect 18328 31968 18380 32020
rect 19616 31968 19668 32020
rect 19800 32011 19852 32020
rect 19800 31977 19809 32011
rect 19809 31977 19843 32011
rect 19843 31977 19852 32011
rect 19800 31968 19852 31977
rect 20628 32011 20680 32020
rect 20628 31977 20637 32011
rect 20637 31977 20671 32011
rect 20671 31977 20680 32011
rect 20628 31968 20680 31977
rect 22376 31968 22428 32020
rect 22652 31968 22704 32020
rect 24032 32011 24084 32020
rect 24032 31977 24041 32011
rect 24041 31977 24075 32011
rect 24075 31977 24084 32011
rect 24032 31968 24084 31977
rect 17408 31900 17460 31952
rect 18420 31900 18472 31952
rect 19524 31900 19576 31952
rect 20536 31900 20588 31952
rect 21916 31943 21968 31952
rect 21916 31909 21925 31943
rect 21925 31909 21959 31943
rect 21959 31909 21968 31943
rect 21916 31900 21968 31909
rect 19432 31832 19484 31884
rect 21088 31875 21140 31884
rect 21088 31841 21097 31875
rect 21097 31841 21131 31875
rect 21131 31841 21140 31875
rect 21088 31832 21140 31841
rect 21180 31875 21232 31884
rect 21180 31841 21189 31875
rect 21189 31841 21223 31875
rect 21223 31841 21232 31875
rect 21180 31832 21232 31841
rect 23296 31832 23348 31884
rect 10692 31696 10744 31748
rect 9128 31671 9180 31680
rect 9128 31637 9137 31671
rect 9137 31637 9171 31671
rect 9171 31637 9180 31671
rect 9128 31628 9180 31637
rect 13728 31696 13780 31748
rect 15660 31696 15712 31748
rect 16672 31696 16724 31748
rect 17684 31807 17736 31816
rect 17684 31773 17693 31807
rect 17693 31773 17727 31807
rect 17727 31773 17736 31807
rect 17684 31764 17736 31773
rect 18880 31696 18932 31748
rect 19248 31696 19300 31748
rect 24492 31696 24544 31748
rect 14004 31628 14056 31680
rect 14648 31671 14700 31680
rect 14648 31637 14657 31671
rect 14657 31637 14691 31671
rect 14691 31637 14700 31671
rect 14648 31628 14700 31637
rect 15108 31628 15160 31680
rect 15936 31628 15988 31680
rect 16580 31628 16632 31680
rect 17500 31628 17552 31680
rect 17776 31628 17828 31680
rect 20352 31628 20404 31680
rect 21364 31628 21416 31680
rect 21640 31628 21692 31680
rect 22100 31628 22152 31680
rect 23848 31628 23900 31680
rect 24952 31628 25004 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 9128 31424 9180 31476
rect 15660 31424 15712 31476
rect 13912 31356 13964 31408
rect 16028 31399 16080 31408
rect 16028 31365 16037 31399
rect 16037 31365 16071 31399
rect 16071 31365 16080 31399
rect 16028 31356 16080 31365
rect 16304 31467 16356 31476
rect 16304 31433 16313 31467
rect 16313 31433 16347 31467
rect 16347 31433 16356 31467
rect 16304 31424 16356 31433
rect 16948 31424 17000 31476
rect 18604 31424 18656 31476
rect 18696 31424 18748 31476
rect 20720 31424 20772 31476
rect 20996 31424 21048 31476
rect 21180 31467 21232 31476
rect 21180 31433 21189 31467
rect 21189 31433 21223 31467
rect 21223 31433 21232 31467
rect 21180 31424 21232 31433
rect 23296 31424 23348 31476
rect 3700 31288 3752 31340
rect 11336 31288 11388 31340
rect 12348 31288 12400 31340
rect 3976 31263 4028 31272
rect 3976 31229 3985 31263
rect 3985 31229 4019 31263
rect 4019 31229 4028 31263
rect 3976 31220 4028 31229
rect 4896 31263 4948 31272
rect 4896 31229 4905 31263
rect 4905 31229 4939 31263
rect 4939 31229 4948 31263
rect 4896 31220 4948 31229
rect 7012 31220 7064 31272
rect 7656 31263 7708 31272
rect 7656 31229 7665 31263
rect 7665 31229 7699 31263
rect 7699 31229 7708 31263
rect 7656 31220 7708 31229
rect 5264 31152 5316 31204
rect 8300 31220 8352 31272
rect 14924 31220 14976 31272
rect 7840 31152 7892 31204
rect 11244 31084 11296 31136
rect 12072 31084 12124 31136
rect 17224 31331 17276 31340
rect 17224 31297 17233 31331
rect 17233 31297 17267 31331
rect 17267 31297 17276 31331
rect 17224 31288 17276 31297
rect 15476 31263 15528 31272
rect 15476 31229 15485 31263
rect 15485 31229 15519 31263
rect 15519 31229 15528 31263
rect 15476 31220 15528 31229
rect 20904 31356 20956 31408
rect 23388 31356 23440 31408
rect 24492 31356 24544 31408
rect 24952 31399 25004 31408
rect 24952 31365 24961 31399
rect 24961 31365 24995 31399
rect 24995 31365 25004 31399
rect 24952 31356 25004 31365
rect 18696 31331 18748 31340
rect 18696 31297 18705 31331
rect 18705 31297 18739 31331
rect 18739 31297 18748 31331
rect 18696 31288 18748 31297
rect 16304 31152 16356 31204
rect 16672 31152 16724 31204
rect 17776 31152 17828 31204
rect 14096 31084 14148 31136
rect 14464 31084 14516 31136
rect 14648 31084 14700 31136
rect 15936 31084 15988 31136
rect 18972 31220 19024 31272
rect 21272 31263 21324 31272
rect 21272 31229 21281 31263
rect 21281 31229 21315 31263
rect 21315 31229 21324 31263
rect 21272 31220 21324 31229
rect 22100 31263 22152 31272
rect 22100 31229 22109 31263
rect 22109 31229 22143 31263
rect 22143 31229 22152 31263
rect 22100 31220 22152 31229
rect 23480 31263 23532 31272
rect 23480 31229 23489 31263
rect 23489 31229 23523 31263
rect 23523 31229 23532 31263
rect 23480 31220 23532 31229
rect 25504 31220 25556 31272
rect 19616 31084 19668 31136
rect 20720 31127 20772 31136
rect 20720 31093 20729 31127
rect 20729 31093 20763 31127
rect 20763 31093 20772 31127
rect 20720 31084 20772 31093
rect 22652 31084 22704 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 7656 30880 7708 30932
rect 8484 30880 8536 30932
rect 12164 30880 12216 30932
rect 14280 30880 14332 30932
rect 16672 30880 16724 30932
rect 17132 30923 17184 30932
rect 17132 30889 17141 30923
rect 17141 30889 17175 30923
rect 17175 30889 17184 30923
rect 17132 30880 17184 30889
rect 17868 30880 17920 30932
rect 6920 30744 6972 30796
rect 11152 30787 11204 30796
rect 11152 30753 11161 30787
rect 11161 30753 11195 30787
rect 11195 30753 11204 30787
rect 11152 30744 11204 30753
rect 11428 30787 11480 30796
rect 11428 30753 11437 30787
rect 11437 30753 11471 30787
rect 11471 30753 11480 30787
rect 11428 30744 11480 30753
rect 15844 30855 15896 30864
rect 15844 30821 15853 30855
rect 15853 30821 15887 30855
rect 15887 30821 15896 30855
rect 15844 30812 15896 30821
rect 17500 30812 17552 30864
rect 13912 30744 13964 30796
rect 14648 30787 14700 30796
rect 14648 30753 14657 30787
rect 14657 30753 14691 30787
rect 14691 30753 14700 30787
rect 14648 30744 14700 30753
rect 16028 30744 16080 30796
rect 16948 30744 17000 30796
rect 17868 30744 17920 30796
rect 7748 30676 7800 30728
rect 15200 30676 15252 30728
rect 10692 30608 10744 30660
rect 10876 30608 10928 30660
rect 18880 30719 18932 30728
rect 18880 30685 18889 30719
rect 18889 30685 18923 30719
rect 18923 30685 18932 30719
rect 18880 30676 18932 30685
rect 21180 30880 21232 30932
rect 22928 30812 22980 30864
rect 20076 30744 20128 30796
rect 23480 30744 23532 30796
rect 22836 30676 22888 30728
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 8392 30540 8444 30592
rect 11336 30540 11388 30592
rect 11888 30583 11940 30592
rect 11888 30549 11897 30583
rect 11897 30549 11931 30583
rect 11931 30549 11940 30583
rect 11888 30540 11940 30549
rect 12440 30540 12492 30592
rect 13728 30540 13780 30592
rect 15108 30540 15160 30592
rect 16304 30583 16356 30592
rect 16304 30549 16313 30583
rect 16313 30549 16347 30583
rect 16347 30549 16356 30583
rect 16304 30540 16356 30549
rect 17868 30608 17920 30660
rect 19708 30608 19760 30660
rect 19800 30651 19852 30660
rect 19800 30617 19809 30651
rect 19809 30617 19843 30651
rect 19843 30617 19852 30651
rect 19800 30608 19852 30617
rect 18328 30540 18380 30592
rect 19524 30540 19576 30592
rect 21088 30540 21140 30592
rect 21364 30540 21416 30592
rect 23296 30583 23348 30592
rect 23296 30549 23305 30583
rect 23305 30549 23339 30583
rect 23339 30549 23348 30583
rect 23296 30540 23348 30549
rect 23940 30540 23992 30592
rect 24860 30540 24912 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 9772 30336 9824 30388
rect 15476 30336 15528 30388
rect 16304 30336 16356 30388
rect 17408 30336 17460 30388
rect 17776 30336 17828 30388
rect 18328 30336 18380 30388
rect 25228 30336 25280 30388
rect 4344 30268 4396 30320
rect 8668 30268 8720 30320
rect 11888 30268 11940 30320
rect 12716 30268 12768 30320
rect 14740 30268 14792 30320
rect 8576 30200 8628 30252
rect 8852 30200 8904 30252
rect 11060 30200 11112 30252
rect 9588 30064 9640 30116
rect 9956 30107 10008 30116
rect 9956 30073 9965 30107
rect 9965 30073 9999 30107
rect 9999 30073 10008 30107
rect 9956 30064 10008 30073
rect 8668 30039 8720 30048
rect 8668 30005 8677 30039
rect 8677 30005 8711 30039
rect 8711 30005 8720 30039
rect 8668 29996 8720 30005
rect 8852 30039 8904 30048
rect 8852 30005 8861 30039
rect 8861 30005 8895 30039
rect 8895 30005 8904 30039
rect 8852 29996 8904 30005
rect 9864 29996 9916 30048
rect 11336 30132 11388 30184
rect 11888 30064 11940 30116
rect 17132 30268 17184 30320
rect 16948 30200 17000 30252
rect 19708 30268 19760 30320
rect 17500 30175 17552 30184
rect 17500 30141 17509 30175
rect 17509 30141 17543 30175
rect 17543 30141 17552 30175
rect 17500 30132 17552 30141
rect 19892 30200 19944 30252
rect 20444 30243 20496 30252
rect 20444 30209 20453 30243
rect 20453 30209 20487 30243
rect 20487 30209 20496 30243
rect 20444 30200 20496 30209
rect 24952 30268 25004 30320
rect 25412 30268 25464 30320
rect 23664 30243 23716 30252
rect 23664 30209 23673 30243
rect 23673 30209 23707 30243
rect 23707 30209 23716 30243
rect 23664 30200 23716 30209
rect 24492 30243 24544 30252
rect 24492 30209 24501 30243
rect 24501 30209 24535 30243
rect 24535 30209 24544 30243
rect 24492 30200 24544 30209
rect 17132 30064 17184 30116
rect 19248 30132 19300 30184
rect 19432 30132 19484 30184
rect 20904 30175 20956 30184
rect 20904 30141 20913 30175
rect 20913 30141 20947 30175
rect 20947 30141 20956 30175
rect 20904 30132 20956 30141
rect 19800 30064 19852 30116
rect 20260 30064 20312 30116
rect 20536 30064 20588 30116
rect 11796 30039 11848 30048
rect 11796 30005 11805 30039
rect 11805 30005 11839 30039
rect 11839 30005 11848 30039
rect 11796 29996 11848 30005
rect 12348 30039 12400 30048
rect 12348 30005 12357 30039
rect 12357 30005 12391 30039
rect 12391 30005 12400 30039
rect 12348 29996 12400 30005
rect 14372 29996 14424 30048
rect 18420 29996 18472 30048
rect 19984 29996 20036 30048
rect 20444 29996 20496 30048
rect 21916 29996 21968 30048
rect 24032 29996 24084 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 5080 29792 5132 29844
rect 8576 29792 8628 29844
rect 11888 29835 11940 29844
rect 11888 29801 11897 29835
rect 11897 29801 11931 29835
rect 11931 29801 11940 29835
rect 11888 29792 11940 29801
rect 13912 29792 13964 29844
rect 15292 29792 15344 29844
rect 16580 29792 16632 29844
rect 17684 29792 17736 29844
rect 18052 29792 18104 29844
rect 21824 29792 21876 29844
rect 23296 29792 23348 29844
rect 25412 29835 25464 29844
rect 25412 29801 25421 29835
rect 25421 29801 25455 29835
rect 25455 29801 25464 29835
rect 25412 29792 25464 29801
rect 4068 29699 4120 29708
rect 4068 29665 4077 29699
rect 4077 29665 4111 29699
rect 4111 29665 4120 29699
rect 4068 29656 4120 29665
rect 11244 29699 11296 29708
rect 11244 29665 11253 29699
rect 11253 29665 11287 29699
rect 11287 29665 11296 29699
rect 11244 29656 11296 29665
rect 11520 29699 11572 29708
rect 11520 29665 11529 29699
rect 11529 29665 11563 29699
rect 11563 29665 11572 29699
rect 11520 29656 11572 29665
rect 3516 29520 3568 29572
rect 6184 29520 6236 29572
rect 17224 29656 17276 29708
rect 18052 29656 18104 29708
rect 18420 29699 18472 29708
rect 18420 29665 18429 29699
rect 18429 29665 18463 29699
rect 18463 29665 18472 29699
rect 18420 29656 18472 29665
rect 18880 29656 18932 29708
rect 19432 29656 19484 29708
rect 19800 29699 19852 29708
rect 19800 29665 19809 29699
rect 19809 29665 19843 29699
rect 19843 29665 19852 29699
rect 19800 29656 19852 29665
rect 16764 29520 16816 29572
rect 17868 29520 17920 29572
rect 18420 29520 18472 29572
rect 20812 29588 20864 29640
rect 20996 29724 21048 29776
rect 22192 29656 22244 29708
rect 19800 29520 19852 29572
rect 10324 29452 10376 29504
rect 10876 29452 10928 29504
rect 16948 29452 17000 29504
rect 19064 29452 19116 29504
rect 19984 29452 20036 29504
rect 21824 29520 21876 29572
rect 22928 29699 22980 29708
rect 22928 29665 22937 29699
rect 22937 29665 22971 29699
rect 22971 29665 22980 29699
rect 22928 29656 22980 29665
rect 23480 29656 23532 29708
rect 22744 29588 22796 29640
rect 24676 29588 24728 29640
rect 21456 29452 21508 29504
rect 21640 29495 21692 29504
rect 21640 29461 21649 29495
rect 21649 29461 21683 29495
rect 21683 29461 21692 29495
rect 21640 29452 21692 29461
rect 21916 29452 21968 29504
rect 24952 29520 25004 29572
rect 24676 29452 24728 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 3976 29248 4028 29300
rect 8392 29291 8444 29300
rect 8392 29257 8401 29291
rect 8401 29257 8435 29291
rect 8435 29257 8444 29291
rect 8392 29248 8444 29257
rect 8576 29248 8628 29300
rect 9128 29248 9180 29300
rect 15568 29248 15620 29300
rect 15844 29291 15896 29300
rect 15844 29257 15853 29291
rect 15853 29257 15887 29291
rect 15887 29257 15896 29291
rect 15844 29248 15896 29257
rect 20536 29248 20588 29300
rect 21640 29248 21692 29300
rect 3608 29112 3660 29164
rect 7656 29155 7708 29164
rect 7656 29121 7665 29155
rect 7665 29121 7699 29155
rect 7699 29121 7708 29155
rect 7656 29112 7708 29121
rect 10324 29155 10376 29164
rect 10324 29121 10333 29155
rect 10333 29121 10367 29155
rect 10367 29121 10376 29155
rect 10324 29112 10376 29121
rect 11060 29112 11112 29164
rect 7380 28976 7432 29028
rect 8944 29087 8996 29096
rect 8944 29053 8953 29087
rect 8953 29053 8987 29087
rect 8987 29053 8996 29087
rect 8944 29044 8996 29053
rect 14188 29180 14240 29232
rect 15384 29180 15436 29232
rect 15660 29180 15712 29232
rect 17040 29180 17092 29232
rect 20904 29180 20956 29232
rect 23756 29180 23808 29232
rect 24768 29223 24820 29232
rect 24768 29189 24777 29223
rect 24777 29189 24811 29223
rect 24811 29189 24820 29223
rect 24768 29180 24820 29189
rect 12348 29155 12400 29164
rect 12348 29121 12357 29155
rect 12357 29121 12391 29155
rect 12391 29121 12400 29155
rect 12348 29112 12400 29121
rect 15568 29112 15620 29164
rect 16856 29112 16908 29164
rect 17500 29112 17552 29164
rect 9404 28976 9456 29028
rect 11428 28976 11480 29028
rect 14096 29087 14148 29096
rect 14096 29053 14105 29087
rect 14105 29053 14139 29087
rect 14139 29053 14148 29087
rect 14096 29044 14148 29053
rect 15936 29087 15988 29096
rect 15936 29053 15945 29087
rect 15945 29053 15979 29087
rect 15979 29053 15988 29087
rect 15936 29044 15988 29053
rect 12624 28976 12676 29028
rect 15384 29019 15436 29028
rect 15384 28985 15393 29019
rect 15393 28985 15427 29019
rect 15427 28985 15436 29019
rect 15384 28976 15436 28985
rect 15660 28976 15712 29028
rect 16764 29019 16816 29028
rect 16764 28985 16773 29019
rect 16773 28985 16807 29019
rect 16807 28985 16816 29019
rect 16764 28976 16816 28985
rect 17776 29044 17828 29096
rect 19064 29155 19116 29164
rect 19064 29121 19073 29155
rect 19073 29121 19107 29155
rect 19107 29121 19116 29155
rect 19064 29112 19116 29121
rect 19800 29112 19852 29164
rect 7012 28951 7064 28960
rect 7012 28917 7021 28951
rect 7021 28917 7055 28951
rect 7055 28917 7064 28951
rect 7012 28908 7064 28917
rect 9680 28951 9732 28960
rect 9680 28917 9689 28951
rect 9689 28917 9723 28951
rect 9723 28917 9732 28951
rect 9680 28908 9732 28917
rect 17500 28951 17552 28960
rect 17500 28917 17509 28951
rect 17509 28917 17543 28951
rect 17543 28917 17552 28951
rect 17500 28908 17552 28917
rect 18328 28976 18380 29028
rect 19432 29044 19484 29096
rect 18420 28908 18472 28960
rect 19892 28976 19944 29028
rect 22376 29044 22428 29096
rect 23940 29155 23992 29164
rect 23940 29121 23949 29155
rect 23949 29121 23983 29155
rect 23983 29121 23992 29155
rect 23940 29112 23992 29121
rect 23296 28976 23348 29028
rect 24308 29019 24360 29028
rect 24308 28985 24317 29019
rect 24317 28985 24351 29019
rect 24351 28985 24360 29019
rect 24308 28976 24360 28985
rect 20536 28951 20588 28960
rect 20536 28917 20545 28951
rect 20545 28917 20579 28951
rect 20579 28917 20588 28951
rect 20536 28908 20588 28917
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 18420 28704 18472 28756
rect 11060 28636 11112 28688
rect 4160 28568 4212 28620
rect 5724 28611 5776 28620
rect 5724 28577 5733 28611
rect 5733 28577 5767 28611
rect 5767 28577 5776 28611
rect 5724 28568 5776 28577
rect 12348 28568 12400 28620
rect 12808 28611 12860 28620
rect 12808 28577 12817 28611
rect 12817 28577 12851 28611
rect 12851 28577 12860 28611
rect 12808 28568 12860 28577
rect 14096 28568 14148 28620
rect 14740 28611 14792 28620
rect 14740 28577 14749 28611
rect 14749 28577 14783 28611
rect 14783 28577 14792 28611
rect 14740 28568 14792 28577
rect 16580 28611 16632 28620
rect 16580 28577 16589 28611
rect 16589 28577 16623 28611
rect 16623 28577 16632 28611
rect 16580 28568 16632 28577
rect 17592 28568 17644 28620
rect 18788 28636 18840 28688
rect 18972 28704 19024 28756
rect 22560 28704 22612 28756
rect 22744 28704 22796 28756
rect 18236 28611 18288 28620
rect 18236 28577 18245 28611
rect 18245 28577 18279 28611
rect 18279 28577 18288 28611
rect 18236 28568 18288 28577
rect 18420 28568 18472 28620
rect 19064 28568 19116 28620
rect 20536 28568 20588 28620
rect 8576 28543 8628 28552
rect 8576 28509 8585 28543
rect 8585 28509 8619 28543
rect 8619 28509 8628 28543
rect 8576 28500 8628 28509
rect 9772 28543 9824 28552
rect 9772 28509 9781 28543
rect 9781 28509 9815 28543
rect 9815 28509 9824 28543
rect 9772 28500 9824 28509
rect 11520 28500 11572 28552
rect 3424 28432 3476 28484
rect 7748 28432 7800 28484
rect 17500 28500 17552 28552
rect 15752 28432 15804 28484
rect 22192 28500 22244 28552
rect 24400 28500 24452 28552
rect 7656 28364 7708 28416
rect 10876 28364 10928 28416
rect 13452 28364 13504 28416
rect 13544 28364 13596 28416
rect 14740 28364 14792 28416
rect 15568 28407 15620 28416
rect 15568 28373 15577 28407
rect 15577 28373 15611 28407
rect 15611 28373 15620 28407
rect 15568 28364 15620 28373
rect 17040 28364 17092 28416
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 17592 28364 17644 28373
rect 17684 28364 17736 28416
rect 18236 28364 18288 28416
rect 18420 28364 18472 28416
rect 19248 28364 19300 28416
rect 19432 28407 19484 28416
rect 19432 28373 19441 28407
rect 19441 28373 19475 28407
rect 19475 28373 19484 28407
rect 19432 28364 19484 28373
rect 21548 28432 21600 28484
rect 22468 28432 22520 28484
rect 23020 28432 23072 28484
rect 25136 28432 25188 28484
rect 23480 28364 23532 28416
rect 24308 28364 24360 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 7840 28160 7892 28212
rect 12808 28160 12860 28212
rect 13452 28160 13504 28212
rect 15660 28160 15712 28212
rect 16580 28160 16632 28212
rect 17684 28160 17736 28212
rect 18236 28160 18288 28212
rect 18420 28160 18472 28212
rect 18972 28203 19024 28212
rect 18972 28169 18981 28203
rect 18981 28169 19015 28203
rect 19015 28169 19024 28203
rect 19708 28203 19760 28212
rect 18972 28160 19024 28169
rect 19708 28169 19717 28203
rect 19717 28169 19751 28203
rect 19751 28169 19760 28203
rect 19708 28160 19760 28169
rect 19892 28160 19944 28212
rect 7012 28092 7064 28144
rect 7748 28092 7800 28144
rect 13360 28092 13412 28144
rect 14464 28092 14516 28144
rect 17500 28092 17552 28144
rect 21180 28092 21232 28144
rect 6828 27999 6880 28008
rect 6828 27965 6837 27999
rect 6837 27965 6871 27999
rect 6871 27965 6880 27999
rect 6828 27956 6880 27965
rect 7748 27956 7800 28008
rect 12348 28067 12400 28076
rect 12348 28033 12357 28067
rect 12357 28033 12391 28067
rect 12391 28033 12400 28067
rect 12348 28024 12400 28033
rect 9772 27956 9824 28008
rect 12440 27956 12492 28008
rect 14280 27820 14332 27872
rect 15936 28024 15988 28076
rect 17868 28067 17920 28076
rect 16304 27888 16356 27940
rect 17868 28033 17877 28067
rect 17877 28033 17911 28067
rect 17911 28033 17920 28067
rect 17868 28024 17920 28033
rect 19248 28024 19300 28076
rect 18604 27956 18656 28008
rect 18880 27956 18932 28008
rect 19708 27956 19760 28008
rect 21364 28024 21416 28076
rect 23296 28160 23348 28212
rect 24124 28092 24176 28144
rect 22468 28024 22520 28076
rect 21180 27999 21232 28008
rect 21180 27965 21189 27999
rect 21189 27965 21223 27999
rect 21223 27965 21232 27999
rect 21180 27956 21232 27965
rect 23020 27956 23072 28008
rect 23572 27999 23624 28008
rect 23572 27965 23581 27999
rect 23581 27965 23615 27999
rect 23615 27965 23624 27999
rect 23572 27956 23624 27965
rect 15016 27863 15068 27872
rect 15016 27829 15025 27863
rect 15025 27829 15059 27863
rect 15059 27829 15068 27863
rect 15016 27820 15068 27829
rect 16396 27820 16448 27872
rect 18328 27820 18380 27872
rect 18880 27820 18932 27872
rect 19248 27820 19300 27872
rect 19708 27820 19760 27872
rect 22008 27888 22060 27940
rect 20628 27820 20680 27872
rect 23388 27820 23440 27872
rect 24584 27931 24636 27940
rect 24584 27897 24593 27931
rect 24593 27897 24627 27931
rect 24627 27897 24636 27931
rect 24584 27888 24636 27897
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 9680 27616 9732 27668
rect 12348 27616 12400 27668
rect 14096 27616 14148 27668
rect 16856 27616 16908 27668
rect 19800 27616 19852 27668
rect 12256 27548 12308 27600
rect 17408 27548 17460 27600
rect 17684 27548 17736 27600
rect 20260 27548 20312 27600
rect 2780 27523 2832 27532
rect 2780 27489 2789 27523
rect 2789 27489 2823 27523
rect 2823 27489 2832 27523
rect 2780 27480 2832 27489
rect 3608 27480 3660 27532
rect 3884 27480 3936 27532
rect 7656 27480 7708 27532
rect 12072 27480 12124 27532
rect 4252 27344 4304 27396
rect 5908 27344 5960 27396
rect 6552 27344 6604 27396
rect 9312 27455 9364 27464
rect 9312 27421 9321 27455
rect 9321 27421 9355 27455
rect 9355 27421 9364 27455
rect 9312 27412 9364 27421
rect 9496 27344 9548 27396
rect 11152 27344 11204 27396
rect 13636 27480 13688 27532
rect 14924 27480 14976 27532
rect 16120 27480 16172 27532
rect 17592 27480 17644 27532
rect 14188 27412 14240 27464
rect 16580 27412 16632 27464
rect 17868 27412 17920 27464
rect 18236 27480 18288 27532
rect 4528 27276 4580 27328
rect 7104 27276 7156 27328
rect 8852 27276 8904 27328
rect 15108 27344 15160 27396
rect 15476 27387 15528 27396
rect 15476 27353 15485 27387
rect 15485 27353 15519 27387
rect 15519 27353 15528 27387
rect 15476 27344 15528 27353
rect 18880 27412 18932 27464
rect 19800 27455 19852 27464
rect 19800 27421 19809 27455
rect 19809 27421 19843 27455
rect 19843 27421 19852 27455
rect 19800 27412 19852 27421
rect 20076 27480 20128 27532
rect 22560 27480 22612 27532
rect 23848 27480 23900 27532
rect 21364 27412 21416 27464
rect 23388 27455 23440 27464
rect 23388 27421 23397 27455
rect 23397 27421 23431 27455
rect 23431 27421 23440 27455
rect 23388 27412 23440 27421
rect 24308 27412 24360 27464
rect 11980 27319 12032 27328
rect 11980 27285 11989 27319
rect 11989 27285 12023 27319
rect 12023 27285 12032 27319
rect 11980 27276 12032 27285
rect 12716 27276 12768 27328
rect 13452 27319 13504 27328
rect 13452 27285 13461 27319
rect 13461 27285 13495 27319
rect 13495 27285 13504 27319
rect 13452 27276 13504 27285
rect 14188 27319 14240 27328
rect 14188 27285 14197 27319
rect 14197 27285 14231 27319
rect 14231 27285 14240 27319
rect 14188 27276 14240 27285
rect 14464 27276 14516 27328
rect 14832 27276 14884 27328
rect 20536 27344 20588 27396
rect 21272 27344 21324 27396
rect 22560 27344 22612 27396
rect 17500 27319 17552 27328
rect 17500 27285 17509 27319
rect 17509 27285 17543 27319
rect 17543 27285 17552 27319
rect 17500 27276 17552 27285
rect 19340 27276 19392 27328
rect 19708 27319 19760 27328
rect 19708 27285 19717 27319
rect 19717 27285 19751 27319
rect 19751 27285 19760 27319
rect 19708 27276 19760 27285
rect 20168 27319 20220 27328
rect 20168 27285 20177 27319
rect 20177 27285 20211 27319
rect 20211 27285 20220 27319
rect 20168 27276 20220 27285
rect 20904 27319 20956 27328
rect 20904 27285 20913 27319
rect 20913 27285 20947 27319
rect 20947 27285 20956 27319
rect 20904 27276 20956 27285
rect 22192 27276 22244 27328
rect 23480 27276 23532 27328
rect 24492 27276 24544 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 3516 27072 3568 27124
rect 6552 27115 6604 27124
rect 6552 27081 6561 27115
rect 6561 27081 6595 27115
rect 6595 27081 6604 27115
rect 6552 27072 6604 27081
rect 7840 27072 7892 27124
rect 7748 27004 7800 27056
rect 11980 27072 12032 27124
rect 13728 27072 13780 27124
rect 11704 27004 11756 27056
rect 3332 26979 3384 26988
rect 3332 26945 3376 26979
rect 3376 26945 3384 26979
rect 3332 26936 3384 26945
rect 3792 26936 3844 26988
rect 8576 26936 8628 26988
rect 9036 26936 9088 26988
rect 3608 26868 3660 26920
rect 6184 26868 6236 26920
rect 4436 26775 4488 26784
rect 4436 26741 4445 26775
rect 4445 26741 4479 26775
rect 4479 26741 4488 26775
rect 4436 26732 4488 26741
rect 9036 26775 9088 26784
rect 9036 26741 9045 26775
rect 9045 26741 9079 26775
rect 9079 26741 9088 26775
rect 9036 26732 9088 26741
rect 11888 26936 11940 26988
rect 11152 26911 11204 26920
rect 11152 26877 11161 26911
rect 11161 26877 11195 26911
rect 11195 26877 11204 26911
rect 11152 26868 11204 26877
rect 11244 26868 11296 26920
rect 9772 26800 9824 26852
rect 13636 27004 13688 27056
rect 14924 27004 14976 27056
rect 15660 27047 15712 27056
rect 15660 27013 15669 27047
rect 15669 27013 15703 27047
rect 15703 27013 15712 27047
rect 15660 27004 15712 27013
rect 18420 27072 18472 27124
rect 20904 27072 20956 27124
rect 21364 27115 21416 27124
rect 21364 27081 21373 27115
rect 21373 27081 21407 27115
rect 21407 27081 21416 27115
rect 21364 27072 21416 27081
rect 23296 27072 23348 27124
rect 23848 27115 23900 27124
rect 23848 27081 23857 27115
rect 23857 27081 23891 27115
rect 23891 27081 23900 27115
rect 23848 27072 23900 27081
rect 20352 27004 20404 27056
rect 14464 26936 14516 26988
rect 12440 26868 12492 26920
rect 15016 26868 15068 26920
rect 17592 26936 17644 26988
rect 17776 26936 17828 26988
rect 20444 26979 20496 26988
rect 20444 26945 20453 26979
rect 20453 26945 20487 26979
rect 20487 26945 20496 26979
rect 20444 26936 20496 26945
rect 16028 26868 16080 26920
rect 16764 26868 16816 26920
rect 17316 26911 17368 26920
rect 17316 26877 17325 26911
rect 17325 26877 17359 26911
rect 17359 26877 17368 26911
rect 17316 26868 17368 26877
rect 15108 26800 15160 26852
rect 17684 26868 17736 26920
rect 11152 26732 11204 26784
rect 14464 26732 14516 26784
rect 14740 26732 14792 26784
rect 15016 26732 15068 26784
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 17316 26732 17368 26784
rect 19432 26868 19484 26920
rect 19524 26911 19576 26920
rect 19524 26877 19533 26911
rect 19533 26877 19567 26911
rect 19567 26877 19576 26911
rect 19524 26868 19576 26877
rect 20076 26868 20128 26920
rect 19248 26800 19300 26852
rect 21732 26936 21784 26988
rect 22744 26936 22796 26988
rect 23572 27004 23624 27056
rect 23296 26936 23348 26988
rect 20812 26868 20864 26920
rect 21456 26868 21508 26920
rect 22100 26911 22152 26920
rect 22100 26877 22109 26911
rect 22109 26877 22143 26911
rect 22143 26877 22152 26911
rect 22100 26868 22152 26877
rect 22468 26800 22520 26852
rect 19432 26732 19484 26784
rect 19708 26732 19760 26784
rect 23388 26800 23440 26852
rect 22652 26732 22704 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 3792 26571 3844 26580
rect 3792 26537 3801 26571
rect 3801 26537 3835 26571
rect 3835 26537 3844 26571
rect 3792 26528 3844 26537
rect 5908 26528 5960 26580
rect 8852 26528 8904 26580
rect 14188 26528 14240 26580
rect 11428 26460 11480 26512
rect 12992 26460 13044 26512
rect 7104 26435 7156 26444
rect 7104 26401 7113 26435
rect 7113 26401 7147 26435
rect 7147 26401 7156 26435
rect 7104 26392 7156 26401
rect 7748 26392 7800 26444
rect 4436 26324 4488 26376
rect 6828 26367 6880 26376
rect 6828 26333 6837 26367
rect 6837 26333 6871 26367
rect 6871 26333 6880 26367
rect 6828 26324 6880 26333
rect 11060 26435 11112 26444
rect 11060 26401 11069 26435
rect 11069 26401 11103 26435
rect 11103 26401 11112 26435
rect 11060 26392 11112 26401
rect 11152 26435 11204 26444
rect 11152 26401 11161 26435
rect 11161 26401 11195 26435
rect 11195 26401 11204 26435
rect 11152 26392 11204 26401
rect 11704 26392 11756 26444
rect 14280 26460 14332 26512
rect 14556 26460 14608 26512
rect 15016 26460 15068 26512
rect 15476 26528 15528 26580
rect 16396 26528 16448 26580
rect 16672 26460 16724 26512
rect 17316 26460 17368 26512
rect 20352 26571 20404 26580
rect 20352 26537 20361 26571
rect 20361 26537 20395 26571
rect 20395 26537 20404 26571
rect 20352 26528 20404 26537
rect 20628 26528 20680 26580
rect 19708 26460 19760 26512
rect 20812 26460 20864 26512
rect 14832 26392 14884 26444
rect 15660 26392 15712 26444
rect 11244 26367 11296 26376
rect 11244 26333 11253 26367
rect 11253 26333 11287 26367
rect 11287 26333 11296 26367
rect 11244 26324 11296 26333
rect 14740 26324 14792 26376
rect 17592 26392 17644 26444
rect 21732 26392 21784 26444
rect 23112 26435 23164 26444
rect 23112 26401 23121 26435
rect 23121 26401 23155 26435
rect 23155 26401 23164 26435
rect 23112 26392 23164 26401
rect 19248 26324 19300 26376
rect 22192 26324 22244 26376
rect 22560 26324 22612 26376
rect 22744 26324 22796 26376
rect 23664 26324 23716 26376
rect 24032 26324 24084 26376
rect 9220 26256 9272 26308
rect 10048 26256 10100 26308
rect 11612 26256 11664 26308
rect 14924 26256 14976 26308
rect 16764 26256 16816 26308
rect 5540 26231 5592 26240
rect 5540 26197 5549 26231
rect 5549 26197 5583 26231
rect 5583 26197 5592 26231
rect 5540 26188 5592 26197
rect 13360 26231 13412 26240
rect 13360 26197 13369 26231
rect 13369 26197 13403 26231
rect 13403 26197 13412 26231
rect 13360 26188 13412 26197
rect 14648 26188 14700 26240
rect 15200 26188 15252 26240
rect 17132 26188 17184 26240
rect 17776 26188 17828 26240
rect 22376 26256 22428 26308
rect 23388 26256 23440 26308
rect 23756 26299 23808 26308
rect 23756 26265 23765 26299
rect 23765 26265 23799 26299
rect 23799 26265 23808 26299
rect 23756 26256 23808 26265
rect 24124 26256 24176 26308
rect 22560 26231 22612 26240
rect 22560 26197 22569 26231
rect 22569 26197 22603 26231
rect 22603 26197 22612 26231
rect 22560 26188 22612 26197
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 3424 25984 3476 26036
rect 5540 25984 5592 26036
rect 12992 26027 13044 26036
rect 12992 25993 13001 26027
rect 13001 25993 13035 26027
rect 13035 25993 13044 26027
rect 12992 25984 13044 25993
rect 13268 25984 13320 26036
rect 15936 25984 15988 26036
rect 3424 25848 3476 25900
rect 6828 25916 6880 25968
rect 8576 25916 8628 25968
rect 9220 25916 9272 25968
rect 13544 25916 13596 25968
rect 16580 25984 16632 26036
rect 18328 26027 18380 26036
rect 18328 25993 18337 26027
rect 18337 25993 18371 26027
rect 18371 25993 18380 26027
rect 18328 25984 18380 25993
rect 19064 25984 19116 26036
rect 16120 25916 16172 25968
rect 7748 25823 7800 25832
rect 7748 25789 7757 25823
rect 7757 25789 7791 25823
rect 7791 25789 7800 25823
rect 7748 25780 7800 25789
rect 8852 25780 8904 25832
rect 11888 25848 11940 25900
rect 12348 25848 12400 25900
rect 19156 25916 19208 25968
rect 19524 25984 19576 26036
rect 20444 25959 20496 25968
rect 20444 25925 20453 25959
rect 20453 25925 20487 25959
rect 20487 25925 20496 25959
rect 20444 25916 20496 25925
rect 12532 25780 12584 25832
rect 17132 25848 17184 25900
rect 19432 25848 19484 25900
rect 23204 25984 23256 26036
rect 22284 25916 22336 25968
rect 24492 25959 24544 25968
rect 24492 25925 24501 25959
rect 24501 25925 24535 25959
rect 24535 25925 24544 25959
rect 24492 25916 24544 25925
rect 16028 25823 16080 25832
rect 16028 25789 16037 25823
rect 16037 25789 16071 25823
rect 16071 25789 16080 25823
rect 16028 25780 16080 25789
rect 9680 25712 9732 25764
rect 4160 25644 4212 25696
rect 5816 25687 5868 25696
rect 5816 25653 5825 25687
rect 5825 25653 5859 25687
rect 5859 25653 5868 25687
rect 5816 25644 5868 25653
rect 12808 25644 12860 25696
rect 13268 25644 13320 25696
rect 13636 25644 13688 25696
rect 18328 25644 18380 25696
rect 19340 25823 19392 25832
rect 19340 25789 19349 25823
rect 19349 25789 19383 25823
rect 19383 25789 19392 25823
rect 19340 25780 19392 25789
rect 22836 25780 22888 25832
rect 23204 25848 23256 25900
rect 23388 25848 23440 25900
rect 24768 25823 24820 25832
rect 24768 25789 24777 25823
rect 24777 25789 24811 25823
rect 24811 25789 24820 25823
rect 24768 25780 24820 25789
rect 18696 25712 18748 25764
rect 20904 25712 20956 25764
rect 19432 25644 19484 25696
rect 19524 25644 19576 25696
rect 19708 25644 19760 25696
rect 19892 25644 19944 25696
rect 22376 25687 22428 25696
rect 22376 25653 22385 25687
rect 22385 25653 22419 25687
rect 22419 25653 22428 25687
rect 22376 25644 22428 25653
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 4160 25440 4212 25492
rect 4436 25483 4488 25492
rect 4436 25449 4445 25483
rect 4445 25449 4479 25483
rect 4479 25449 4488 25483
rect 4436 25440 4488 25449
rect 11428 25440 11480 25492
rect 13360 25440 13412 25492
rect 16028 25440 16080 25492
rect 12072 25372 12124 25424
rect 14372 25372 14424 25424
rect 6828 25304 6880 25356
rect 7104 25304 7156 25356
rect 7840 25304 7892 25356
rect 8852 25304 8904 25356
rect 9496 25304 9548 25356
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 12808 25304 12860 25356
rect 14740 25304 14792 25356
rect 3792 25236 3844 25288
rect 4436 25236 4488 25288
rect 6276 25236 6328 25288
rect 7748 25236 7800 25288
rect 8300 25236 8352 25288
rect 10232 25236 10284 25288
rect 12532 25279 12584 25288
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 14648 25236 14700 25288
rect 16028 25236 16080 25288
rect 21916 25372 21968 25424
rect 17224 25304 17276 25356
rect 18696 25304 18748 25356
rect 18880 25304 18932 25356
rect 20168 25236 20220 25288
rect 21272 25304 21324 25356
rect 22008 25304 22060 25356
rect 22468 25304 22520 25356
rect 24308 25304 24360 25356
rect 21640 25236 21692 25288
rect 23480 25236 23532 25288
rect 23940 25236 23992 25288
rect 24860 25279 24912 25288
rect 24860 25245 24869 25279
rect 24869 25245 24903 25279
rect 24903 25245 24912 25279
rect 24860 25236 24912 25245
rect 5816 25168 5868 25220
rect 7656 25168 7708 25220
rect 3332 25100 3384 25152
rect 6368 25100 6420 25152
rect 9496 25143 9548 25152
rect 9496 25109 9505 25143
rect 9505 25109 9539 25143
rect 9539 25109 9548 25143
rect 9496 25100 9548 25109
rect 10232 25143 10284 25152
rect 10232 25109 10241 25143
rect 10241 25109 10275 25143
rect 10275 25109 10284 25143
rect 10232 25100 10284 25109
rect 14096 25168 14148 25220
rect 15384 25168 15436 25220
rect 16764 25168 16816 25220
rect 17776 25168 17828 25220
rect 20720 25168 20772 25220
rect 20904 25211 20956 25220
rect 20904 25177 20913 25211
rect 20913 25177 20947 25211
rect 20947 25177 20956 25211
rect 20904 25168 20956 25177
rect 22100 25168 22152 25220
rect 22468 25168 22520 25220
rect 11428 25100 11480 25152
rect 13728 25100 13780 25152
rect 15476 25100 15528 25152
rect 15844 25100 15896 25152
rect 19708 25100 19760 25152
rect 20444 25100 20496 25152
rect 21732 25100 21784 25152
rect 22284 25100 22336 25152
rect 23940 25143 23992 25152
rect 23940 25109 23949 25143
rect 23949 25109 23983 25143
rect 23983 25109 23992 25143
rect 23940 25100 23992 25109
rect 24032 25100 24084 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 7196 24896 7248 24948
rect 7656 24939 7708 24948
rect 7656 24905 7665 24939
rect 7665 24905 7699 24939
rect 7699 24905 7708 24939
rect 7656 24896 7708 24905
rect 9496 24896 9548 24948
rect 16764 24939 16816 24948
rect 16764 24905 16773 24939
rect 16773 24905 16807 24939
rect 16807 24905 16816 24939
rect 16764 24896 16816 24905
rect 19892 24939 19944 24948
rect 19892 24905 19901 24939
rect 19901 24905 19935 24939
rect 19935 24905 19944 24939
rect 19892 24896 19944 24905
rect 22284 24896 22336 24948
rect 9680 24871 9732 24880
rect 9680 24837 9689 24871
rect 9689 24837 9723 24871
rect 9723 24837 9732 24871
rect 9680 24828 9732 24837
rect 6552 24760 6604 24812
rect 9312 24760 9364 24812
rect 2872 24735 2924 24744
rect 2872 24701 2881 24735
rect 2881 24701 2915 24735
rect 2915 24701 2924 24735
rect 2872 24692 2924 24701
rect 3332 24692 3384 24744
rect 9220 24692 9272 24744
rect 11980 24760 12032 24812
rect 4344 24624 4396 24676
rect 4528 24556 4580 24608
rect 6368 24599 6420 24608
rect 6368 24565 6377 24599
rect 6377 24565 6411 24599
rect 6411 24565 6420 24599
rect 6368 24556 6420 24565
rect 11152 24599 11204 24608
rect 11152 24565 11161 24599
rect 11161 24565 11195 24599
rect 11195 24565 11204 24599
rect 11152 24556 11204 24565
rect 11704 24599 11756 24608
rect 11704 24565 11713 24599
rect 11713 24565 11747 24599
rect 11747 24565 11756 24599
rect 11704 24556 11756 24565
rect 11980 24556 12032 24608
rect 12348 24556 12400 24608
rect 14832 24760 14884 24812
rect 15844 24803 15896 24812
rect 15844 24769 15853 24803
rect 15853 24769 15887 24803
rect 15887 24769 15896 24803
rect 15844 24760 15896 24769
rect 16120 24760 16172 24812
rect 16396 24760 16448 24812
rect 19984 24803 20036 24812
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 20996 24803 21048 24812
rect 20996 24769 21005 24803
rect 21005 24769 21039 24803
rect 21039 24769 21048 24803
rect 20996 24760 21048 24769
rect 21180 24760 21232 24812
rect 17684 24692 17736 24744
rect 18696 24735 18748 24744
rect 18696 24701 18705 24735
rect 18705 24701 18739 24735
rect 18739 24701 18748 24735
rect 18696 24692 18748 24701
rect 17132 24624 17184 24676
rect 14832 24556 14884 24608
rect 16580 24556 16632 24608
rect 20352 24692 20404 24744
rect 23848 24760 23900 24812
rect 19156 24624 19208 24676
rect 22836 24624 22888 24676
rect 24676 24735 24728 24744
rect 24676 24701 24685 24735
rect 24685 24701 24719 24735
rect 24719 24701 24728 24735
rect 24676 24692 24728 24701
rect 24860 24624 24912 24676
rect 19340 24556 19392 24608
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 6092 24352 6144 24404
rect 6276 24352 6328 24404
rect 7104 24259 7156 24268
rect 7104 24225 7113 24259
rect 7113 24225 7147 24259
rect 7147 24225 7156 24259
rect 7104 24216 7156 24225
rect 8392 24216 8444 24268
rect 14924 24352 14976 24404
rect 15752 24352 15804 24404
rect 18696 24352 18748 24404
rect 10324 24259 10376 24268
rect 10324 24225 10333 24259
rect 10333 24225 10367 24259
rect 10367 24225 10376 24259
rect 10324 24216 10376 24225
rect 12440 24216 12492 24268
rect 17132 24259 17184 24268
rect 17132 24225 17141 24259
rect 17141 24225 17175 24259
rect 17175 24225 17184 24259
rect 17132 24216 17184 24225
rect 20536 24216 20588 24268
rect 3608 24148 3660 24200
rect 4160 24148 4212 24200
rect 7656 24148 7708 24200
rect 9312 24148 9364 24200
rect 11428 24191 11480 24200
rect 11428 24157 11437 24191
rect 11437 24157 11471 24191
rect 11471 24157 11480 24191
rect 11428 24148 11480 24157
rect 17868 24148 17920 24200
rect 19340 24148 19392 24200
rect 6368 24080 6420 24132
rect 1768 24012 1820 24064
rect 4620 24012 4672 24064
rect 11704 24123 11756 24132
rect 11704 24089 11713 24123
rect 11713 24089 11747 24123
rect 11747 24089 11756 24123
rect 11704 24080 11756 24089
rect 12348 24080 12400 24132
rect 16396 24080 16448 24132
rect 7472 24012 7524 24064
rect 8852 24012 8904 24064
rect 9956 24012 10008 24064
rect 13820 24012 13872 24064
rect 16028 24012 16080 24064
rect 23388 24352 23440 24404
rect 21640 24327 21692 24336
rect 21640 24293 21649 24327
rect 21649 24293 21683 24327
rect 21683 24293 21692 24327
rect 21640 24284 21692 24293
rect 24032 24191 24084 24200
rect 24032 24157 24041 24191
rect 24041 24157 24075 24191
rect 24075 24157 24084 24191
rect 24032 24148 24084 24157
rect 22836 24123 22888 24132
rect 22836 24089 22845 24123
rect 22845 24089 22879 24123
rect 22879 24089 22888 24123
rect 22836 24080 22888 24089
rect 24400 24080 24452 24132
rect 22744 24012 22796 24064
rect 23296 24012 23348 24064
rect 23388 24012 23440 24064
rect 24676 24055 24728 24064
rect 24676 24021 24685 24055
rect 24685 24021 24719 24055
rect 24719 24021 24728 24055
rect 24676 24012 24728 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 4252 23808 4304 23860
rect 9128 23808 9180 23860
rect 9956 23851 10008 23860
rect 9956 23817 9965 23851
rect 9965 23817 9999 23851
rect 9999 23817 10008 23851
rect 9956 23808 10008 23817
rect 10692 23851 10744 23860
rect 10692 23817 10701 23851
rect 10701 23817 10735 23851
rect 10735 23817 10744 23851
rect 10692 23808 10744 23817
rect 12072 23808 12124 23860
rect 16120 23808 16172 23860
rect 16580 23808 16632 23860
rect 17500 23808 17552 23860
rect 20996 23808 21048 23860
rect 21548 23808 21600 23860
rect 23572 23808 23624 23860
rect 4068 23715 4120 23724
rect 4068 23681 4112 23715
rect 4112 23681 4120 23715
rect 4068 23672 4120 23681
rect 11152 23740 11204 23792
rect 20904 23740 20956 23792
rect 21088 23740 21140 23792
rect 24676 23740 24728 23792
rect 11336 23672 11388 23724
rect 12256 23672 12308 23724
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 11888 23647 11940 23656
rect 11888 23613 11897 23647
rect 11897 23613 11931 23647
rect 11931 23613 11940 23647
rect 11888 23604 11940 23613
rect 13728 23604 13780 23656
rect 15752 23647 15804 23656
rect 15752 23613 15761 23647
rect 15761 23613 15795 23647
rect 15795 23613 15804 23647
rect 15752 23604 15804 23613
rect 19064 23672 19116 23724
rect 19340 23715 19392 23724
rect 19340 23681 19349 23715
rect 19349 23681 19383 23715
rect 19383 23681 19392 23715
rect 19340 23672 19392 23681
rect 21272 23672 21324 23724
rect 22376 23672 22428 23724
rect 16028 23604 16080 23656
rect 19616 23647 19668 23656
rect 19616 23613 19625 23647
rect 19625 23613 19659 23647
rect 19659 23613 19668 23647
rect 19616 23604 19668 23613
rect 20628 23604 20680 23656
rect 22192 23604 22244 23656
rect 16580 23536 16632 23588
rect 7472 23468 7524 23520
rect 13360 23468 13412 23520
rect 16396 23468 16448 23520
rect 23296 23604 23348 23656
rect 23296 23468 23348 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 4436 23307 4488 23316
rect 4436 23273 4445 23307
rect 4445 23273 4479 23307
rect 4479 23273 4488 23307
rect 4436 23264 4488 23273
rect 15200 23264 15252 23316
rect 16764 23264 16816 23316
rect 18696 23264 18748 23316
rect 19616 23264 19668 23316
rect 3424 23196 3476 23248
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 2780 23128 2832 23137
rect 3424 23103 3476 23112
rect 3424 23069 3433 23103
rect 3433 23069 3467 23103
rect 3467 23069 3476 23103
rect 3424 23060 3476 23069
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7656 23128 7708 23180
rect 9680 23196 9732 23248
rect 10324 23196 10376 23248
rect 8392 23171 8444 23180
rect 8392 23137 8401 23171
rect 8401 23137 8435 23171
rect 8435 23137 8444 23171
rect 8392 23128 8444 23137
rect 10232 23171 10284 23180
rect 10232 23137 10241 23171
rect 10241 23137 10275 23171
rect 10275 23137 10284 23171
rect 10232 23128 10284 23137
rect 11336 23128 11388 23180
rect 9772 23060 9824 23112
rect 2780 22992 2832 23044
rect 3516 22992 3568 23044
rect 4436 22924 4488 22976
rect 5816 22967 5868 22976
rect 5816 22933 5825 22967
rect 5825 22933 5859 22967
rect 5859 22933 5868 22967
rect 5816 22924 5868 22933
rect 7472 22992 7524 23044
rect 12532 23035 12584 23044
rect 12532 23001 12541 23035
rect 12541 23001 12575 23035
rect 12575 23001 12584 23035
rect 12532 22992 12584 23001
rect 7840 22924 7892 22976
rect 8484 22924 8536 22976
rect 9588 22967 9640 22976
rect 9588 22933 9597 22967
rect 9597 22933 9631 22967
rect 9631 22933 9640 22967
rect 9588 22924 9640 22933
rect 10508 22924 10560 22976
rect 11060 22924 11112 22976
rect 13820 23128 13872 23180
rect 14556 23171 14608 23180
rect 14556 23137 14565 23171
rect 14565 23137 14599 23171
rect 14599 23137 14608 23171
rect 14556 23128 14608 23137
rect 17408 23196 17460 23248
rect 21088 23196 21140 23248
rect 17776 23128 17828 23180
rect 22744 23196 22796 23248
rect 21732 23171 21784 23180
rect 21732 23137 21741 23171
rect 21741 23137 21775 23171
rect 21775 23137 21784 23171
rect 21732 23128 21784 23137
rect 13728 23060 13780 23112
rect 18604 23060 18656 23112
rect 20812 23060 20864 23112
rect 21548 23060 21600 23112
rect 23388 23060 23440 23112
rect 24124 23060 24176 23112
rect 17500 22992 17552 23044
rect 19064 22992 19116 23044
rect 15844 22924 15896 22976
rect 16212 22924 16264 22976
rect 16764 22967 16816 22976
rect 16764 22933 16773 22967
rect 16773 22933 16807 22967
rect 16807 22933 16816 22967
rect 16764 22924 16816 22933
rect 18696 22924 18748 22976
rect 18880 22924 18932 22976
rect 20352 22967 20404 22976
rect 20352 22933 20361 22967
rect 20361 22933 20395 22967
rect 20395 22933 20404 22967
rect 20352 22924 20404 22933
rect 22192 22967 22244 22976
rect 22192 22933 22201 22967
rect 22201 22933 22235 22967
rect 22235 22933 22244 22967
rect 22192 22924 22244 22933
rect 25228 22967 25280 22976
rect 25228 22933 25237 22967
rect 25237 22933 25271 22967
rect 25271 22933 25280 22967
rect 25228 22924 25280 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 3516 22720 3568 22772
rect 5816 22720 5868 22772
rect 8852 22720 8904 22772
rect 10508 22763 10560 22772
rect 10508 22729 10517 22763
rect 10517 22729 10551 22763
rect 10551 22729 10560 22763
rect 10508 22720 10560 22729
rect 11520 22720 11572 22772
rect 8392 22652 8444 22704
rect 4436 22584 4488 22636
rect 4528 22584 4580 22636
rect 5540 22584 5592 22636
rect 8852 22584 8904 22636
rect 7656 22516 7708 22568
rect 8208 22516 8260 22568
rect 10784 22448 10836 22500
rect 4252 22380 4304 22432
rect 6276 22380 6328 22432
rect 11336 22380 11388 22432
rect 12532 22720 12584 22772
rect 13912 22720 13964 22772
rect 13360 22652 13412 22704
rect 14464 22652 14516 22704
rect 15016 22652 15068 22704
rect 15200 22652 15252 22704
rect 17960 22720 18012 22772
rect 19432 22763 19484 22772
rect 19432 22729 19441 22763
rect 19441 22729 19475 22763
rect 19475 22729 19484 22763
rect 19432 22720 19484 22729
rect 20536 22720 20588 22772
rect 15844 22584 15896 22636
rect 12808 22559 12860 22568
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 19340 22652 19392 22704
rect 20076 22652 20128 22704
rect 20352 22652 20404 22704
rect 22008 22652 22060 22704
rect 24124 22652 24176 22704
rect 17132 22584 17184 22636
rect 19064 22584 19116 22636
rect 20996 22584 21048 22636
rect 21088 22584 21140 22636
rect 18696 22516 18748 22568
rect 23848 22559 23900 22568
rect 23848 22525 23857 22559
rect 23857 22525 23891 22559
rect 23891 22525 23900 22559
rect 23848 22516 23900 22525
rect 12532 22423 12584 22432
rect 12532 22389 12541 22423
rect 12541 22389 12575 22423
rect 12575 22389 12584 22423
rect 12532 22380 12584 22389
rect 12716 22380 12768 22432
rect 14464 22380 14516 22432
rect 15108 22380 15160 22432
rect 16672 22380 16724 22432
rect 20628 22448 20680 22500
rect 23296 22380 23348 22432
rect 24768 22516 24820 22568
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 4620 22219 4672 22228
rect 4620 22185 4650 22219
rect 4650 22185 4672 22219
rect 4620 22176 4672 22185
rect 15200 22176 15252 22228
rect 19432 22176 19484 22228
rect 20352 22176 20404 22228
rect 23848 22176 23900 22228
rect 12532 22108 12584 22160
rect 5356 22040 5408 22092
rect 7012 22040 7064 22092
rect 7104 22083 7156 22092
rect 7104 22049 7113 22083
rect 7113 22049 7147 22083
rect 7147 22049 7156 22083
rect 7104 22040 7156 22049
rect 11428 22040 11480 22092
rect 12808 22040 12860 22092
rect 13728 22108 13780 22160
rect 9220 21972 9272 22024
rect 15016 22108 15068 22160
rect 15844 22151 15896 22160
rect 15844 22117 15853 22151
rect 15853 22117 15887 22151
rect 15887 22117 15896 22151
rect 15844 22108 15896 22117
rect 14648 22040 14700 22092
rect 17960 22108 18012 22160
rect 18328 22108 18380 22160
rect 18696 22108 18748 22160
rect 19248 22108 19300 22160
rect 18420 22040 18472 22092
rect 18604 22040 18656 22092
rect 23204 22040 23256 22092
rect 14372 21972 14424 22024
rect 15660 22015 15712 22024
rect 15660 21981 15669 22015
rect 15669 21981 15703 22015
rect 15703 21981 15712 22015
rect 15660 21972 15712 21981
rect 16764 22015 16816 22024
rect 16764 21981 16773 22015
rect 16773 21981 16807 22015
rect 16807 21981 16816 22015
rect 16764 21972 16816 21981
rect 6368 21904 6420 21956
rect 7472 21904 7524 21956
rect 8484 21904 8536 21956
rect 10784 21947 10836 21956
rect 10784 21913 10793 21947
rect 10793 21913 10827 21947
rect 10827 21913 10836 21947
rect 10784 21904 10836 21913
rect 11796 21904 11848 21956
rect 6276 21836 6328 21888
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 6920 21879 6972 21888
rect 6920 21845 6929 21879
rect 6929 21845 6963 21879
rect 6963 21845 6972 21879
rect 6920 21836 6972 21845
rect 7012 21879 7064 21888
rect 7012 21845 7021 21879
rect 7021 21845 7055 21879
rect 7055 21845 7064 21879
rect 7012 21836 7064 21845
rect 8576 21836 8628 21888
rect 9588 21836 9640 21888
rect 12440 21879 12492 21888
rect 12440 21845 12449 21879
rect 12449 21845 12483 21879
rect 12483 21845 12492 21879
rect 12440 21836 12492 21845
rect 12716 21836 12768 21888
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 13636 21904 13688 21956
rect 15292 21904 15344 21956
rect 13820 21836 13872 21888
rect 16488 21904 16540 21956
rect 16672 21879 16724 21888
rect 16672 21845 16681 21879
rect 16681 21845 16715 21879
rect 16715 21845 16724 21879
rect 16672 21836 16724 21845
rect 19432 21972 19484 22024
rect 24952 21972 25004 22024
rect 20720 21904 20772 21956
rect 21548 21947 21600 21956
rect 21548 21913 21557 21947
rect 21557 21913 21591 21947
rect 21591 21913 21600 21947
rect 21548 21904 21600 21913
rect 17316 21836 17368 21888
rect 18328 21836 18380 21888
rect 19064 21836 19116 21888
rect 19432 21836 19484 21888
rect 20904 21836 20956 21888
rect 22008 21904 22060 21956
rect 22836 21904 22888 21956
rect 24308 21904 24360 21956
rect 22376 21836 22428 21888
rect 23572 21836 23624 21888
rect 24124 21879 24176 21888
rect 24124 21845 24133 21879
rect 24133 21845 24167 21879
rect 24167 21845 24176 21879
rect 24124 21836 24176 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 6368 21675 6420 21684
rect 6368 21641 6377 21675
rect 6377 21641 6411 21675
rect 6411 21641 6420 21675
rect 6368 21632 6420 21641
rect 6920 21632 6972 21684
rect 7840 21632 7892 21684
rect 10324 21632 10376 21684
rect 3332 21564 3384 21616
rect 8300 21564 8352 21616
rect 4252 21539 4304 21548
rect 4252 21505 4261 21539
rect 4261 21505 4295 21539
rect 4295 21505 4304 21539
rect 4252 21496 4304 21505
rect 2872 21471 2924 21480
rect 2872 21437 2881 21471
rect 2881 21437 2915 21471
rect 2915 21437 2924 21471
rect 2872 21428 2924 21437
rect 4068 21471 4120 21480
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 9036 21496 9088 21548
rect 8208 21428 8260 21480
rect 9588 21564 9640 21616
rect 8576 21360 8628 21412
rect 1676 21292 1728 21344
rect 10140 21428 10192 21480
rect 11152 21564 11204 21616
rect 11796 21632 11848 21684
rect 15200 21632 15252 21684
rect 16856 21632 16908 21684
rect 18420 21632 18472 21684
rect 11612 21496 11664 21548
rect 12440 21564 12492 21616
rect 13268 21564 13320 21616
rect 13912 21564 13964 21616
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 11428 21360 11480 21412
rect 14464 21496 14516 21548
rect 17500 21564 17552 21616
rect 19432 21632 19484 21684
rect 19708 21632 19760 21684
rect 20904 21632 20956 21684
rect 22192 21632 22244 21684
rect 22560 21632 22612 21684
rect 20260 21564 20312 21616
rect 22836 21564 22888 21616
rect 23480 21607 23532 21616
rect 23480 21573 23489 21607
rect 23489 21573 23523 21607
rect 23523 21573 23532 21607
rect 23480 21564 23532 21573
rect 23572 21564 23624 21616
rect 13268 21360 13320 21412
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 10416 21335 10468 21344
rect 10416 21301 10425 21335
rect 10425 21301 10459 21335
rect 10459 21301 10468 21335
rect 10416 21292 10468 21301
rect 11612 21335 11664 21344
rect 11612 21301 11621 21335
rect 11621 21301 11655 21335
rect 11655 21301 11664 21335
rect 11612 21292 11664 21301
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 12440 21335 12492 21344
rect 12440 21301 12449 21335
rect 12449 21301 12483 21335
rect 12483 21301 12492 21335
rect 12440 21292 12492 21301
rect 13360 21292 13412 21344
rect 14740 21471 14792 21480
rect 14740 21437 14749 21471
rect 14749 21437 14783 21471
rect 14783 21437 14792 21471
rect 14740 21428 14792 21437
rect 13912 21360 13964 21412
rect 15292 21496 15344 21548
rect 15752 21471 15804 21480
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 18328 21496 18380 21548
rect 20076 21539 20128 21548
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 20536 21539 20588 21548
rect 20536 21505 20545 21539
rect 20545 21505 20579 21539
rect 20579 21505 20588 21539
rect 20536 21496 20588 21505
rect 22652 21496 22704 21548
rect 23204 21539 23256 21548
rect 23204 21505 23213 21539
rect 23213 21505 23247 21539
rect 23247 21505 23256 21539
rect 23204 21496 23256 21505
rect 17960 21471 18012 21480
rect 17960 21437 17969 21471
rect 17969 21437 18003 21471
rect 18003 21437 18012 21471
rect 17960 21428 18012 21437
rect 18604 21428 18656 21480
rect 13820 21335 13872 21344
rect 13820 21301 13829 21335
rect 13829 21301 13863 21335
rect 13863 21301 13872 21335
rect 13820 21292 13872 21301
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 14004 21292 14056 21301
rect 14280 21335 14332 21344
rect 14280 21301 14289 21335
rect 14289 21301 14323 21335
rect 14323 21301 14332 21335
rect 14280 21292 14332 21301
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 17500 21292 17552 21344
rect 17868 21292 17920 21344
rect 19248 21292 19300 21344
rect 21640 21292 21692 21344
rect 24952 21335 25004 21344
rect 24952 21301 24961 21335
rect 24961 21301 24995 21335
rect 24995 21301 25004 21335
rect 24952 21292 25004 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 7104 21131 7156 21140
rect 7104 21097 7113 21131
rect 7113 21097 7147 21131
rect 7147 21097 7156 21131
rect 7104 21088 7156 21097
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 9312 21088 9364 21140
rect 1308 20952 1360 21004
rect 5356 20995 5408 21004
rect 5356 20961 5365 20995
rect 5365 20961 5399 20995
rect 5399 20961 5408 20995
rect 5356 20952 5408 20961
rect 8392 20952 8444 21004
rect 9772 20952 9824 21004
rect 10140 20952 10192 21004
rect 10416 20952 10468 21004
rect 11612 21088 11664 21140
rect 15292 21088 15344 21140
rect 15752 21088 15804 21140
rect 15936 21020 15988 21072
rect 12440 20952 12492 21004
rect 12808 20952 12860 21004
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 7104 20884 7156 20936
rect 8576 20884 8628 20936
rect 8944 20884 8996 20936
rect 9312 20884 9364 20936
rect 5632 20859 5684 20868
rect 5632 20825 5641 20859
rect 5641 20825 5675 20859
rect 5675 20825 5684 20859
rect 5632 20816 5684 20825
rect 6368 20816 6420 20868
rect 8484 20816 8536 20868
rect 7840 20748 7892 20800
rect 8668 20748 8720 20800
rect 8944 20748 8996 20800
rect 9588 20748 9640 20800
rect 11244 20884 11296 20936
rect 12624 20884 12676 20936
rect 18512 21088 18564 21140
rect 22008 21088 22060 21140
rect 23572 21088 23624 21140
rect 19524 21020 19576 21072
rect 17960 20995 18012 21004
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 18788 20995 18840 21004
rect 18788 20961 18797 20995
rect 18797 20961 18831 20995
rect 18831 20961 18840 20995
rect 18788 20952 18840 20961
rect 20812 20952 20864 21004
rect 22652 20952 22704 21004
rect 24860 20952 24912 21004
rect 24492 20884 24544 20936
rect 14464 20816 14516 20868
rect 16856 20816 16908 20868
rect 19708 20816 19760 20868
rect 20168 20816 20220 20868
rect 25228 20816 25280 20868
rect 10968 20748 11020 20800
rect 11704 20791 11756 20800
rect 11704 20757 11713 20791
rect 11713 20757 11747 20791
rect 11747 20757 11756 20791
rect 11704 20748 11756 20757
rect 12532 20748 12584 20800
rect 13820 20748 13872 20800
rect 16948 20748 17000 20800
rect 17132 20791 17184 20800
rect 17132 20757 17141 20791
rect 17141 20757 17175 20791
rect 17175 20757 17184 20791
rect 17132 20748 17184 20757
rect 19340 20748 19392 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 3424 20544 3476 20596
rect 4344 20587 4396 20596
rect 4344 20553 4353 20587
rect 4353 20553 4387 20587
rect 4387 20553 4396 20587
rect 4344 20544 4396 20553
rect 8852 20587 8904 20596
rect 8852 20553 8861 20587
rect 8861 20553 8895 20587
rect 8895 20553 8904 20587
rect 8852 20544 8904 20553
rect 10324 20544 10376 20596
rect 11060 20544 11112 20596
rect 11704 20544 11756 20596
rect 14464 20544 14516 20596
rect 14740 20544 14792 20596
rect 16488 20544 16540 20596
rect 19524 20587 19576 20596
rect 19524 20553 19533 20587
rect 19533 20553 19567 20587
rect 19567 20553 19576 20587
rect 19524 20544 19576 20553
rect 21548 20544 21600 20596
rect 6368 20476 6420 20528
rect 11980 20476 12032 20528
rect 6736 20408 6788 20460
rect 8392 20408 8444 20460
rect 8944 20408 8996 20460
rect 14096 20476 14148 20528
rect 6000 20340 6052 20392
rect 9128 20340 9180 20392
rect 9312 20383 9364 20392
rect 9312 20349 9321 20383
rect 9321 20349 9355 20383
rect 9355 20349 9364 20383
rect 9312 20340 9364 20349
rect 10876 20383 10928 20392
rect 10876 20349 10885 20383
rect 10885 20349 10919 20383
rect 10919 20349 10928 20383
rect 10876 20340 10928 20349
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 9680 20272 9732 20324
rect 14556 20408 14608 20460
rect 18512 20476 18564 20528
rect 19984 20476 20036 20528
rect 15016 20340 15068 20392
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 18788 20408 18840 20460
rect 22284 20451 22336 20460
rect 22284 20417 22293 20451
rect 22293 20417 22327 20451
rect 22327 20417 22336 20451
rect 22284 20408 22336 20417
rect 24860 20408 24912 20460
rect 25136 20451 25188 20460
rect 25136 20417 25145 20451
rect 25145 20417 25179 20451
rect 25179 20417 25188 20451
rect 25136 20408 25188 20417
rect 15752 20272 15804 20324
rect 18604 20315 18656 20324
rect 18604 20281 18613 20315
rect 18613 20281 18647 20315
rect 18647 20281 18656 20315
rect 18604 20272 18656 20281
rect 19340 20383 19392 20392
rect 19340 20349 19349 20383
rect 19349 20349 19383 20383
rect 19383 20349 19392 20383
rect 19340 20340 19392 20349
rect 24768 20383 24820 20392
rect 24768 20349 24777 20383
rect 24777 20349 24811 20383
rect 24811 20349 24820 20383
rect 24768 20340 24820 20349
rect 21272 20272 21324 20324
rect 6920 20204 6972 20256
rect 10508 20204 10560 20256
rect 10600 20204 10652 20256
rect 14740 20247 14792 20256
rect 14740 20213 14749 20247
rect 14749 20213 14783 20247
rect 14783 20213 14792 20247
rect 14740 20204 14792 20213
rect 16948 20204 17000 20256
rect 17684 20204 17736 20256
rect 19616 20204 19668 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 5632 20000 5684 20052
rect 7012 20000 7064 20052
rect 9036 20000 9088 20052
rect 5172 19932 5224 19984
rect 11704 20000 11756 20052
rect 14648 20000 14700 20052
rect 20996 20000 21048 20052
rect 23572 20000 23624 20052
rect 11244 19932 11296 19984
rect 8208 19864 8260 19916
rect 10232 19864 10284 19916
rect 16488 19932 16540 19984
rect 18880 19932 18932 19984
rect 15108 19864 15160 19916
rect 18328 19864 18380 19916
rect 6920 19796 6972 19848
rect 10508 19796 10560 19848
rect 12716 19796 12768 19848
rect 16580 19796 16632 19848
rect 19800 19864 19852 19916
rect 24860 19864 24912 19916
rect 19156 19796 19208 19848
rect 21916 19796 21968 19848
rect 23756 19796 23808 19848
rect 24400 19796 24452 19848
rect 7656 19660 7708 19712
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 10508 19703 10560 19712
rect 10508 19669 10517 19703
rect 10517 19669 10551 19703
rect 10551 19669 10560 19703
rect 10508 19660 10560 19669
rect 13544 19728 13596 19780
rect 15108 19728 15160 19780
rect 17132 19728 17184 19780
rect 17868 19728 17920 19780
rect 22376 19728 22428 19780
rect 12256 19660 12308 19712
rect 12716 19660 12768 19712
rect 13452 19703 13504 19712
rect 13452 19669 13461 19703
rect 13461 19669 13495 19703
rect 13495 19669 13504 19703
rect 13452 19660 13504 19669
rect 18788 19660 18840 19712
rect 22652 19660 22704 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 4068 19456 4120 19508
rect 7748 19456 7800 19508
rect 10140 19456 10192 19508
rect 10876 19456 10928 19508
rect 15200 19456 15252 19508
rect 2780 19388 2832 19440
rect 8484 19388 8536 19440
rect 11980 19388 12032 19440
rect 12716 19388 12768 19440
rect 13452 19388 13504 19440
rect 5540 19252 5592 19304
rect 7564 19363 7616 19372
rect 7564 19329 7573 19363
rect 7573 19329 7607 19363
rect 7607 19329 7616 19363
rect 7564 19320 7616 19329
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 10692 19320 10744 19372
rect 14464 19320 14516 19372
rect 15108 19388 15160 19440
rect 18972 19456 19024 19508
rect 19064 19388 19116 19440
rect 20168 19388 20220 19440
rect 23572 19388 23624 19440
rect 24124 19388 24176 19440
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 9404 19252 9456 19304
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12348 19295 12400 19304
rect 12348 19261 12357 19295
rect 12357 19261 12391 19295
rect 12391 19261 12400 19295
rect 12348 19252 12400 19261
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 16672 19320 16724 19372
rect 17408 19320 17460 19372
rect 24400 19320 24452 19372
rect 16120 19252 16172 19304
rect 1768 19184 1820 19236
rect 21088 19252 21140 19304
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 21456 19184 21508 19236
rect 7104 19116 7156 19168
rect 11612 19116 11664 19168
rect 16488 19116 16540 19168
rect 18696 19116 18748 19168
rect 20444 19116 20496 19168
rect 23756 19159 23808 19168
rect 23756 19125 23765 19159
rect 23765 19125 23799 19159
rect 23799 19125 23808 19159
rect 23756 19116 23808 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 6000 18955 6052 18964
rect 6000 18921 6009 18955
rect 6009 18921 6043 18955
rect 6043 18921 6052 18955
rect 6000 18912 6052 18921
rect 9128 18955 9180 18964
rect 9128 18921 9137 18955
rect 9137 18921 9171 18955
rect 9171 18921 9180 18955
rect 9128 18912 9180 18921
rect 10508 18912 10560 18964
rect 11428 18955 11480 18964
rect 11428 18921 11437 18955
rect 11437 18921 11471 18955
rect 11471 18921 11480 18955
rect 11428 18912 11480 18921
rect 15200 18912 15252 18964
rect 16488 18912 16540 18964
rect 16672 18955 16724 18964
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 19432 18912 19484 18964
rect 6276 18844 6328 18896
rect 1308 18776 1360 18828
rect 6644 18819 6696 18828
rect 6644 18785 6653 18819
rect 6653 18785 6687 18819
rect 6687 18785 6696 18819
rect 6644 18776 6696 18785
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 10692 18844 10744 18896
rect 13636 18844 13688 18896
rect 16212 18844 16264 18896
rect 19892 18844 19944 18896
rect 20352 18912 20404 18964
rect 22284 18955 22336 18964
rect 22284 18921 22293 18955
rect 22293 18921 22327 18955
rect 22327 18921 22336 18955
rect 22284 18912 22336 18921
rect 10508 18776 10560 18828
rect 11060 18776 11112 18828
rect 12348 18776 12400 18828
rect 14648 18776 14700 18828
rect 7288 18640 7340 18692
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 10232 18708 10284 18760
rect 8852 18640 8904 18692
rect 9496 18640 9548 18692
rect 11152 18640 11204 18692
rect 12072 18640 12124 18692
rect 14740 18708 14792 18760
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 17224 18776 17276 18828
rect 19708 18776 19760 18828
rect 21088 18776 21140 18828
rect 24032 18819 24084 18828
rect 24032 18785 24041 18819
rect 24041 18785 24075 18819
rect 24075 18785 24084 18819
rect 24032 18776 24084 18785
rect 16396 18708 16448 18760
rect 16672 18708 16724 18760
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 19800 18708 19852 18760
rect 24584 18751 24636 18760
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 12532 18640 12584 18692
rect 13360 18640 13412 18692
rect 20076 18640 20128 18692
rect 23480 18640 23532 18692
rect 7104 18572 7156 18624
rect 10140 18572 10192 18624
rect 10324 18572 10376 18624
rect 11888 18615 11940 18624
rect 11888 18581 11897 18615
rect 11897 18581 11931 18615
rect 11931 18581 11940 18615
rect 11888 18572 11940 18581
rect 14004 18572 14056 18624
rect 15936 18615 15988 18624
rect 15936 18581 15945 18615
rect 15945 18581 15979 18615
rect 15979 18581 15988 18615
rect 15936 18572 15988 18581
rect 19432 18572 19484 18624
rect 19984 18572 20036 18624
rect 20168 18615 20220 18624
rect 20168 18581 20177 18615
rect 20177 18581 20211 18615
rect 20211 18581 20220 18615
rect 20168 18572 20220 18581
rect 21180 18572 21232 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 8576 18368 8628 18420
rect 9036 18368 9088 18420
rect 9772 18368 9824 18420
rect 10876 18368 10928 18420
rect 11152 18411 11204 18420
rect 11152 18377 11161 18411
rect 11161 18377 11195 18411
rect 11195 18377 11204 18411
rect 11152 18368 11204 18377
rect 12072 18368 12124 18420
rect 13820 18368 13872 18420
rect 14648 18368 14700 18420
rect 14740 18411 14792 18420
rect 14740 18377 14749 18411
rect 14749 18377 14783 18411
rect 14783 18377 14792 18411
rect 14740 18368 14792 18377
rect 19340 18368 19392 18420
rect 19984 18368 20036 18420
rect 20904 18368 20956 18420
rect 14280 18300 14332 18352
rect 8484 18232 8536 18284
rect 9496 18232 9548 18284
rect 10968 18232 11020 18284
rect 6552 18207 6604 18216
rect 6552 18173 6561 18207
rect 6561 18173 6595 18207
rect 6595 18173 6604 18207
rect 6552 18164 6604 18173
rect 7472 18164 7524 18216
rect 9864 18164 9916 18216
rect 10508 18164 10560 18216
rect 11152 18164 11204 18216
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 15936 18232 15988 18284
rect 18328 18300 18380 18352
rect 20352 18300 20404 18352
rect 19432 18232 19484 18284
rect 20536 18232 20588 18284
rect 13636 18164 13688 18216
rect 14188 18164 14240 18216
rect 17960 18164 18012 18216
rect 21088 18164 21140 18216
rect 23756 18300 23808 18352
rect 25136 18343 25188 18352
rect 25136 18309 25145 18343
rect 25145 18309 25179 18343
rect 25179 18309 25188 18343
rect 25136 18300 25188 18309
rect 22744 18232 22796 18284
rect 9404 18028 9456 18080
rect 20628 18096 20680 18148
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 23480 18139 23532 18148
rect 23480 18105 23489 18139
rect 23489 18105 23523 18139
rect 23523 18105 23532 18139
rect 23480 18096 23532 18105
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 11980 18028 12032 18080
rect 13912 18028 13964 18080
rect 19800 18071 19852 18080
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 23296 18028 23348 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 5816 17824 5868 17876
rect 6644 17824 6696 17876
rect 7288 17867 7340 17876
rect 7288 17833 7297 17867
rect 7297 17833 7331 17867
rect 7331 17833 7340 17867
rect 7288 17824 7340 17833
rect 12072 17824 12124 17876
rect 17960 17824 18012 17876
rect 23572 17867 23624 17876
rect 23572 17833 23581 17867
rect 23581 17833 23615 17867
rect 23615 17833 23624 17867
rect 23572 17824 23624 17833
rect 24584 17824 24636 17876
rect 10324 17756 10376 17808
rect 12256 17756 12308 17808
rect 14648 17756 14700 17808
rect 6552 17688 6604 17740
rect 6460 17620 6512 17672
rect 7748 17731 7800 17740
rect 7748 17697 7757 17731
rect 7757 17697 7791 17731
rect 7791 17697 7800 17731
rect 7748 17688 7800 17697
rect 7840 17731 7892 17740
rect 7840 17697 7849 17731
rect 7849 17697 7883 17731
rect 7883 17697 7892 17731
rect 7840 17688 7892 17697
rect 12440 17688 12492 17740
rect 14464 17688 14516 17740
rect 14740 17731 14792 17740
rect 14740 17697 14749 17731
rect 14749 17697 14783 17731
rect 14783 17697 14792 17731
rect 14740 17688 14792 17697
rect 14924 17756 14976 17808
rect 18788 17756 18840 17808
rect 24124 17799 24176 17808
rect 24124 17765 24133 17799
rect 24133 17765 24167 17799
rect 24167 17765 24176 17799
rect 24124 17756 24176 17765
rect 7564 17620 7616 17672
rect 8300 17620 8352 17672
rect 11796 17663 11848 17672
rect 5356 17595 5408 17604
rect 5356 17561 5365 17595
rect 5365 17561 5399 17595
rect 5399 17561 5408 17595
rect 5356 17552 5408 17561
rect 11796 17629 11805 17663
rect 11805 17629 11839 17663
rect 11839 17629 11848 17663
rect 11796 17620 11848 17629
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 11152 17552 11204 17604
rect 13636 17552 13688 17604
rect 16764 17620 16816 17672
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 17132 17620 17184 17672
rect 17316 17620 17368 17672
rect 18328 17620 18380 17672
rect 21088 17688 21140 17740
rect 23756 17620 23808 17672
rect 7656 17527 7708 17536
rect 7656 17493 7665 17527
rect 7665 17493 7699 17527
rect 7699 17493 7708 17527
rect 7656 17484 7708 17493
rect 8484 17484 8536 17536
rect 8944 17484 8996 17536
rect 10508 17484 10560 17536
rect 12624 17484 12676 17536
rect 20628 17552 20680 17604
rect 21180 17552 21232 17604
rect 22100 17595 22152 17604
rect 22100 17561 22109 17595
rect 22109 17561 22143 17595
rect 22143 17561 22152 17595
rect 22100 17552 22152 17561
rect 14924 17484 14976 17536
rect 15200 17484 15252 17536
rect 16672 17484 16724 17536
rect 17868 17484 17920 17536
rect 19432 17484 19484 17536
rect 19708 17484 19760 17536
rect 22468 17484 22520 17536
rect 25228 17527 25280 17536
rect 25228 17493 25237 17527
rect 25237 17493 25271 17527
rect 25271 17493 25280 17527
rect 25228 17484 25280 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 5356 17323 5408 17332
rect 5356 17289 5365 17323
rect 5365 17289 5399 17323
rect 5399 17289 5408 17323
rect 5356 17280 5408 17289
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 7656 17280 7708 17332
rect 9588 17280 9640 17332
rect 9864 17280 9916 17332
rect 10968 17280 11020 17332
rect 11428 17280 11480 17332
rect 4068 17212 4120 17264
rect 11612 17212 11664 17264
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6644 17144 6696 17196
rect 10048 17144 10100 17196
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 8576 17119 8628 17128
rect 8576 17085 8585 17119
rect 8585 17085 8619 17119
rect 8619 17085 8628 17119
rect 8576 17076 8628 17085
rect 9404 17076 9456 17128
rect 10508 17076 10560 17128
rect 8484 17008 8536 17060
rect 9312 17008 9364 17060
rect 2780 16940 2832 16992
rect 6460 16940 6512 16992
rect 6644 16940 6696 16992
rect 7748 16940 7800 16992
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 12808 17323 12860 17332
rect 12808 17289 12817 17323
rect 12817 17289 12851 17323
rect 12851 17289 12860 17323
rect 12808 17280 12860 17289
rect 13820 17280 13872 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 16856 17323 16908 17332
rect 16856 17289 16865 17323
rect 16865 17289 16899 17323
rect 16899 17289 16908 17323
rect 16856 17280 16908 17289
rect 13544 17212 13596 17264
rect 18420 17280 18472 17332
rect 18972 17280 19024 17332
rect 21456 17323 21508 17332
rect 21456 17289 21465 17323
rect 21465 17289 21499 17323
rect 21499 17289 21508 17323
rect 21456 17280 21508 17289
rect 22100 17280 22152 17332
rect 17868 17212 17920 17264
rect 18696 17212 18748 17264
rect 19708 17212 19760 17264
rect 12624 17076 12676 17128
rect 13728 17076 13780 17128
rect 13820 17076 13872 17128
rect 19248 17144 19300 17196
rect 20720 17144 20772 17196
rect 25136 17255 25188 17264
rect 25136 17221 25145 17255
rect 25145 17221 25179 17255
rect 25179 17221 25188 17255
rect 25136 17212 25188 17221
rect 14556 17119 14608 17128
rect 14556 17085 14565 17119
rect 14565 17085 14599 17119
rect 14599 17085 14608 17119
rect 14556 17076 14608 17085
rect 15660 17119 15712 17128
rect 15660 17085 15669 17119
rect 15669 17085 15703 17119
rect 15703 17085 15712 17119
rect 15660 17076 15712 17085
rect 16396 17076 16448 17128
rect 21088 17076 21140 17128
rect 21272 17076 21324 17128
rect 23664 17144 23716 17196
rect 11980 17008 12032 17060
rect 18788 17008 18840 17060
rect 20260 17008 20312 17060
rect 18604 16940 18656 16992
rect 23388 17051 23440 17060
rect 23388 17017 23397 17051
rect 23397 17017 23431 17051
rect 23431 17017 23440 17051
rect 23388 17008 23440 17017
rect 22836 16940 22888 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 6000 16736 6052 16788
rect 7840 16736 7892 16788
rect 8484 16736 8536 16788
rect 16396 16779 16448 16788
rect 16396 16745 16405 16779
rect 16405 16745 16439 16779
rect 16439 16745 16448 16779
rect 16396 16736 16448 16745
rect 18696 16779 18748 16788
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 20628 16736 20680 16788
rect 22468 16736 22520 16788
rect 8668 16711 8720 16720
rect 6920 16600 6972 16652
rect 8668 16677 8677 16711
rect 8677 16677 8711 16711
rect 8711 16677 8720 16711
rect 8668 16668 8720 16677
rect 9496 16668 9548 16720
rect 8300 16600 8352 16652
rect 9220 16600 9272 16652
rect 1768 16575 1820 16584
rect 1768 16541 1777 16575
rect 1777 16541 1811 16575
rect 1811 16541 1820 16575
rect 1768 16532 1820 16541
rect 9496 16575 9548 16584
rect 9496 16541 9505 16575
rect 9505 16541 9539 16575
rect 9539 16541 9548 16575
rect 9496 16532 9548 16541
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 12624 16600 12676 16652
rect 13360 16600 13412 16652
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 17592 16600 17644 16652
rect 17868 16600 17920 16652
rect 22192 16600 22244 16652
rect 25228 16736 25280 16788
rect 24032 16668 24084 16720
rect 11520 16532 11572 16584
rect 13452 16532 13504 16584
rect 18512 16532 18564 16584
rect 20812 16532 20864 16584
rect 20996 16532 21048 16584
rect 1308 16464 1360 16516
rect 6920 16464 6972 16516
rect 7656 16507 7708 16516
rect 7656 16473 7665 16507
rect 7665 16473 7699 16507
rect 7699 16473 7708 16507
rect 7656 16464 7708 16473
rect 7564 16396 7616 16448
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 16488 16464 16540 16516
rect 21180 16464 21232 16516
rect 22468 16464 22520 16516
rect 12808 16396 12860 16448
rect 19340 16439 19392 16448
rect 19340 16405 19349 16439
rect 19349 16405 19383 16439
rect 19383 16405 19392 16439
rect 19340 16396 19392 16405
rect 19984 16396 20036 16448
rect 20812 16396 20864 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 6736 16192 6788 16244
rect 7748 16235 7800 16244
rect 7748 16201 7757 16235
rect 7757 16201 7791 16235
rect 7791 16201 7800 16235
rect 7748 16192 7800 16201
rect 10692 16235 10744 16244
rect 10692 16201 10701 16235
rect 10701 16201 10735 16235
rect 10735 16201 10744 16235
rect 10692 16192 10744 16201
rect 19892 16235 19944 16244
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 20168 16192 20220 16244
rect 11796 16124 11848 16176
rect 15108 16124 15160 16176
rect 17500 16124 17552 16176
rect 20996 16124 21048 16176
rect 7840 16056 7892 16108
rect 8484 15988 8536 16040
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 11704 16056 11756 16108
rect 12348 16099 12400 16108
rect 12348 16065 12357 16099
rect 12357 16065 12391 16099
rect 12391 16065 12400 16099
rect 12348 16056 12400 16065
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 24308 16056 24360 16108
rect 8852 15963 8904 15972
rect 8852 15929 8861 15963
rect 8861 15929 8895 15963
rect 8895 15929 8904 15963
rect 8852 15920 8904 15929
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 11612 15988 11664 16040
rect 18420 15988 18472 16040
rect 19156 16031 19208 16040
rect 19156 15997 19165 16031
rect 19165 15997 19199 16031
rect 19199 15997 19208 16031
rect 19156 15988 19208 15997
rect 19800 16031 19852 16040
rect 19800 15997 19809 16031
rect 19809 15997 19843 16031
rect 19843 15997 19852 16031
rect 19800 15988 19852 15997
rect 12808 15920 12860 15972
rect 14096 15920 14148 15972
rect 21456 15988 21508 16040
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 23572 15920 23624 15972
rect 10048 15852 10100 15904
rect 16488 15852 16540 15904
rect 17592 15852 17644 15904
rect 18696 15895 18748 15904
rect 18696 15861 18705 15895
rect 18705 15861 18739 15895
rect 18739 15861 18748 15895
rect 18696 15852 18748 15861
rect 21364 15852 21416 15904
rect 22652 15852 22704 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 7656 15648 7708 15700
rect 8392 15648 8444 15700
rect 14556 15648 14608 15700
rect 7288 15444 7340 15496
rect 8576 15580 8628 15632
rect 10876 15580 10928 15632
rect 11704 15512 11756 15564
rect 12440 15512 12492 15564
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 17224 15648 17276 15700
rect 18512 15648 18564 15700
rect 20904 15648 20956 15700
rect 22284 15648 22336 15700
rect 9404 15444 9456 15496
rect 10600 15444 10652 15496
rect 14556 15444 14608 15496
rect 7012 15308 7064 15360
rect 7564 15308 7616 15360
rect 11060 15308 11112 15360
rect 11244 15351 11296 15360
rect 11244 15317 11253 15351
rect 11253 15317 11287 15351
rect 11287 15317 11296 15351
rect 11244 15308 11296 15317
rect 11704 15351 11756 15360
rect 11704 15317 11713 15351
rect 11713 15317 11747 15351
rect 11747 15317 11756 15351
rect 11704 15308 11756 15317
rect 15016 15376 15068 15428
rect 15108 15419 15160 15428
rect 15108 15385 15117 15419
rect 15117 15385 15151 15419
rect 15151 15385 15160 15419
rect 15108 15376 15160 15385
rect 14556 15308 14608 15360
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 17592 15444 17644 15496
rect 18788 15512 18840 15564
rect 20812 15555 20864 15564
rect 20812 15521 20821 15555
rect 20821 15521 20855 15555
rect 20855 15521 20864 15555
rect 20812 15512 20864 15521
rect 21180 15512 21232 15564
rect 18328 15444 18380 15496
rect 18696 15444 18748 15496
rect 19156 15444 19208 15496
rect 21548 15444 21600 15496
rect 22744 15487 22796 15496
rect 22744 15453 22753 15487
rect 22753 15453 22787 15487
rect 22787 15453 22796 15487
rect 22744 15444 22796 15453
rect 16212 15419 16264 15428
rect 16212 15385 16221 15419
rect 16221 15385 16255 15419
rect 16255 15385 16264 15419
rect 16212 15376 16264 15385
rect 19340 15376 19392 15428
rect 25504 15376 25556 15428
rect 18696 15308 18748 15360
rect 19524 15308 19576 15360
rect 20996 15351 21048 15360
rect 20996 15317 21005 15351
rect 21005 15317 21039 15351
rect 21039 15317 21048 15351
rect 20996 15308 21048 15317
rect 21732 15308 21784 15360
rect 21916 15308 21968 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 6828 15104 6880 15156
rect 7012 15079 7064 15088
rect 7012 15045 7021 15079
rect 7021 15045 7055 15079
rect 7055 15045 7064 15079
rect 7012 15036 7064 15045
rect 11888 15104 11940 15156
rect 14096 15147 14148 15156
rect 14096 15113 14105 15147
rect 14105 15113 14139 15147
rect 14139 15113 14148 15147
rect 14096 15104 14148 15113
rect 16212 15104 16264 15156
rect 17500 15147 17552 15156
rect 10784 15036 10836 15088
rect 12440 15036 12492 15088
rect 12716 15036 12768 15088
rect 13452 15036 13504 15088
rect 15016 15079 15068 15088
rect 15016 15045 15025 15079
rect 15025 15045 15059 15079
rect 15059 15045 15068 15079
rect 15016 15036 15068 15045
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 18420 15104 18472 15156
rect 19064 15104 19116 15156
rect 11520 14968 11572 15020
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 7104 14900 7156 14952
rect 7656 14900 7708 14952
rect 11152 14943 11204 14952
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 12348 14900 12400 14952
rect 14188 14943 14240 14952
rect 14188 14909 14197 14943
rect 14197 14909 14231 14943
rect 14231 14909 14240 14943
rect 14188 14900 14240 14909
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 16672 14900 16724 14952
rect 17224 14900 17276 14952
rect 18512 15036 18564 15088
rect 19800 15036 19852 15088
rect 20720 15104 20772 15156
rect 21824 15104 21876 15156
rect 24400 15104 24452 15156
rect 18328 14968 18380 15020
rect 21640 14968 21692 15020
rect 22376 15036 22428 15088
rect 18604 14900 18656 14952
rect 19432 14900 19484 14952
rect 19800 14900 19852 14952
rect 21824 14943 21876 14952
rect 21824 14909 21833 14943
rect 21833 14909 21867 14943
rect 21867 14909 21876 14943
rect 21824 14900 21876 14909
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 14832 14875 14884 14884
rect 14832 14841 14841 14875
rect 14841 14841 14875 14875
rect 14875 14841 14884 14875
rect 14832 14832 14884 14841
rect 16580 14832 16632 14884
rect 8300 14764 8352 14816
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 9680 14764 9732 14816
rect 15568 14764 15620 14816
rect 18696 14832 18748 14884
rect 21180 14832 21232 14884
rect 23848 14832 23900 14884
rect 20628 14764 20680 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 7288 14560 7340 14612
rect 7656 14560 7708 14612
rect 11244 14560 11296 14612
rect 12624 14560 12676 14612
rect 15660 14560 15712 14612
rect 16304 14560 16356 14612
rect 20996 14560 21048 14612
rect 8300 14424 8352 14476
rect 11152 14424 11204 14476
rect 6276 14288 6328 14340
rect 6828 14288 6880 14340
rect 10048 14288 10100 14340
rect 10140 14331 10192 14340
rect 10140 14297 10149 14331
rect 10149 14297 10183 14331
rect 10183 14297 10192 14331
rect 10140 14288 10192 14297
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 13728 14492 13780 14544
rect 18696 14492 18748 14544
rect 16028 14424 16080 14476
rect 17408 14424 17460 14476
rect 18328 14424 18380 14476
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 14648 14356 14700 14408
rect 14004 14288 14056 14340
rect 8944 14220 8996 14229
rect 11888 14220 11940 14272
rect 15568 14356 15620 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 22836 14356 22888 14408
rect 16488 14288 16540 14340
rect 22376 14288 22428 14340
rect 23940 14288 23992 14340
rect 16396 14220 16448 14272
rect 19708 14220 19760 14272
rect 22836 14263 22888 14272
rect 22836 14229 22845 14263
rect 22845 14229 22879 14263
rect 22879 14229 22888 14263
rect 22836 14220 22888 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 6828 14016 6880 14068
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 8300 13948 8352 14000
rect 8944 14016 8996 14068
rect 11244 14016 11296 14068
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12808 14016 12860 14068
rect 14740 14016 14792 14068
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 19524 14016 19576 14068
rect 22008 14016 22060 14068
rect 10784 13948 10836 14000
rect 15292 13948 15344 14000
rect 15752 13991 15804 14000
rect 15752 13957 15761 13991
rect 15761 13957 15795 13991
rect 15795 13957 15804 13991
rect 15752 13948 15804 13957
rect 17868 13991 17920 14000
rect 17868 13957 17877 13991
rect 17877 13957 17911 13991
rect 17911 13957 17920 13991
rect 17868 13948 17920 13957
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 13360 13880 13412 13932
rect 14280 13880 14332 13932
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 18788 13923 18840 13932
rect 18788 13889 18797 13923
rect 18797 13889 18831 13923
rect 18831 13889 18840 13923
rect 18788 13880 18840 13889
rect 22100 13880 22152 13932
rect 22836 13923 22888 13932
rect 22836 13889 22845 13923
rect 22845 13889 22879 13923
rect 22879 13889 22888 13923
rect 22836 13880 22888 13889
rect 23480 13880 23532 13932
rect 940 13812 992 13864
rect 8208 13855 8260 13864
rect 8208 13821 8217 13855
rect 8217 13821 8251 13855
rect 8251 13821 8260 13855
rect 8208 13812 8260 13821
rect 8760 13812 8812 13864
rect 8944 13812 8996 13864
rect 9404 13744 9456 13796
rect 11704 13744 11756 13796
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 15568 13812 15620 13864
rect 15844 13812 15896 13864
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 18328 13812 18380 13864
rect 14648 13744 14700 13796
rect 19340 13744 19392 13796
rect 21456 13812 21508 13864
rect 20720 13744 20772 13796
rect 10508 13676 10560 13728
rect 14740 13719 14792 13728
rect 14740 13685 14749 13719
rect 14749 13685 14783 13719
rect 14783 13685 14792 13719
rect 14740 13676 14792 13685
rect 16120 13676 16172 13728
rect 19524 13676 19576 13728
rect 19800 13676 19852 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 8208 13472 8260 13524
rect 11060 13472 11112 13524
rect 8484 13268 8536 13320
rect 14372 13472 14424 13524
rect 17776 13472 17828 13524
rect 20996 13472 21048 13524
rect 15384 13404 15436 13456
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 12900 13379 12952 13388
rect 12900 13345 12909 13379
rect 12909 13345 12943 13379
rect 12943 13345 12952 13379
rect 12900 13336 12952 13345
rect 13728 13336 13780 13388
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 14924 13336 14976 13388
rect 14004 13268 14056 13320
rect 14648 13268 14700 13320
rect 17408 13404 17460 13456
rect 17316 13336 17368 13388
rect 17500 13268 17552 13320
rect 20720 13268 20772 13320
rect 20904 13268 20956 13320
rect 22376 13336 22428 13388
rect 22192 13268 22244 13320
rect 19156 13200 19208 13252
rect 16488 13132 16540 13184
rect 20352 13243 20404 13252
rect 20352 13209 20361 13243
rect 20361 13209 20395 13243
rect 20395 13209 20404 13243
rect 20352 13200 20404 13209
rect 20996 13200 21048 13252
rect 25504 13200 25556 13252
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 11244 12971 11296 12980
rect 11244 12937 11253 12971
rect 11253 12937 11287 12971
rect 11287 12937 11296 12971
rect 11244 12928 11296 12937
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 13360 12928 13412 12980
rect 15200 12928 15252 12980
rect 15476 12928 15528 12980
rect 17132 12928 17184 12980
rect 18788 12928 18840 12980
rect 21732 12928 21784 12980
rect 14648 12860 14700 12912
rect 15568 12903 15620 12912
rect 15568 12869 15577 12903
rect 15577 12869 15611 12903
rect 15611 12869 15620 12903
rect 15568 12860 15620 12869
rect 19524 12860 19576 12912
rect 14372 12792 14424 12844
rect 16396 12792 16448 12844
rect 24216 12860 24268 12912
rect 24584 12860 24636 12912
rect 20996 12835 21048 12844
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 22376 12835 22428 12844
rect 22376 12801 22385 12835
rect 22385 12801 22419 12835
rect 22419 12801 22428 12835
rect 22376 12792 22428 12801
rect 23296 12792 23348 12844
rect 23388 12792 23440 12844
rect 10784 12724 10836 12776
rect 15568 12724 15620 12776
rect 17776 12724 17828 12776
rect 12808 12699 12860 12708
rect 12808 12665 12817 12699
rect 12817 12665 12851 12699
rect 12851 12665 12860 12699
rect 12808 12656 12860 12665
rect 16856 12656 16908 12708
rect 13452 12631 13504 12640
rect 13452 12597 13461 12631
rect 13461 12597 13495 12631
rect 13495 12597 13504 12631
rect 13452 12588 13504 12597
rect 13728 12588 13780 12640
rect 18052 12656 18104 12708
rect 21088 12724 21140 12776
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22100 12724 22152 12733
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 20996 12656 21048 12708
rect 21364 12656 21416 12708
rect 22836 12656 22888 12708
rect 20444 12588 20496 12640
rect 23296 12588 23348 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 16028 12427 16080 12436
rect 16028 12393 16037 12427
rect 16037 12393 16071 12427
rect 16071 12393 16080 12427
rect 16028 12384 16080 12393
rect 2780 12316 2832 12368
rect 5908 12316 5960 12368
rect 8300 12248 8352 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 11244 12248 11296 12300
rect 10600 12044 10652 12096
rect 12164 12248 12216 12300
rect 20076 12316 20128 12368
rect 25044 12316 25096 12368
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 21364 12248 21416 12300
rect 22376 12248 22428 12300
rect 22652 12248 22704 12300
rect 12256 12180 12308 12232
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 15660 12180 15712 12232
rect 16488 12180 16540 12232
rect 18880 12180 18932 12232
rect 21732 12180 21784 12232
rect 17316 12112 17368 12164
rect 20904 12112 20956 12164
rect 21456 12112 21508 12164
rect 11244 12044 11296 12096
rect 19524 12044 19576 12096
rect 24860 12044 24912 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 9864 11840 9916 11892
rect 11980 11840 12032 11892
rect 7840 11704 7892 11756
rect 11060 11704 11112 11756
rect 11428 11704 11480 11756
rect 14280 11840 14332 11892
rect 19708 11840 19760 11892
rect 20996 11883 21048 11892
rect 20996 11849 21005 11883
rect 21005 11849 21039 11883
rect 21039 11849 21048 11883
rect 20996 11840 21048 11849
rect 15660 11772 15712 11824
rect 16948 11772 17000 11824
rect 10600 11679 10652 11688
rect 10600 11645 10609 11679
rect 10609 11645 10643 11679
rect 10643 11645 10652 11679
rect 10600 11636 10652 11645
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 13912 11636 13964 11688
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 18880 11772 18932 11824
rect 20536 11772 20588 11824
rect 22100 11815 22152 11824
rect 22100 11781 22109 11815
rect 22109 11781 22143 11815
rect 22143 11781 22152 11815
rect 22100 11772 22152 11781
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 17500 11704 17552 11756
rect 19892 11704 19944 11756
rect 21180 11704 21232 11756
rect 23848 11704 23900 11756
rect 19432 11636 19484 11688
rect 16488 11568 16540 11620
rect 22560 11568 22612 11620
rect 23388 11568 23440 11620
rect 13544 11500 13596 11552
rect 13728 11500 13780 11552
rect 15200 11500 15252 11552
rect 19892 11543 19944 11552
rect 19892 11509 19901 11543
rect 19901 11509 19935 11543
rect 19935 11509 19944 11543
rect 19892 11500 19944 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 12440 11296 12492 11348
rect 12992 11296 13044 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 15292 11296 15344 11348
rect 19064 11296 19116 11348
rect 19432 11339 19484 11348
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 12532 11228 12584 11280
rect 12164 11160 12216 11212
rect 12716 11160 12768 11212
rect 20628 11228 20680 11280
rect 15660 11160 15712 11212
rect 20812 11160 20864 11212
rect 19064 11092 19116 11144
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 20536 11092 20588 11144
rect 11244 11024 11296 11076
rect 12256 11024 12308 11076
rect 12992 11024 13044 11076
rect 14280 11067 14332 11076
rect 14280 11033 14289 11067
rect 14289 11033 14323 11067
rect 14323 11033 14332 11067
rect 14280 11024 14332 11033
rect 15568 10956 15620 11008
rect 16120 11024 16172 11076
rect 19616 11024 19668 11076
rect 21272 11024 21324 11076
rect 21548 11067 21600 11076
rect 21548 11033 21557 11067
rect 21557 11033 21591 11067
rect 21591 11033 21600 11067
rect 21548 11024 21600 11033
rect 16396 10999 16448 11008
rect 16396 10965 16405 10999
rect 16405 10965 16439 10999
rect 16439 10965 16448 10999
rect 16396 10956 16448 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 9956 10752 10008 10804
rect 12992 10752 13044 10804
rect 11980 10548 12032 10600
rect 15568 10752 15620 10804
rect 15200 10684 15252 10736
rect 16396 10684 16448 10736
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 15384 10548 15436 10600
rect 13544 10480 13596 10532
rect 19892 10616 19944 10668
rect 20444 10659 20496 10668
rect 20444 10625 20453 10659
rect 20453 10625 20487 10659
rect 20487 10625 20496 10659
rect 20444 10616 20496 10625
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 23940 10480 23992 10532
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 19892 10412 19944 10464
rect 21456 10412 21508 10464
rect 23480 10455 23532 10464
rect 23480 10421 23489 10455
rect 23489 10421 23523 10455
rect 23523 10421 23532 10455
rect 23480 10412 23532 10421
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 18972 10004 19024 10056
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 22836 10047 22888 10056
rect 22836 10013 22845 10047
rect 22845 10013 22879 10047
rect 22879 10013 22888 10047
rect 22836 10004 22888 10013
rect 24952 10004 25004 10056
rect 17040 9979 17092 9988
rect 17040 9945 17049 9979
rect 17049 9945 17083 9979
rect 17083 9945 17092 9979
rect 17040 9936 17092 9945
rect 22928 9936 22980 9988
rect 22192 9911 22244 9920
rect 22192 9877 22201 9911
rect 22201 9877 22235 9911
rect 22235 9877 22244 9911
rect 22192 9868 22244 9877
rect 23204 9868 23256 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 22836 9707 22888 9716
rect 22836 9673 22845 9707
rect 22845 9673 22879 9707
rect 22879 9673 22888 9707
rect 22836 9664 22888 9673
rect 12624 9596 12676 9648
rect 13452 9528 13504 9580
rect 13728 9528 13780 9580
rect 19892 9528 19944 9580
rect 23296 9571 23348 9580
rect 23296 9537 23305 9571
rect 23305 9537 23339 9571
rect 23339 9537 23348 9571
rect 23296 9528 23348 9537
rect 23940 9571 23992 9580
rect 23940 9537 23949 9571
rect 23949 9537 23983 9571
rect 23983 9537 23992 9571
rect 23940 9528 23992 9537
rect 2872 9460 2924 9512
rect 5724 9460 5776 9512
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 19432 9324 19484 9376
rect 24584 9324 24636 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 16764 8916 16816 8968
rect 20352 8916 20404 8968
rect 23388 8916 23440 8968
rect 25044 8916 25096 8968
rect 21824 8848 21876 8900
rect 7748 8780 7800 8832
rect 17776 8780 17828 8832
rect 23940 8823 23992 8832
rect 23940 8789 23949 8823
rect 23949 8789 23983 8823
rect 23983 8789 23992 8823
rect 23940 8780 23992 8789
rect 24032 8780 24084 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 7840 8576 7892 8628
rect 21916 8508 21968 8560
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 5540 8440 5592 8492
rect 11520 8372 11572 8424
rect 11888 8372 11940 8424
rect 23480 8440 23532 8492
rect 22652 8415 22704 8424
rect 22652 8381 22661 8415
rect 22661 8381 22695 8415
rect 22695 8381 22704 8415
rect 22652 8372 22704 8381
rect 20996 8304 21048 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 8300 7896 8352 7948
rect 23296 7939 23348 7948
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 21456 7828 21508 7880
rect 21640 7828 21692 7880
rect 24860 7871 24912 7880
rect 24860 7837 24869 7871
rect 24869 7837 24903 7871
rect 24903 7837 24912 7871
rect 24860 7828 24912 7837
rect 4252 7803 4304 7812
rect 4252 7769 4261 7803
rect 4261 7769 4295 7803
rect 4295 7769 4304 7803
rect 4252 7760 4304 7769
rect 8576 7760 8628 7812
rect 15936 7760 15988 7812
rect 22008 7760 22060 7812
rect 21732 7735 21784 7744
rect 21732 7701 21741 7735
rect 21741 7701 21775 7735
rect 21775 7701 21784 7735
rect 21732 7692 21784 7701
rect 24124 7692 24176 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 4252 7488 4304 7540
rect 15476 7420 15528 7472
rect 23388 7420 23440 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 20628 7395 20680 7404
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 23388 7284 23440 7336
rect 16304 7216 16356 7268
rect 20260 7148 20312 7200
rect 20352 7148 20404 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 24860 6808 24912 6860
rect 17224 6740 17276 6792
rect 3148 6604 3200 6656
rect 6184 6604 6236 6656
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 24584 6740 24636 6792
rect 21916 6715 21968 6724
rect 21916 6681 21925 6715
rect 21925 6681 21959 6715
rect 21959 6681 21968 6715
rect 21916 6672 21968 6681
rect 21456 6604 21508 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 3976 6400 4028 6452
rect 21640 6400 21692 6452
rect 19708 6332 19760 6384
rect 2780 6264 2832 6316
rect 21456 6307 21508 6316
rect 21456 6273 21465 6307
rect 21465 6273 21499 6307
rect 21499 6273 21508 6307
rect 21456 6264 21508 6273
rect 22008 6264 22060 6316
rect 23940 6307 23992 6316
rect 23940 6273 23949 6307
rect 23949 6273 23983 6307
rect 23983 6273 23992 6307
rect 23940 6264 23992 6273
rect 22284 6196 22336 6248
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 22836 6128 22888 6180
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 21916 5720 21968 5772
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 21548 5652 21600 5704
rect 22192 5652 22244 5704
rect 21364 5627 21416 5636
rect 21364 5593 21373 5627
rect 21373 5593 21407 5627
rect 21407 5593 21416 5627
rect 21364 5584 21416 5593
rect 23020 5584 23072 5636
rect 19984 5516 20036 5568
rect 21456 5516 21508 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 2780 5312 2832 5364
rect 1676 5176 1728 5228
rect 3976 5176 4028 5228
rect 23020 5244 23072 5296
rect 20996 5219 21048 5228
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 21824 5176 21876 5228
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 5540 5040 5592 5092
rect 19708 5108 19760 5160
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 21824 5040 21876 5092
rect 1676 4972 1728 5024
rect 9496 4972 9548 5024
rect 13360 4972 13412 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 9128 4700 9180 4752
rect 8300 4632 8352 4684
rect 13452 4632 13504 4684
rect 13636 4632 13688 4684
rect 22100 4700 22152 4752
rect 2504 4564 2556 4616
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 21732 4564 21784 4616
rect 20352 4539 20404 4548
rect 20352 4505 20361 4539
rect 20361 4505 20395 4539
rect 20395 4505 20404 4539
rect 20352 4496 20404 4505
rect 2044 4428 2096 4480
rect 20076 4428 20128 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 1400 4088 1452 4140
rect 7564 4088 7616 4140
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 3424 4020 3476 4072
rect 3884 4020 3936 4072
rect 7472 4020 7524 4072
rect 10416 4020 10468 4072
rect 11612 4020 11664 4072
rect 13452 4020 13504 4072
rect 15844 4020 15896 4072
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 20260 4088 20312 4140
rect 22192 4131 22244 4140
rect 22192 4097 22201 4131
rect 22201 4097 22235 4131
rect 22235 4097 22244 4131
rect 22192 4088 22244 4097
rect 4804 3952 4856 4004
rect 9588 3952 9640 4004
rect 16396 3952 16448 4004
rect 17500 4020 17552 4072
rect 20444 4020 20496 4072
rect 21548 3952 21600 4004
rect 2688 3884 2740 3936
rect 4068 3884 4120 3936
rect 4252 3884 4304 3936
rect 6092 3884 6144 3936
rect 6736 3884 6788 3936
rect 8760 3884 8812 3936
rect 9404 3884 9456 3936
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 10968 3884 11020 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 8944 3680 8996 3732
rect 9220 3723 9272 3732
rect 9220 3689 9229 3723
rect 9229 3689 9263 3723
rect 9263 3689 9272 3723
rect 9220 3680 9272 3689
rect 10048 3723 10100 3732
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 22652 3680 22704 3732
rect 24952 3680 25004 3732
rect 5264 3655 5316 3664
rect 5264 3621 5273 3655
rect 5273 3621 5307 3655
rect 5307 3621 5316 3655
rect 5264 3612 5316 3621
rect 16120 3612 16172 3664
rect 7472 3544 7524 3596
rect 8300 3544 8352 3596
rect 14648 3544 14700 3596
rect 16028 3544 16080 3596
rect 17868 3544 17920 3596
rect 2412 3519 2464 3528
rect 2412 3485 2421 3519
rect 2421 3485 2455 3519
rect 2455 3485 2464 3519
rect 2412 3476 2464 3485
rect 3516 3476 3568 3528
rect 2780 3408 2832 3460
rect 6092 3476 6144 3528
rect 6460 3476 6512 3528
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 9772 3476 9824 3528
rect 10876 3476 10928 3528
rect 14188 3476 14240 3528
rect 16580 3476 16632 3528
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 18328 3476 18380 3528
rect 20812 3476 20864 3528
rect 12716 3451 12768 3460
rect 12716 3417 12725 3451
rect 12725 3417 12759 3451
rect 12759 3417 12768 3451
rect 12716 3408 12768 3417
rect 14924 3408 14976 3460
rect 18972 3408 19024 3460
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3332 3340 3384 3349
rect 4988 3340 5040 3392
rect 6828 3340 6880 3392
rect 7840 3340 7892 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 11244 3340 11296 3392
rect 22008 3340 22060 3392
rect 23388 3340 23440 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 2412 3136 2464 3188
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 7380 3136 7432 3188
rect 8392 3179 8444 3188
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 11060 3136 11112 3188
rect 19340 3136 19392 3188
rect 7196 3068 7248 3120
rect 9588 3068 9640 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 3884 3000 3936 3052
rect 5356 3000 5408 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8300 3000 8352 3052
rect 8668 3000 8720 3052
rect 9036 3000 9088 3052
rect 10508 3000 10560 3052
rect 10968 3000 11020 3052
rect 11244 3000 11296 3052
rect 14832 3068 14884 3120
rect 18604 3068 18656 3120
rect 20352 3068 20404 3120
rect 21456 3068 21508 3120
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 16488 3000 16540 3052
rect 17684 3000 17736 3052
rect 18512 3000 18564 3052
rect 4160 2932 4212 2984
rect 9496 2932 9548 2984
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 14188 2932 14240 2984
rect 15660 2932 15712 2984
rect 18328 2932 18380 2984
rect 20720 3000 20772 3052
rect 22560 3000 22612 3052
rect 13912 2864 13964 2916
rect 17132 2864 17184 2916
rect 21180 2932 21232 2984
rect 22468 2932 22520 2984
rect 21364 2864 21416 2916
rect 22652 2864 22704 2916
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 11336 2796 11388 2848
rect 16764 2796 16816 2848
rect 19892 2796 19944 2848
rect 20812 2796 20864 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 2872 2592 2924 2644
rect 4068 2635 4120 2644
rect 4068 2601 4077 2635
rect 4077 2601 4111 2635
rect 4111 2601 4120 2635
rect 4068 2592 4120 2601
rect 14464 2592 14516 2644
rect 18512 2635 18564 2644
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 24676 2635 24728 2644
rect 24676 2601 24685 2635
rect 24685 2601 24719 2635
rect 24719 2601 24728 2635
rect 24676 2592 24728 2601
rect 10600 2456 10652 2508
rect 13636 2524 13688 2576
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 4620 2388 4672 2440
rect 7196 2388 7248 2440
rect 7564 2388 7616 2440
rect 8944 2388 8996 2440
rect 10140 2388 10192 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 11980 2456 12032 2508
rect 14556 2456 14608 2508
rect 15292 2456 15344 2508
rect 17776 2456 17828 2508
rect 12072 2388 12124 2440
rect 12808 2388 12860 2440
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 20720 2456 20772 2508
rect 25044 2388 25096 2440
rect 5724 2320 5776 2372
rect 13820 2320 13872 2372
rect 24124 2320 24176 2372
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 12256 2252 12308 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 8944 2048 8996 2100
rect 13912 2048 13964 2100
rect 12256 1980 12308 2032
rect 17316 1980 17368 2032
rect 7104 1912 7156 1964
rect 13728 1912 13780 1964
rect 11152 1844 11204 1896
rect 12348 1844 12400 1896
<< metal2 >>
rect 1490 56200 1546 57000
rect 1858 56200 1914 57000
rect 2226 56200 2282 57000
rect 2594 56200 2650 57000
rect 2962 56200 3018 57000
rect 3330 56200 3386 57000
rect 3698 56200 3754 57000
rect 4066 56200 4122 57000
rect 4434 56200 4490 57000
rect 4802 56200 4858 57000
rect 5170 56200 5226 57000
rect 5276 56222 5488 56250
rect 1504 49298 1532 56200
rect 1584 52896 1636 52902
rect 1584 52838 1636 52844
rect 1596 50930 1624 52838
rect 1584 50924 1636 50930
rect 1584 50866 1636 50872
rect 1872 49910 1900 56200
rect 2240 50386 2268 56200
rect 2412 53440 2464 53446
rect 2412 53382 2464 53388
rect 2424 53106 2452 53382
rect 2412 53100 2464 53106
rect 2412 53042 2464 53048
rect 2608 52986 2636 56200
rect 2976 55214 3004 56200
rect 2884 55186 3004 55214
rect 2608 52958 2820 52986
rect 2792 50998 2820 52958
rect 2884 51474 2912 55186
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2962 53000 3018 53009
rect 2962 52935 2964 52944
rect 3016 52935 3018 52944
rect 2964 52906 3016 52912
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 3344 52086 3372 56200
rect 3712 52698 3740 56200
rect 3974 55448 4030 55457
rect 3974 55383 4030 55392
rect 3988 55214 4016 55383
rect 3896 55186 4016 55214
rect 3700 52692 3752 52698
rect 3700 52634 3752 52640
rect 3424 52488 3476 52494
rect 3424 52430 3476 52436
rect 3332 52080 3384 52086
rect 3332 52022 3384 52028
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2872 51468 2924 51474
rect 2872 51410 2924 51416
rect 3436 51066 3464 52430
rect 3896 52086 3924 55186
rect 3976 54120 4028 54126
rect 3976 54062 4028 54068
rect 3988 53786 4016 54062
rect 3976 53780 4028 53786
rect 3976 53722 4028 53728
rect 4080 52986 4108 56200
rect 4252 53100 4304 53106
rect 4252 53042 4304 53048
rect 4080 52958 4200 52986
rect 3884 52080 3936 52086
rect 3884 52022 3936 52028
rect 3976 51264 4028 51270
rect 3976 51206 4028 51212
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 2780 50992 2832 50998
rect 2780 50934 2832 50940
rect 3700 50924 3752 50930
rect 3700 50866 3752 50872
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 3330 50416 3386 50425
rect 2228 50380 2280 50386
rect 3330 50351 3386 50360
rect 2228 50322 2280 50328
rect 1860 49904 1912 49910
rect 1860 49846 1912 49852
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 1492 49292 1544 49298
rect 1492 49234 1544 49240
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 1308 43308 1360 43314
rect 1308 43250 1360 43256
rect 1320 43217 1348 43250
rect 1306 43208 1362 43217
rect 1306 43143 1362 43152
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 3344 41414 3372 50351
rect 3424 49836 3476 49842
rect 3424 49778 3476 49784
rect 3436 42294 3464 49778
rect 3516 49088 3568 49094
rect 3516 49030 3568 49036
rect 3528 43110 3556 49030
rect 3516 43104 3568 43110
rect 3516 43046 3568 43052
rect 3424 42288 3476 42294
rect 3424 42230 3476 42236
rect 3712 41750 3740 50866
rect 3988 50318 4016 51206
rect 4172 50998 4200 52958
rect 4264 52698 4292 53042
rect 4448 53038 4476 56200
rect 4436 53032 4488 53038
rect 4436 52974 4488 52980
rect 4252 52692 4304 52698
rect 4252 52634 4304 52640
rect 4620 52352 4672 52358
rect 4620 52294 4672 52300
rect 4632 51406 4660 52294
rect 4816 52086 4844 56200
rect 5184 56114 5212 56200
rect 5276 56114 5304 56222
rect 5184 56086 5304 56114
rect 5460 53428 5488 56222
rect 5538 56200 5594 57000
rect 5906 56200 5962 57000
rect 6274 56200 6330 57000
rect 6642 56200 6698 57000
rect 7010 56200 7066 57000
rect 7378 56200 7434 57000
rect 7746 56200 7802 57000
rect 7852 56222 8064 56250
rect 5552 53582 5580 56200
rect 5632 54188 5684 54194
rect 5632 54130 5684 54136
rect 5540 53576 5592 53582
rect 5540 53518 5592 53524
rect 5460 53400 5580 53428
rect 4988 52624 5040 52630
rect 4988 52566 5040 52572
rect 4804 52080 4856 52086
rect 4804 52022 4856 52028
rect 4804 51944 4856 51950
rect 4804 51886 4856 51892
rect 4620 51400 4672 51406
rect 4620 51342 4672 51348
rect 4160 50992 4212 50998
rect 4160 50934 4212 50940
rect 3884 50312 3936 50318
rect 3884 50254 3936 50260
rect 3976 50312 4028 50318
rect 3976 50254 4028 50260
rect 3792 43172 3844 43178
rect 3792 43114 3844 43120
rect 3700 41744 3752 41750
rect 3700 41686 3752 41692
rect 3344 41386 3464 41414
rect 1308 41132 1360 41138
rect 1308 41074 1360 41080
rect 1320 40769 1348 41074
rect 3436 41002 3464 41386
rect 3424 40996 3476 41002
rect 3424 40938 3476 40944
rect 3700 40928 3752 40934
rect 3700 40870 3752 40876
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 1306 40760 1362 40769
rect 2950 40763 3258 40772
rect 1306 40695 1362 40704
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 1308 38344 1360 38350
rect 1306 38312 1308 38321
rect 1360 38312 1362 38321
rect 1306 38247 1362 38256
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1596 35873 1624 36110
rect 1582 35864 1638 35873
rect 1582 35799 1638 35808
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 1216 33516 1268 33522
rect 1216 33458 1268 33464
rect 1228 33425 1256 33458
rect 1214 33416 1270 33425
rect 1214 33351 1270 33360
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 3712 31346 3740 40870
rect 3700 31340 3752 31346
rect 3700 31282 3752 31288
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2778 30968 2834 30977
rect 2950 30971 3258 30980
rect 2778 30903 2834 30912
rect 2792 27538 2820 30903
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 3516 29572 3568 29578
rect 3516 29514 3568 29520
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2870 28520 2926 28529
rect 2870 28455 2926 28464
rect 3424 28484 3476 28490
rect 2780 27532 2832 27538
rect 2780 27474 2832 27480
rect 2778 26072 2834 26081
rect 2778 26007 2834 26016
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 1320 21010 1348 21111
rect 1308 21004 1360 21010
rect 1308 20946 1360 20952
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18737 1348 18770
rect 1688 18766 1716 21286
rect 1780 20942 1808 24006
rect 2792 23186 2820 26007
rect 2884 24750 2912 28455
rect 3424 28426 3476 28432
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 3344 25158 3372 26930
rect 3436 26042 3464 28426
rect 3528 27130 3556 29514
rect 3608 29164 3660 29170
rect 3608 29106 3660 29112
rect 3620 27538 3648 29106
rect 3608 27532 3660 27538
rect 3608 27474 3660 27480
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3620 26926 3648 27474
rect 3804 26994 3832 43114
rect 3896 42294 3924 50254
rect 4252 50176 4304 50182
rect 4252 50118 4304 50124
rect 4264 49910 4292 50118
rect 4252 49904 4304 49910
rect 4252 49846 4304 49852
rect 4066 48104 4122 48113
rect 4066 48039 4122 48048
rect 3974 45656 4030 45665
rect 3974 45591 3976 45600
rect 4028 45591 4030 45600
rect 3976 45562 4028 45568
rect 3884 42288 3936 42294
rect 3884 42230 3936 42236
rect 4080 41274 4108 48039
rect 4816 42770 4844 51886
rect 4804 42764 4856 42770
rect 4804 42706 4856 42712
rect 5000 42362 5028 52566
rect 5552 51474 5580 53400
rect 5540 51468 5592 51474
rect 5540 51410 5592 51416
rect 5540 51332 5592 51338
rect 5540 51274 5592 51280
rect 5552 51066 5580 51274
rect 5540 51060 5592 51066
rect 5540 51002 5592 51008
rect 5448 50924 5500 50930
rect 5448 50866 5500 50872
rect 5460 42770 5488 50866
rect 5644 50386 5672 54130
rect 5920 53786 5948 56200
rect 6000 54188 6052 54194
rect 6000 54130 6052 54136
rect 5908 53780 5960 53786
rect 5908 53722 5960 53728
rect 5632 50380 5684 50386
rect 5632 50322 5684 50328
rect 5908 44872 5960 44878
rect 5908 44814 5960 44820
rect 5448 42764 5500 42770
rect 5448 42706 5500 42712
rect 5264 42560 5316 42566
rect 5264 42502 5316 42508
rect 4988 42356 5040 42362
rect 4988 42298 5040 42304
rect 4344 42220 4396 42226
rect 4344 42162 4396 42168
rect 4356 41818 4384 42162
rect 4896 42152 4948 42158
rect 4896 42094 4948 42100
rect 4344 41812 4396 41818
rect 4344 41754 4396 41760
rect 4068 41268 4120 41274
rect 4068 41210 4120 41216
rect 4068 38208 4120 38214
rect 4068 38150 4120 38156
rect 3884 33312 3936 33318
rect 3884 33254 3936 33260
rect 3896 27538 3924 33254
rect 3976 31272 4028 31278
rect 3976 31214 4028 31220
rect 3988 29306 4016 31214
rect 4080 29714 4108 38150
rect 4160 36032 4212 36038
rect 4160 35974 4212 35980
rect 4068 29708 4120 29714
rect 4068 29650 4120 29656
rect 3976 29300 4028 29306
rect 3976 29242 4028 29248
rect 4172 28626 4200 35974
rect 4356 30326 4384 41754
rect 4528 35624 4580 35630
rect 4528 35566 4580 35572
rect 4540 35290 4568 35566
rect 4528 35284 4580 35290
rect 4528 35226 4580 35232
rect 4908 34746 4936 42094
rect 5080 41540 5132 41546
rect 5080 41482 5132 41488
rect 4896 34740 4948 34746
rect 4896 34682 4948 34688
rect 4896 31272 4948 31278
rect 4896 31214 4948 31220
rect 4344 30320 4396 30326
rect 4344 30262 4396 30268
rect 4160 28620 4212 28626
rect 4160 28562 4212 28568
rect 3884 27532 3936 27538
rect 3884 27474 3936 27480
rect 4252 27396 4304 27402
rect 4252 27338 4304 27344
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 3424 26036 3476 26042
rect 3424 25978 3476 25984
rect 3424 25900 3476 25906
rect 3424 25842 3476 25848
rect 3332 25152 3384 25158
rect 3332 25094 3384 25100
rect 3344 24750 3372 25094
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2870 23624 2926 23633
rect 2870 23559 2926 23568
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 2792 19446 2820 22986
rect 2884 21486 2912 23559
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3344 21622 3372 24686
rect 3436 23254 3464 25842
rect 3620 24206 3648 26862
rect 3804 26586 3832 26930
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 3804 25294 3832 26522
rect 4160 25696 4212 25702
rect 4160 25638 4212 25644
rect 4172 25498 4200 25638
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 3792 25288 3844 25294
rect 3792 25230 3844 25236
rect 4172 24206 4200 25434
rect 3608 24200 3660 24206
rect 3608 24142 3660 24148
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4264 23866 4292 27338
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4436 26784 4488 26790
rect 4436 26726 4488 26732
rect 4448 26382 4476 26726
rect 4436 26376 4488 26382
rect 4436 26318 4488 26324
rect 4448 25498 4476 26318
rect 4436 25492 4488 25498
rect 4436 25434 4488 25440
rect 4436 25288 4488 25294
rect 4436 25230 4488 25236
rect 4344 24676 4396 24682
rect 4344 24618 4396 24624
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 3436 20602 3464 23054
rect 3516 23044 3568 23050
rect 3516 22986 3568 22992
rect 3528 22778 3556 22986
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 4080 21486 4108 23666
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4264 21554 4292 22374
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 4080 19514 4108 21422
rect 4356 20602 4384 24618
rect 4448 23322 4476 25230
rect 4540 24614 4568 27270
rect 4908 26353 4936 31214
rect 5092 29850 5120 41482
rect 5276 31210 5304 42502
rect 5448 39432 5500 39438
rect 5448 39374 5500 39380
rect 5356 39364 5408 39370
rect 5356 39306 5408 39312
rect 5368 39098 5396 39306
rect 5356 39092 5408 39098
rect 5356 39034 5408 39040
rect 5460 38418 5488 39374
rect 5920 39098 5948 44814
rect 6012 44538 6040 54130
rect 6184 53100 6236 53106
rect 6184 53042 6236 53048
rect 6092 50924 6144 50930
rect 6092 50866 6144 50872
rect 6104 45082 6132 50866
rect 6196 46102 6224 53042
rect 6288 53038 6316 56200
rect 6276 53032 6328 53038
rect 6276 52974 6328 52980
rect 6552 52896 6604 52902
rect 6552 52838 6604 52844
rect 6564 52154 6592 52838
rect 6656 52562 6684 56200
rect 6736 53576 6788 53582
rect 6736 53518 6788 53524
rect 6644 52556 6696 52562
rect 6644 52498 6696 52504
rect 6552 52148 6604 52154
rect 6552 52090 6604 52096
rect 6460 52012 6512 52018
rect 6460 51954 6512 51960
rect 6184 46096 6236 46102
rect 6184 46038 6236 46044
rect 6092 45076 6144 45082
rect 6092 45018 6144 45024
rect 6000 44532 6052 44538
rect 6000 44474 6052 44480
rect 6472 44470 6500 51954
rect 6644 51400 6696 51406
rect 6644 51342 6696 51348
rect 6552 45280 6604 45286
rect 6552 45222 6604 45228
rect 6564 44962 6592 45222
rect 6656 45082 6684 51342
rect 6748 50998 6776 53518
rect 6828 52488 6880 52494
rect 6828 52430 6880 52436
rect 6736 50992 6788 50998
rect 6736 50934 6788 50940
rect 6840 46646 6868 52430
rect 7024 51474 7052 56200
rect 7392 53514 7420 56200
rect 7380 53508 7432 53514
rect 7380 53450 7432 53456
rect 7288 53440 7340 53446
rect 7288 53382 7340 53388
rect 7196 53100 7248 53106
rect 7196 53042 7248 53048
rect 7208 52154 7236 53042
rect 7196 52148 7248 52154
rect 7196 52090 7248 52096
rect 7012 51468 7064 51474
rect 7012 51410 7064 51416
rect 6828 46640 6880 46646
rect 6828 46582 6880 46588
rect 6644 45076 6696 45082
rect 6644 45018 6696 45024
rect 7300 45014 7328 53382
rect 7760 52562 7788 56200
rect 7852 54194 7880 56222
rect 8036 56114 8064 56222
rect 8114 56200 8170 57000
rect 8482 56200 8538 57000
rect 8850 56200 8906 57000
rect 9218 56200 9274 57000
rect 9586 56200 9642 57000
rect 9954 56200 10010 57000
rect 10322 56200 10378 57000
rect 10690 56200 10746 57000
rect 11058 56200 11114 57000
rect 11426 56200 11482 57000
rect 11794 56200 11850 57000
rect 12162 56200 12218 57000
rect 12530 56200 12586 57000
rect 12898 56200 12954 57000
rect 13266 56200 13322 57000
rect 13634 56200 13690 57000
rect 14002 56200 14058 57000
rect 14370 56200 14426 57000
rect 14738 56200 14794 57000
rect 15106 56200 15162 57000
rect 15474 56200 15530 57000
rect 15842 56200 15898 57000
rect 16210 56200 16266 57000
rect 16578 56200 16634 57000
rect 16946 56200 17002 57000
rect 17314 56200 17370 57000
rect 17682 56200 17738 57000
rect 18050 56200 18106 57000
rect 18156 56222 18368 56250
rect 8128 56114 8156 56200
rect 8036 56086 8156 56114
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 7840 54188 7892 54194
rect 7840 54130 7892 54136
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 8392 53100 8444 53106
rect 8392 53042 8444 53048
rect 7840 52964 7892 52970
rect 7840 52906 7892 52912
rect 7748 52556 7800 52562
rect 7748 52498 7800 52504
rect 7852 51074 7880 52906
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7576 51046 7880 51074
rect 7472 50312 7524 50318
rect 7472 50254 7524 50260
rect 7484 47258 7512 50254
rect 7472 47252 7524 47258
rect 7472 47194 7524 47200
rect 7380 46368 7432 46374
rect 7380 46310 7432 46316
rect 7288 45008 7340 45014
rect 6564 44934 6684 44962
rect 7288 44950 7340 44956
rect 6656 44810 6684 44934
rect 6644 44804 6696 44810
rect 6644 44746 6696 44752
rect 7288 44804 7340 44810
rect 7288 44746 7340 44752
rect 6460 44464 6512 44470
rect 6460 44406 6512 44412
rect 6368 42560 6420 42566
rect 6368 42502 6420 42508
rect 6380 42265 6408 42502
rect 6366 42256 6422 42265
rect 6366 42191 6422 42200
rect 6184 42016 6236 42022
rect 6184 41958 6236 41964
rect 5908 39092 5960 39098
rect 5908 39034 5960 39040
rect 6000 38956 6052 38962
rect 6000 38898 6052 38904
rect 6092 38956 6144 38962
rect 6092 38898 6144 38904
rect 5448 38412 5500 38418
rect 5448 38354 5500 38360
rect 5460 38010 5488 38354
rect 6012 38010 6040 38898
rect 5448 38004 5500 38010
rect 5448 37946 5500 37952
rect 6000 38004 6052 38010
rect 6000 37946 6052 37952
rect 5540 37800 5592 37806
rect 5540 37742 5592 37748
rect 5552 36242 5580 37742
rect 6000 37324 6052 37330
rect 6000 37266 6052 37272
rect 5540 36236 5592 36242
rect 5540 36178 5592 36184
rect 5552 34474 5580 36178
rect 5908 35760 5960 35766
rect 5908 35702 5960 35708
rect 5920 35086 5948 35702
rect 6012 35630 6040 37266
rect 6000 35624 6052 35630
rect 6000 35566 6052 35572
rect 5908 35080 5960 35086
rect 5908 35022 5960 35028
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5540 34468 5592 34474
rect 5540 34410 5592 34416
rect 5644 34066 5672 34546
rect 5816 34536 5868 34542
rect 5816 34478 5868 34484
rect 5632 34060 5684 34066
rect 5632 34002 5684 34008
rect 5828 32910 5856 34478
rect 6012 33998 6040 35566
rect 6104 34746 6132 38898
rect 6092 34740 6144 34746
rect 6092 34682 6144 34688
rect 6000 33992 6052 33998
rect 6000 33934 6052 33940
rect 6196 33658 6224 41958
rect 6552 41540 6604 41546
rect 6552 41482 6604 41488
rect 6564 41018 6592 41482
rect 6656 41154 6684 44746
rect 6828 44396 6880 44402
rect 6828 44338 6880 44344
rect 6656 41126 6776 41154
rect 6564 40990 6684 41018
rect 6656 40934 6684 40990
rect 6644 40928 6696 40934
rect 6644 40870 6696 40876
rect 6656 39846 6684 40870
rect 6644 39840 6696 39846
rect 6644 39782 6696 39788
rect 6552 38412 6604 38418
rect 6552 38354 6604 38360
rect 6644 38412 6696 38418
rect 6748 38400 6776 41126
rect 6696 38372 6776 38400
rect 6644 38354 6696 38360
rect 6368 38276 6420 38282
rect 6368 38218 6420 38224
rect 6380 37942 6408 38218
rect 6368 37936 6420 37942
rect 6368 37878 6420 37884
rect 6380 36854 6408 37878
rect 6564 37398 6592 38354
rect 6552 37392 6604 37398
rect 6552 37334 6604 37340
rect 6368 36848 6420 36854
rect 6368 36790 6420 36796
rect 6564 36174 6592 37334
rect 6840 36582 6868 44338
rect 7300 44198 7328 44746
rect 7288 44192 7340 44198
rect 7288 44134 7340 44140
rect 7104 40656 7156 40662
rect 7104 40598 7156 40604
rect 7012 38888 7064 38894
rect 7012 38830 7064 38836
rect 6828 36576 6880 36582
rect 6828 36518 6880 36524
rect 7024 36378 7052 38830
rect 7116 37806 7144 40598
rect 7196 40520 7248 40526
rect 7196 40462 7248 40468
rect 7208 39642 7236 40462
rect 7196 39636 7248 39642
rect 7196 39578 7248 39584
rect 7104 37800 7156 37806
rect 7104 37742 7156 37748
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 6552 36168 6604 36174
rect 6552 36110 6604 36116
rect 6564 35834 6592 36110
rect 6920 36100 6972 36106
rect 6920 36042 6972 36048
rect 6932 35834 6960 36042
rect 6552 35828 6604 35834
rect 6552 35770 6604 35776
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 6564 35154 6592 35770
rect 7012 35488 7064 35494
rect 7116 35476 7144 37742
rect 7064 35448 7144 35476
rect 7012 35430 7064 35436
rect 6552 35148 6604 35154
rect 6552 35090 6604 35096
rect 6564 34542 6592 35090
rect 7024 35018 7052 35430
rect 7012 35012 7064 35018
rect 7012 34954 7064 34960
rect 6736 34672 6788 34678
rect 6736 34614 6788 34620
rect 6552 34536 6604 34542
rect 6552 34478 6604 34484
rect 6184 33652 6236 33658
rect 6184 33594 6236 33600
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5828 32434 5856 32846
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 5264 31204 5316 31210
rect 5264 31146 5316 31152
rect 5080 29844 5132 29850
rect 5080 29786 5132 29792
rect 6184 29572 6236 29578
rect 6184 29514 6236 29520
rect 5724 28620 5776 28626
rect 5724 28562 5776 28568
rect 4894 26344 4950 26353
rect 4894 26279 4950 26288
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4448 23066 4476 23258
rect 4448 23038 4568 23066
rect 4436 22976 4488 22982
rect 4436 22918 4488 22924
rect 4448 22642 4476 22918
rect 4540 22642 4568 23038
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 4528 22636 4580 22642
rect 4528 22578 4580 22584
rect 4632 22234 4660 24006
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 1768 19236 1820 19242
rect 1768 19178 1820 19184
rect 1676 18760 1728 18766
rect 1306 18728 1362 18737
rect 1676 18702 1728 18708
rect 1306 18663 1362 18672
rect 1780 16590 1808 19178
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 4080 17270 4108 19450
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 2792 13938 2820 16934
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 940 13864 992 13870
rect 938 13832 940 13841
rect 992 13832 994 13841
rect 938 13767 994 13776
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2792 11393 2820 12310
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2778 11384 2834 11393
rect 2950 11387 3258 11396
rect 2778 11319 2834 11328
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 8945 2912 9454
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2870 8936 2926 8945
rect 2870 8871 2926 8880
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4264 7546 4292 7754
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6497 3188 6598
rect 3146 6488 3202 6497
rect 3988 6458 4016 7346
rect 4908 6914 4936 26279
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5552 26042 5580 26182
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5368 21010 5396 22034
rect 5356 21004 5408 21010
rect 5356 20946 5408 20952
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 4816 6886 4936 6914
rect 3146 6423 3202 6432
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2792 5370 2820 6258
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 1688 5030 1716 5170
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 3398 1440 4082
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 1601 1440 3334
rect 1398 1592 1454 1601
rect 1398 1527 1454 1536
rect 1688 800 1716 4966
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3988 4826 4016 5170
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 3058 1808 3334
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2056 800 2084 4422
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2424 3194 2452 3470
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2516 3074 2544 4558
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 4066 4040 4122 4049
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2424 3046 2544 3074
rect 2424 800 2452 3046
rect 2700 2446 2728 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3330 3496 3386 3505
rect 2780 3460 2832 3466
rect 3330 3431 3386 3440
rect 2780 3402 2832 3408
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2792 800 2820 3402
rect 3344 3398 3372 3431
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2884 2650 2912 2994
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3160 870 3280 898
rect 3160 800 3188 870
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3252 762 3280 870
rect 3436 762 3464 4014
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3528 800 3556 3470
rect 3896 3058 3924 4014
rect 4066 3975 4122 3984
rect 4080 3942 4108 3975
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3896 800 3924 2994
rect 4172 2990 4200 4558
rect 4816 4010 4844 6886
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4066 2680 4122 2689
rect 4066 2615 4068 2624
rect 4120 2615 4122 2624
rect 4068 2586 4120 2592
rect 4264 2446 4292 3878
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4264 800 4292 2382
rect 4632 800 4660 2382
rect 5000 800 5028 3334
rect 5184 3194 5212 19926
rect 5552 19310 5580 22578
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5644 20058 5672 20810
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5368 17338 5396 17546
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5736 9518 5764 28562
rect 5908 27396 5960 27402
rect 5908 27338 5960 27344
rect 5920 26586 5948 27338
rect 6196 26926 6224 29514
rect 6552 27396 6604 27402
rect 6552 27338 6604 27344
rect 6564 27130 6592 27338
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 5908 26580 5960 26586
rect 5908 26522 5960 26528
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5828 25226 5856 25638
rect 5816 25220 5868 25226
rect 5816 25162 5868 25168
rect 5816 22976 5868 22982
rect 5816 22918 5868 22924
rect 5828 22778 5856 22918
rect 5816 22772 5868 22778
rect 5816 22714 5868 22720
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5552 5098 5580 8434
rect 5828 6914 5856 17818
rect 5920 12374 5948 26522
rect 6092 24404 6144 24410
rect 6092 24346 6144 24352
rect 6104 23186 6132 24346
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6012 18970 6040 20334
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6012 16794 6040 17138
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5828 6886 5948 6914
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5264 3664 5316 3670
rect 5262 3632 5264 3641
rect 5316 3632 5318 3641
rect 5262 3567 5318 3576
rect 5920 3194 5948 6886
rect 6196 6662 6224 26862
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6288 24410 6316 25230
rect 6368 25152 6420 25158
rect 6368 25094 6420 25100
rect 6380 24614 6408 25094
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 6276 24404 6328 24410
rect 6276 24346 6328 24352
rect 6380 24138 6408 24550
rect 6368 24132 6420 24138
rect 6368 24074 6420 24080
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6288 21894 6316 22374
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6288 18902 6316 21830
rect 6380 21690 6408 21898
rect 6564 21894 6592 24754
rect 6748 22094 6776 34614
rect 6828 34536 6880 34542
rect 6828 34478 6880 34484
rect 6840 34202 6868 34478
rect 6828 34196 6880 34202
rect 6828 34138 6880 34144
rect 6920 32224 6972 32230
rect 6920 32166 6972 32172
rect 6932 32026 6960 32166
rect 6920 32020 6972 32026
rect 6920 31962 6972 31968
rect 6932 30802 6960 31962
rect 7024 31278 7052 34954
rect 7104 33380 7156 33386
rect 7104 33322 7156 33328
rect 7116 32978 7144 33322
rect 7104 32972 7156 32978
rect 7104 32914 7156 32920
rect 7116 32230 7144 32914
rect 7300 32230 7328 44134
rect 7392 39098 7420 46310
rect 7576 43994 7604 51046
rect 7840 50992 7892 50998
rect 7840 50934 7892 50940
rect 7748 49836 7800 49842
rect 7748 49778 7800 49784
rect 7656 44872 7708 44878
rect 7656 44814 7708 44820
rect 7564 43988 7616 43994
rect 7564 43930 7616 43936
rect 7564 41608 7616 41614
rect 7564 41550 7616 41556
rect 7576 41206 7604 41550
rect 7564 41200 7616 41206
rect 7564 41142 7616 41148
rect 7576 39642 7604 41142
rect 7564 39636 7616 39642
rect 7564 39578 7616 39584
rect 7576 39370 7604 39578
rect 7564 39364 7616 39370
rect 7564 39306 7616 39312
rect 7380 39092 7432 39098
rect 7380 39034 7432 39040
rect 7472 38208 7524 38214
rect 7472 38150 7524 38156
rect 7484 36922 7512 38150
rect 7668 37466 7696 44814
rect 7760 43450 7788 49778
rect 7852 45082 7880 50934
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7840 45076 7892 45082
rect 7840 45018 7892 45024
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 8404 44470 8432 53042
rect 8496 51950 8524 56200
rect 8864 53650 8892 56200
rect 8852 53644 8904 53650
rect 8852 53586 8904 53592
rect 8576 53576 8628 53582
rect 8576 53518 8628 53524
rect 9128 53576 9180 53582
rect 9128 53518 9180 53524
rect 8484 51944 8536 51950
rect 8484 51886 8536 51892
rect 8484 51400 8536 51406
rect 8484 51342 8536 51348
rect 8496 46102 8524 51342
rect 8588 50522 8616 53518
rect 8852 52488 8904 52494
rect 8852 52430 8904 52436
rect 8760 52012 8812 52018
rect 8760 51954 8812 51960
rect 8772 51074 8800 51954
rect 8680 51046 8800 51074
rect 8576 50516 8628 50522
rect 8576 50458 8628 50464
rect 8576 49768 8628 49774
rect 8576 49710 8628 49716
rect 8484 46096 8536 46102
rect 8484 46038 8536 46044
rect 8588 45558 8616 49710
rect 8576 45552 8628 45558
rect 8576 45494 8628 45500
rect 8680 45082 8708 51046
rect 8760 45824 8812 45830
rect 8760 45766 8812 45772
rect 8668 45076 8720 45082
rect 8668 45018 8720 45024
rect 8484 44804 8536 44810
rect 8484 44746 8536 44752
rect 8392 44464 8444 44470
rect 8392 44406 8444 44412
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7748 43444 7800 43450
rect 7748 43386 7800 43392
rect 7840 43308 7892 43314
rect 7840 43250 7892 43256
rect 7748 42560 7800 42566
rect 7748 42502 7800 42508
rect 7760 42158 7788 42502
rect 7748 42152 7800 42158
rect 7748 42094 7800 42100
rect 7852 41414 7880 43250
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 8392 42288 8444 42294
rect 8392 42230 8444 42236
rect 8404 41682 8432 42230
rect 8392 41676 8444 41682
rect 8392 41618 8444 41624
rect 7760 41386 7880 41414
rect 7656 37460 7708 37466
rect 7656 37402 7708 37408
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 7656 36848 7708 36854
rect 7656 36790 7708 36796
rect 7668 36106 7696 36790
rect 7656 36100 7708 36106
rect 7656 36042 7708 36048
rect 7564 35148 7616 35154
rect 7564 35090 7616 35096
rect 7576 33114 7604 35090
rect 7668 34746 7696 36042
rect 7760 35290 7788 41386
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 8404 41070 8432 41618
rect 8116 41064 8168 41070
rect 8116 41006 8168 41012
rect 8392 41064 8444 41070
rect 8392 41006 8444 41012
rect 8128 40730 8156 41006
rect 8116 40724 8168 40730
rect 8116 40666 8168 40672
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 8300 39500 8352 39506
rect 8300 39442 8352 39448
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 8312 38350 8340 39442
rect 8496 38486 8524 44746
rect 8668 43104 8720 43110
rect 8668 43046 8720 43052
rect 8576 42696 8628 42702
rect 8576 42638 8628 42644
rect 8588 41818 8616 42638
rect 8576 41812 8628 41818
rect 8576 41754 8628 41760
rect 8576 39840 8628 39846
rect 8576 39782 8628 39788
rect 8588 38894 8616 39782
rect 8576 38888 8628 38894
rect 8576 38830 8628 38836
rect 8484 38480 8536 38486
rect 8484 38422 8536 38428
rect 8300 38344 8352 38350
rect 8300 38286 8352 38292
rect 8300 38208 8352 38214
rect 8300 38150 8352 38156
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 8312 37942 8340 38150
rect 8300 37936 8352 37942
rect 8300 37878 8352 37884
rect 8496 37244 8524 38422
rect 8680 37874 8708 43046
rect 8772 39386 8800 45766
rect 8864 45014 8892 52430
rect 9140 51882 9168 53518
rect 9232 53038 9260 56200
rect 9600 53564 9628 56200
rect 9968 55214 9996 56200
rect 9876 55186 9996 55214
rect 9876 54126 9904 55186
rect 9956 54188 10008 54194
rect 9956 54130 10008 54136
rect 9864 54120 9916 54126
rect 9864 54062 9916 54068
rect 9600 53536 9720 53564
rect 9496 53100 9548 53106
rect 9496 53042 9548 53048
rect 9220 53032 9272 53038
rect 9220 52974 9272 52980
rect 9312 52420 9364 52426
rect 9312 52362 9364 52368
rect 9128 51876 9180 51882
rect 9128 51818 9180 51824
rect 9036 51400 9088 51406
rect 9036 51342 9088 51348
rect 8944 47048 8996 47054
rect 8944 46990 8996 46996
rect 8852 45008 8904 45014
rect 8852 44950 8904 44956
rect 8956 42566 8984 46990
rect 9048 46714 9076 51342
rect 9220 50924 9272 50930
rect 9220 50866 9272 50872
rect 9232 46714 9260 50866
rect 9324 47802 9352 52362
rect 9404 50312 9456 50318
rect 9404 50254 9456 50260
rect 9312 47796 9364 47802
rect 9312 47738 9364 47744
rect 9036 46708 9088 46714
rect 9036 46650 9088 46656
rect 9220 46708 9272 46714
rect 9220 46650 9272 46656
rect 9128 46572 9180 46578
rect 9128 46514 9180 46520
rect 8944 42560 8996 42566
rect 8944 42502 8996 42508
rect 8852 40996 8904 41002
rect 8852 40938 8904 40944
rect 8864 40458 8892 40938
rect 9036 40588 9088 40594
rect 9036 40530 9088 40536
rect 8852 40452 8904 40458
rect 8852 40394 8904 40400
rect 9048 40390 9076 40530
rect 9036 40384 9088 40390
rect 9036 40326 9088 40332
rect 9048 40118 9076 40326
rect 9036 40112 9088 40118
rect 9036 40054 9088 40060
rect 8772 39358 8892 39386
rect 8760 39296 8812 39302
rect 8760 39238 8812 39244
rect 8772 39098 8800 39238
rect 8760 39092 8812 39098
rect 8760 39034 8812 39040
rect 8864 38978 8892 39358
rect 8772 38950 8892 38978
rect 8668 37868 8720 37874
rect 8668 37810 8720 37816
rect 8576 37800 8628 37806
rect 8772 37754 8800 38950
rect 9048 38826 9076 40054
rect 9140 39642 9168 46514
rect 9312 45552 9364 45558
rect 9312 45494 9364 45500
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9232 44305 9260 44338
rect 9218 44296 9274 44305
rect 9218 44231 9274 44240
rect 9324 43858 9352 45494
rect 9416 43994 9444 50254
rect 9508 49910 9536 53042
rect 9588 52488 9640 52494
rect 9588 52430 9640 52436
rect 9600 50998 9628 52430
rect 9692 52086 9720 53536
rect 9680 52080 9732 52086
rect 9680 52022 9732 52028
rect 9968 51610 9996 54130
rect 10336 53038 10364 56200
rect 10324 53032 10376 53038
rect 10324 52974 10376 52980
rect 10704 52562 10732 56200
rect 11072 53650 11100 56200
rect 11440 54262 11468 56200
rect 11428 54256 11480 54262
rect 11428 54198 11480 54204
rect 11520 54188 11572 54194
rect 11520 54130 11572 54136
rect 11060 53644 11112 53650
rect 11060 53586 11112 53592
rect 10692 52556 10744 52562
rect 10692 52498 10744 52504
rect 10876 52012 10928 52018
rect 10876 51954 10928 51960
rect 9956 51604 10008 51610
rect 9956 51546 10008 51552
rect 9588 50992 9640 50998
rect 9588 50934 9640 50940
rect 10048 49972 10100 49978
rect 10048 49914 10100 49920
rect 9496 49904 9548 49910
rect 9496 49846 9548 49852
rect 10060 47122 10088 49914
rect 10048 47116 10100 47122
rect 10048 47058 10100 47064
rect 9680 45824 9732 45830
rect 9680 45766 9732 45772
rect 9496 45620 9548 45626
rect 9496 45562 9548 45568
rect 9508 44538 9536 45562
rect 9496 44532 9548 44538
rect 9496 44474 9548 44480
rect 9404 43988 9456 43994
rect 9404 43930 9456 43936
rect 9508 43858 9536 44474
rect 9312 43852 9364 43858
rect 9312 43794 9364 43800
rect 9496 43852 9548 43858
rect 9496 43794 9548 43800
rect 9404 43376 9456 43382
rect 9232 43324 9404 43330
rect 9232 43318 9456 43324
rect 9232 43302 9444 43318
rect 9232 42226 9260 43302
rect 9508 43228 9536 43794
rect 9324 43200 9536 43228
rect 9220 42220 9272 42226
rect 9220 42162 9272 42168
rect 9232 41682 9260 42162
rect 9220 41676 9272 41682
rect 9220 41618 9272 41624
rect 9232 40934 9260 41618
rect 9324 41070 9352 43200
rect 9404 42560 9456 42566
rect 9404 42502 9456 42508
rect 9588 42560 9640 42566
rect 9588 42502 9640 42508
rect 9312 41064 9364 41070
rect 9312 41006 9364 41012
rect 9220 40928 9272 40934
rect 9220 40870 9272 40876
rect 9232 40118 9260 40870
rect 9324 40390 9352 41006
rect 9312 40384 9364 40390
rect 9312 40326 9364 40332
rect 9220 40112 9272 40118
rect 9220 40054 9272 40060
rect 9128 39636 9180 39642
rect 9128 39578 9180 39584
rect 9324 38978 9352 40326
rect 9416 39098 9444 42502
rect 9496 42220 9548 42226
rect 9496 42162 9548 42168
rect 9508 41818 9536 42162
rect 9496 41812 9548 41818
rect 9496 41754 9548 41760
rect 9600 39438 9628 42502
rect 9588 39432 9640 39438
rect 9588 39374 9640 39380
rect 9496 39296 9548 39302
rect 9496 39238 9548 39244
rect 9588 39296 9640 39302
rect 9588 39238 9640 39244
rect 9404 39092 9456 39098
rect 9404 39034 9456 39040
rect 9324 38950 9444 38978
rect 9036 38820 9088 38826
rect 9036 38762 9088 38768
rect 8852 38004 8904 38010
rect 8852 37946 8904 37952
rect 8576 37742 8628 37748
rect 8588 37398 8616 37742
rect 8680 37726 8800 37754
rect 8576 37392 8628 37398
rect 8576 37334 8628 37340
rect 8404 37216 8524 37244
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 8300 35760 8352 35766
rect 8300 35702 8352 35708
rect 8312 35290 8340 35702
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 8300 35284 8352 35290
rect 8300 35226 8352 35232
rect 8300 34944 8352 34950
rect 8300 34886 8352 34892
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 7656 34740 7708 34746
rect 7656 34682 7708 34688
rect 7840 33856 7892 33862
rect 7840 33798 7892 33804
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7576 32910 7604 33050
rect 7564 32904 7616 32910
rect 7564 32846 7616 32852
rect 7104 32224 7156 32230
rect 7104 32166 7156 32172
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7668 31754 7696 33594
rect 7748 32360 7800 32366
rect 7748 32302 7800 32308
rect 7576 31726 7696 31754
rect 7012 31272 7064 31278
rect 7012 31214 7064 31220
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 7380 29028 7432 29034
rect 7380 28970 7432 28976
rect 7012 28960 7064 28966
rect 7012 28902 7064 28908
rect 7024 28150 7052 28902
rect 7012 28144 7064 28150
rect 7012 28086 7064 28092
rect 6828 28008 6880 28014
rect 6828 27950 6880 27956
rect 6840 26382 6868 27950
rect 7104 27328 7156 27334
rect 7104 27270 7156 27276
rect 7116 26450 7144 27270
rect 7104 26444 7156 26450
rect 7104 26386 7156 26392
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6840 25974 6868 26318
rect 6828 25968 6880 25974
rect 6828 25910 6880 25916
rect 6840 25362 6868 25910
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 7116 24274 7144 25298
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 7104 24268 7156 24274
rect 7024 24228 7104 24256
rect 7024 22098 7052 24228
rect 7104 24210 7156 24216
rect 6748 22066 6868 22094
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6380 20874 6408 21626
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 6380 20534 6408 20810
rect 6368 20528 6420 20534
rect 6368 20470 6420 20476
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6276 18896 6328 18902
rect 6276 18838 6328 18844
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6564 17746 6592 18158
rect 6656 17882 6684 18770
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6472 16998 6500 17614
rect 6656 17202 6684 17818
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6656 16130 6684 16934
rect 6748 16250 6776 20402
rect 6840 16640 6868 22066
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6932 21690 6960 21830
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19854 6960 20198
rect 7024 20058 7052 21830
rect 7116 21146 7144 22034
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7116 20942 7144 21082
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7116 18630 7144 19110
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 6920 16652 6972 16658
rect 6840 16612 6920 16640
rect 6920 16594 6972 16600
rect 6840 16522 6960 16538
rect 6840 16516 6972 16522
rect 6840 16510 6920 16516
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6840 16130 6868 16510
rect 6920 16458 6972 16464
rect 6656 16102 6868 16130
rect 6840 15162 6868 16102
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6840 14346 6868 15098
rect 7024 15094 7052 15302
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 7116 14958 7144 18566
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6288 7886 6316 14282
rect 6840 14074 6868 14282
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6104 3534 6132 3878
rect 6748 3738 6776 3878
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5368 800 5396 2994
rect 5736 2378 5764 2994
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5736 800 5764 2314
rect 6104 800 6132 3470
rect 6472 2854 6500 3470
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3058 6868 3334
rect 7208 3126 7236 24890
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7300 17882 7328 18634
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7300 14618 7328 15438
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7392 3194 7420 28970
rect 7576 26466 7604 31726
rect 7656 31272 7708 31278
rect 7656 31214 7708 31220
rect 7668 30938 7696 31214
rect 7656 30932 7708 30938
rect 7656 30874 7708 30880
rect 7760 30734 7788 32302
rect 7852 31210 7880 33798
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8312 33674 8340 34886
rect 8404 33844 8432 37216
rect 8680 37194 8708 37726
rect 8668 37188 8720 37194
rect 8668 37130 8720 37136
rect 8576 34740 8628 34746
rect 8576 34682 8628 34688
rect 8588 33998 8616 34682
rect 8576 33992 8628 33998
rect 8576 33934 8628 33940
rect 8404 33816 8616 33844
rect 8312 33646 8524 33674
rect 8392 33516 8444 33522
rect 8392 33458 8444 33464
rect 8404 32978 8432 33458
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 8300 32768 8352 32774
rect 8300 32710 8352 32716
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 8312 32502 8340 32710
rect 8300 32496 8352 32502
rect 8300 32438 8352 32444
rect 8024 32360 8076 32366
rect 8024 32302 8076 32308
rect 8036 31890 8064 32302
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 8300 31272 8352 31278
rect 8300 31214 8352 31220
rect 7840 31204 7892 31210
rect 7840 31146 7892 31152
rect 7748 30728 7800 30734
rect 7748 30670 7800 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 7656 29164 7708 29170
rect 7656 29106 7708 29112
rect 7668 28422 7696 29106
rect 7748 28484 7800 28490
rect 7748 28426 7800 28432
rect 7656 28416 7708 28422
rect 7656 28358 7708 28364
rect 7668 27538 7696 28358
rect 7760 28150 7788 28426
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7748 28144 7800 28150
rect 7748 28086 7800 28092
rect 7760 28014 7788 28086
rect 7748 28008 7800 28014
rect 7748 27950 7800 27956
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7760 27062 7788 27950
rect 7852 27130 7880 28154
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7748 27056 7800 27062
rect 7748 26998 7800 27004
rect 7576 26438 7696 26466
rect 7760 26450 7788 26998
rect 7668 25226 7696 26438
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 7748 25832 7800 25838
rect 7748 25774 7800 25780
rect 7760 25294 7788 25774
rect 7852 25362 7880 27066
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7840 25356 7892 25362
rect 7840 25298 7892 25304
rect 8312 25294 8340 31214
rect 8496 30938 8524 33646
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8404 29306 8432 30534
rect 8588 30258 8616 33816
rect 8680 31754 8708 37130
rect 8864 35714 8892 37946
rect 8944 37664 8996 37670
rect 8944 37606 8996 37612
rect 8956 37262 8984 37606
rect 8944 37256 8996 37262
rect 8944 37198 8996 37204
rect 9048 36854 9076 38762
rect 9220 37324 9272 37330
rect 9220 37266 9272 37272
rect 9312 37324 9364 37330
rect 9312 37266 9364 37272
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9036 36848 9088 36854
rect 9036 36790 9088 36796
rect 8864 35686 8984 35714
rect 8760 35624 8812 35630
rect 8760 35566 8812 35572
rect 8852 35624 8904 35630
rect 8852 35566 8904 35572
rect 8772 34202 8800 35566
rect 8864 34542 8892 35566
rect 8956 35290 8984 35686
rect 8944 35284 8996 35290
rect 8944 35226 8996 35232
rect 8956 35018 8984 35226
rect 8944 35012 8996 35018
rect 8944 34954 8996 34960
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8760 34196 8812 34202
rect 8760 34138 8812 34144
rect 8864 31890 8892 34478
rect 8956 33114 8984 34954
rect 9048 33454 9076 36790
rect 9140 34202 9168 37062
rect 9232 36786 9260 37266
rect 9220 36780 9272 36786
rect 9220 36722 9272 36728
rect 9324 34746 9352 37266
rect 9416 36786 9444 38950
rect 9404 36780 9456 36786
rect 9404 36722 9456 36728
rect 9402 36680 9458 36689
rect 9402 36615 9458 36624
rect 9312 34740 9364 34746
rect 9312 34682 9364 34688
rect 9128 34196 9180 34202
rect 9128 34138 9180 34144
rect 9036 33448 9088 33454
rect 9036 33390 9088 33396
rect 9048 33318 9076 33390
rect 9036 33312 9088 33318
rect 9036 33254 9088 33260
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 9048 32366 9076 33254
rect 9036 32360 9088 32366
rect 9036 32302 9088 32308
rect 8852 31884 8904 31890
rect 8852 31826 8904 31832
rect 8864 31754 8892 31826
rect 8680 31726 8800 31754
rect 8864 31726 8984 31754
rect 8668 30320 8720 30326
rect 8668 30262 8720 30268
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8680 30054 8708 30262
rect 8668 30048 8720 30054
rect 8668 29990 8720 29996
rect 8576 29844 8628 29850
rect 8576 29786 8628 29792
rect 8588 29306 8616 29786
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8576 29300 8628 29306
rect 8576 29242 8628 29248
rect 8576 28552 8628 28558
rect 8576 28494 8628 28500
rect 8588 26994 8616 28494
rect 8576 26988 8628 26994
rect 8576 26930 8628 26936
rect 8588 25974 8616 26930
rect 8576 25968 8628 25974
rect 8576 25910 8628 25916
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 7656 25220 7708 25226
rect 7656 25162 7708 25168
rect 7668 24954 7696 25162
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 8392 24268 8444 24274
rect 8392 24210 8444 24216
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 23526 7512 24006
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7484 23050 7512 23462
rect 7668 23186 7696 24142
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8404 23186 8432 24210
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 8392 23180 8444 23186
rect 8392 23122 8444 23128
rect 7472 23044 7524 23050
rect 7472 22986 7524 22992
rect 7484 21962 7512 22986
rect 7668 22574 7696 23122
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7852 21690 7880 22918
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8404 22710 8432 23122
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8220 21876 8248 22510
rect 8220 21848 8340 21876
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 8312 21622 8340 21848
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 7840 20800 7892 20806
rect 8220 20788 8248 21422
rect 8404 21010 8432 22646
rect 8496 21962 8524 22918
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 8496 21146 8524 21898
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8588 21418 8616 21830
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 8220 20760 8340 20788
rect 7840 20742 7892 20748
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7484 17338 7512 18158
rect 7576 17678 7604 19314
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7668 17626 7696 19654
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7760 17746 7788 19450
rect 7852 19310 7880 20742
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 20482 8340 20760
rect 8220 20454 8340 20482
rect 8404 20466 8432 20946
rect 8496 20874 8524 21082
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8392 20460 8444 20466
rect 8220 19922 8248 20454
rect 8392 20402 8444 20408
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8496 19446 8524 20810
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8588 18426 8616 20878
rect 8680 20806 8708 29990
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7668 17598 7788 17626
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 17338 7696 17478
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7760 17082 7788 17598
rect 7576 17054 7788 17082
rect 7576 16454 7604 17054
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7668 15706 7696 16458
rect 7760 16250 7788 16934
rect 7852 16794 7880 17682
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7852 16114 7880 16730
rect 8312 16658 8340 17614
rect 8496 17542 8524 18226
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 4146 7604 15302
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7668 14618 7696 14894
rect 8312 14822 8340 16594
rect 8404 15706 8432 17070
rect 8496 17066 8524 17478
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8496 16794 8524 17002
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8496 14822 8524 15982
rect 8588 15638 8616 17070
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 8312 14482 8340 14758
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8312 14006 8340 14418
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8220 13530 8248 13806
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8312 12306 8340 13942
rect 8496 13326 8524 14758
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8680 13138 8708 16662
rect 8772 13870 8800 31726
rect 8852 30252 8904 30258
rect 8852 30194 8904 30200
rect 8864 30054 8892 30194
rect 8852 30048 8904 30054
rect 8852 29990 8904 29996
rect 8864 28506 8892 29990
rect 8956 29102 8984 31726
rect 9128 31680 9180 31686
rect 9128 31622 9180 31628
rect 9140 31482 9168 31622
rect 9128 31476 9180 31482
rect 9128 31418 9180 31424
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 8944 29096 8996 29102
rect 8944 29038 8996 29044
rect 8864 28478 8984 28506
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8864 26586 8892 27270
rect 8852 26580 8904 26586
rect 8852 26522 8904 26528
rect 8864 25838 8892 26522
rect 8852 25832 8904 25838
rect 8852 25774 8904 25780
rect 8864 25362 8892 25774
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8864 22778 8892 24006
rect 8852 22772 8904 22778
rect 8852 22714 8904 22720
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8864 20602 8892 22578
rect 8956 20942 8984 28478
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9048 26790 9076 26930
rect 9036 26784 9088 26790
rect 9034 26752 9036 26761
rect 9088 26752 9090 26761
rect 9034 26687 9090 26696
rect 9140 23866 9168 29242
rect 9416 29034 9444 36615
rect 9508 35290 9536 39238
rect 9600 39098 9628 39238
rect 9588 39092 9640 39098
rect 9588 39034 9640 39040
rect 9692 38758 9720 45766
rect 10060 45286 10088 47058
rect 10324 46980 10376 46986
rect 10324 46922 10376 46928
rect 10336 45354 10364 46922
rect 10324 45348 10376 45354
rect 10324 45290 10376 45296
rect 10048 45280 10100 45286
rect 10048 45222 10100 45228
rect 10060 43382 10088 45222
rect 10888 45014 10916 51954
rect 11060 49836 11112 49842
rect 11060 49778 11112 49784
rect 11428 49836 11480 49842
rect 11428 49778 11480 49784
rect 10968 47660 11020 47666
rect 10968 47602 11020 47608
rect 10876 45008 10928 45014
rect 10876 44950 10928 44956
rect 10508 44804 10560 44810
rect 10508 44746 10560 44752
rect 10520 44713 10548 44746
rect 10506 44704 10562 44713
rect 10506 44639 10562 44648
rect 10980 43926 11008 47602
rect 11072 46986 11100 49778
rect 11060 46980 11112 46986
rect 11060 46922 11112 46928
rect 11072 46714 11100 46922
rect 11060 46708 11112 46714
rect 11060 46650 11112 46656
rect 11072 45626 11100 46650
rect 11440 46170 11468 49778
rect 11428 46164 11480 46170
rect 11428 46106 11480 46112
rect 11428 45824 11480 45830
rect 11428 45766 11480 45772
rect 11060 45620 11112 45626
rect 11060 45562 11112 45568
rect 10968 43920 11020 43926
rect 10968 43862 11020 43868
rect 10232 43784 10284 43790
rect 10232 43726 10284 43732
rect 10048 43376 10100 43382
rect 10048 43318 10100 43324
rect 10140 40996 10192 41002
rect 10140 40938 10192 40944
rect 10152 39545 10180 40938
rect 10138 39536 10194 39545
rect 10138 39471 10194 39480
rect 9956 38888 10008 38894
rect 9956 38830 10008 38836
rect 10048 38888 10100 38894
rect 10048 38830 10100 38836
rect 9680 38752 9732 38758
rect 9680 38694 9732 38700
rect 9968 38350 9996 38830
rect 9956 38344 10008 38350
rect 9956 38286 10008 38292
rect 9864 38208 9916 38214
rect 9864 38150 9916 38156
rect 9588 37800 9640 37806
rect 9588 37742 9640 37748
rect 9496 35284 9548 35290
rect 9496 35226 9548 35232
rect 9600 35222 9628 37742
rect 9772 35760 9824 35766
rect 9772 35702 9824 35708
rect 9588 35216 9640 35222
rect 9588 35158 9640 35164
rect 9600 34066 9628 35158
rect 9680 34944 9732 34950
rect 9680 34886 9732 34892
rect 9588 34060 9640 34066
rect 9588 34002 9640 34008
rect 9692 33658 9720 34886
rect 9784 34542 9812 35702
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9784 34202 9812 34478
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9680 33652 9732 33658
rect 9680 33594 9732 33600
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9692 32502 9720 33050
rect 9680 32496 9732 32502
rect 9680 32438 9732 32444
rect 9588 32292 9640 32298
rect 9588 32234 9640 32240
rect 9600 31822 9628 32234
rect 9692 32026 9720 32438
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 9600 30122 9628 31758
rect 9772 30388 9824 30394
rect 9772 30330 9824 30336
rect 9588 30116 9640 30122
rect 9588 30058 9640 30064
rect 9404 29028 9456 29034
rect 9404 28970 9456 28976
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9692 27674 9720 28902
rect 9784 28558 9812 30330
rect 9876 30054 9904 38150
rect 10060 36922 10088 38830
rect 10244 37126 10272 43726
rect 10784 43716 10836 43722
rect 10784 43658 10836 43664
rect 10416 43308 10468 43314
rect 10416 43250 10468 43256
rect 10428 42770 10456 43250
rect 10416 42764 10468 42770
rect 10416 42706 10468 42712
rect 10428 41206 10456 42706
rect 10508 42016 10560 42022
rect 10508 41958 10560 41964
rect 10416 41200 10468 41206
rect 10416 41142 10468 41148
rect 10416 40928 10468 40934
rect 10416 40870 10468 40876
rect 10428 40662 10456 40870
rect 10416 40656 10468 40662
rect 10416 40598 10468 40604
rect 10324 40384 10376 40390
rect 10324 40326 10376 40332
rect 10416 40384 10468 40390
rect 10416 40326 10468 40332
rect 10336 38962 10364 40326
rect 10324 38956 10376 38962
rect 10324 38898 10376 38904
rect 10428 38010 10456 40326
rect 10520 39982 10548 41958
rect 10600 41132 10652 41138
rect 10600 41074 10652 41080
rect 10508 39976 10560 39982
rect 10508 39918 10560 39924
rect 10612 38010 10640 41074
rect 10692 41064 10744 41070
rect 10692 41006 10744 41012
rect 10704 38554 10732 41006
rect 10796 40458 10824 43658
rect 11072 43330 11100 45562
rect 11244 45416 11296 45422
rect 11244 45358 11296 45364
rect 11256 44810 11284 45358
rect 11244 44804 11296 44810
rect 11244 44746 11296 44752
rect 11256 44713 11284 44746
rect 11242 44704 11298 44713
rect 11242 44639 11298 44648
rect 11440 43602 11468 45766
rect 11532 45558 11560 54130
rect 11808 53038 11836 56200
rect 12176 53650 12204 56200
rect 12544 55214 12572 56200
rect 12544 55186 12664 55214
rect 12532 54188 12584 54194
rect 12532 54130 12584 54136
rect 12164 53644 12216 53650
rect 12164 53586 12216 53592
rect 12072 53576 12124 53582
rect 12072 53518 12124 53524
rect 11888 53100 11940 53106
rect 11888 53042 11940 53048
rect 11796 53032 11848 53038
rect 11796 52974 11848 52980
rect 11900 52154 11928 53042
rect 11888 52148 11940 52154
rect 11888 52090 11940 52096
rect 11704 52012 11756 52018
rect 11704 51954 11756 51960
rect 11716 47802 11744 51954
rect 11704 47796 11756 47802
rect 11704 47738 11756 47744
rect 11704 47660 11756 47666
rect 11704 47602 11756 47608
rect 11520 45552 11572 45558
rect 11520 45494 11572 45500
rect 11610 44296 11666 44305
rect 11610 44231 11612 44240
rect 11664 44231 11666 44240
rect 11612 44202 11664 44208
rect 11440 43574 11652 43602
rect 11072 43302 11284 43330
rect 11060 43240 11112 43246
rect 11060 43182 11112 43188
rect 11152 43240 11204 43246
rect 11152 43182 11204 43188
rect 10968 41268 11020 41274
rect 10968 41210 11020 41216
rect 10980 40730 11008 41210
rect 10968 40724 11020 40730
rect 10968 40666 11020 40672
rect 10784 40452 10836 40458
rect 10784 40394 10836 40400
rect 10980 40390 11008 40666
rect 11072 40390 11100 43182
rect 10968 40384 11020 40390
rect 10968 40326 11020 40332
rect 11060 40384 11112 40390
rect 11060 40326 11112 40332
rect 11060 40180 11112 40186
rect 11060 40122 11112 40128
rect 10968 39840 11020 39846
rect 10968 39782 11020 39788
rect 10980 39409 11008 39782
rect 10966 39400 11022 39409
rect 10966 39335 11022 39344
rect 10692 38548 10744 38554
rect 10692 38490 10744 38496
rect 11072 38418 11100 40122
rect 11164 39438 11192 43182
rect 11256 42634 11284 43302
rect 11244 42628 11296 42634
rect 11244 42570 11296 42576
rect 11336 42628 11388 42634
rect 11336 42570 11388 42576
rect 11348 42362 11376 42570
rect 11336 42356 11388 42362
rect 11336 42298 11388 42304
rect 11244 41540 11296 41546
rect 11244 41482 11296 41488
rect 11256 40610 11284 41482
rect 11348 41414 11376 42298
rect 11348 41386 11560 41414
rect 11428 41200 11480 41206
rect 11428 41142 11480 41148
rect 11440 40934 11468 41142
rect 11428 40928 11480 40934
rect 11428 40870 11480 40876
rect 11256 40582 11376 40610
rect 11244 40452 11296 40458
rect 11244 40394 11296 40400
rect 11256 39846 11284 40394
rect 11348 40186 11376 40582
rect 11428 40384 11480 40390
rect 11428 40326 11480 40332
rect 11336 40180 11388 40186
rect 11336 40122 11388 40128
rect 11244 39840 11296 39846
rect 11244 39782 11296 39788
rect 11256 39642 11284 39782
rect 11244 39636 11296 39642
rect 11244 39578 11296 39584
rect 11152 39432 11204 39438
rect 11152 39374 11204 39380
rect 11336 39296 11388 39302
rect 11336 39238 11388 39244
rect 11060 38412 11112 38418
rect 11060 38354 11112 38360
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 10416 38004 10468 38010
rect 10416 37946 10468 37952
rect 10600 38004 10652 38010
rect 10600 37946 10652 37952
rect 10612 37262 10640 37946
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 10232 37120 10284 37126
rect 10232 37062 10284 37068
rect 10612 36922 10640 37198
rect 10876 37120 10928 37126
rect 10876 37062 10928 37068
rect 10048 36916 10100 36922
rect 10048 36858 10100 36864
rect 10600 36916 10652 36922
rect 10600 36858 10652 36864
rect 10060 35154 10088 36858
rect 10324 36712 10376 36718
rect 10324 36654 10376 36660
rect 10336 35834 10364 36654
rect 10324 35828 10376 35834
rect 10324 35770 10376 35776
rect 10336 35154 10364 35770
rect 10692 35692 10744 35698
rect 10692 35634 10744 35640
rect 10048 35148 10100 35154
rect 10048 35090 10100 35096
rect 10324 35148 10376 35154
rect 10324 35090 10376 35096
rect 10336 34678 10364 35090
rect 10704 35018 10732 35634
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10692 35012 10744 35018
rect 10692 34954 10744 34960
rect 10324 34672 10376 34678
rect 10324 34614 10376 34620
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9968 30122 9996 33390
rect 10232 31884 10284 31890
rect 10336 31872 10364 34614
rect 10796 33590 10824 35022
rect 10888 33658 10916 37062
rect 11072 36174 11100 37402
rect 11060 36168 11112 36174
rect 11060 36110 11112 36116
rect 11058 34912 11114 34921
rect 11058 34847 11114 34856
rect 11072 34746 11100 34847
rect 11150 34776 11206 34785
rect 11060 34740 11112 34746
rect 11150 34711 11152 34720
rect 11060 34682 11112 34688
rect 11204 34711 11206 34720
rect 11152 34682 11204 34688
rect 11152 34536 11204 34542
rect 11152 34478 11204 34484
rect 11060 34468 11112 34474
rect 11060 34410 11112 34416
rect 10876 33652 10928 33658
rect 10876 33594 10928 33600
rect 10784 33584 10836 33590
rect 10784 33526 10836 33532
rect 11072 33386 11100 34410
rect 11164 33998 11192 34478
rect 11256 34202 11284 38150
rect 11348 37330 11376 39238
rect 11440 37738 11468 40326
rect 11532 39846 11560 41386
rect 11624 41002 11652 43574
rect 11716 42362 11744 47602
rect 11796 46912 11848 46918
rect 11796 46854 11848 46860
rect 11808 46034 11836 46854
rect 11796 46028 11848 46034
rect 11796 45970 11848 45976
rect 11888 45892 11940 45898
rect 11888 45834 11940 45840
rect 11900 44538 11928 45834
rect 12084 45082 12112 53518
rect 12544 52154 12572 54130
rect 12636 54126 12664 55186
rect 12912 54262 12940 56200
rect 13280 55214 13308 56200
rect 13280 55186 13400 55214
rect 12900 54256 12952 54262
rect 12900 54198 12952 54204
rect 12624 54120 12676 54126
rect 12624 54062 12676 54068
rect 12716 53984 12768 53990
rect 12716 53926 12768 53932
rect 12624 53576 12676 53582
rect 12624 53518 12676 53524
rect 12636 52698 12664 53518
rect 12624 52692 12676 52698
rect 12624 52634 12676 52640
rect 12532 52148 12584 52154
rect 12532 52090 12584 52096
rect 12348 52012 12400 52018
rect 12348 51954 12400 51960
rect 12360 49978 12388 51954
rect 12348 49972 12400 49978
rect 12348 49914 12400 49920
rect 12728 49722 12756 53926
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12808 52488 12860 52494
rect 12808 52430 12860 52436
rect 12636 49694 12756 49722
rect 12440 46368 12492 46374
rect 12440 46310 12492 46316
rect 12532 46368 12584 46374
rect 12532 46310 12584 46316
rect 12452 45554 12480 46310
rect 12544 46034 12572 46310
rect 12532 46028 12584 46034
rect 12532 45970 12584 45976
rect 12452 45526 12572 45554
rect 12256 45484 12308 45490
rect 12256 45426 12308 45432
rect 12164 45348 12216 45354
rect 12164 45290 12216 45296
rect 12176 45098 12204 45290
rect 12268 45286 12296 45426
rect 12256 45280 12308 45286
rect 12254 45248 12256 45257
rect 12308 45248 12310 45257
rect 12254 45183 12310 45192
rect 12072 45076 12124 45082
rect 12176 45070 12296 45098
rect 12072 45018 12124 45024
rect 11888 44532 11940 44538
rect 11888 44474 11940 44480
rect 12268 44266 12296 45070
rect 12544 44878 12572 45526
rect 12532 44872 12584 44878
rect 12532 44814 12584 44820
rect 12348 44328 12400 44334
rect 12348 44270 12400 44276
rect 12256 44260 12308 44266
rect 12256 44202 12308 44208
rect 11704 42356 11756 42362
rect 11704 42298 11756 42304
rect 11796 42220 11848 42226
rect 11796 42162 11848 42168
rect 11704 41608 11756 41614
rect 11704 41550 11756 41556
rect 11612 40996 11664 41002
rect 11612 40938 11664 40944
rect 11716 40050 11744 41550
rect 11704 40044 11756 40050
rect 11704 39986 11756 39992
rect 11520 39840 11572 39846
rect 11520 39782 11572 39788
rect 11532 39506 11560 39782
rect 11520 39500 11572 39506
rect 11520 39442 11572 39448
rect 11704 38888 11756 38894
rect 11704 38830 11756 38836
rect 11716 38350 11744 38830
rect 11808 38554 11836 42162
rect 12072 41540 12124 41546
rect 12072 41482 12124 41488
rect 12084 41274 12112 41482
rect 12072 41268 12124 41274
rect 12072 41210 12124 41216
rect 12268 41070 12296 44202
rect 12360 43994 12388 44270
rect 12636 44010 12664 49694
rect 12820 49434 12848 52430
rect 13372 52426 13400 55186
rect 13648 53174 13676 56200
rect 14016 53582 14044 56200
rect 14004 53576 14056 53582
rect 14004 53518 14056 53524
rect 13636 53168 13688 53174
rect 13636 53110 13688 53116
rect 13648 52698 13676 53110
rect 14384 53106 14412 56200
rect 14752 54330 14780 56200
rect 14740 54324 14792 54330
rect 14740 54266 14792 54272
rect 15120 54176 15148 56200
rect 15200 54188 15252 54194
rect 15120 54148 15200 54176
rect 15200 54130 15252 54136
rect 15016 53984 15068 53990
rect 15016 53926 15068 53932
rect 14648 53440 14700 53446
rect 14648 53382 14700 53388
rect 14372 53100 14424 53106
rect 14372 53042 14424 53048
rect 14004 52964 14056 52970
rect 14004 52906 14056 52912
rect 13636 52692 13688 52698
rect 13636 52634 13688 52640
rect 14016 52601 14044 52906
rect 14002 52592 14058 52601
rect 14002 52527 14058 52536
rect 13360 52420 13412 52426
rect 13360 52362 13412 52368
rect 13372 52154 13400 52362
rect 13360 52148 13412 52154
rect 13360 52090 13412 52096
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12808 49428 12860 49434
rect 12808 49370 12860 49376
rect 13544 49224 13596 49230
rect 13544 49166 13596 49172
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 12808 46912 12860 46918
rect 12808 46854 12860 46860
rect 12716 46028 12768 46034
rect 12716 45970 12768 45976
rect 12728 44334 12756 45970
rect 12820 45830 12848 46854
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 12808 45824 12860 45830
rect 12808 45766 12860 45772
rect 13452 45824 13504 45830
rect 13452 45766 13504 45772
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 12808 44736 12860 44742
rect 12808 44678 12860 44684
rect 12716 44328 12768 44334
rect 12716 44270 12768 44276
rect 12348 43988 12400 43994
rect 12348 43930 12400 43936
rect 12544 43982 12664 44010
rect 12348 43648 12400 43654
rect 12348 43590 12400 43596
rect 12256 41064 12308 41070
rect 12256 41006 12308 41012
rect 11980 40928 12032 40934
rect 11980 40870 12032 40876
rect 11992 40526 12020 40870
rect 12072 40588 12124 40594
rect 12072 40530 12124 40536
rect 11980 40520 12032 40526
rect 11980 40462 12032 40468
rect 11980 40112 12032 40118
rect 11980 40054 12032 40060
rect 11992 39506 12020 40054
rect 11980 39500 12032 39506
rect 11900 39460 11980 39488
rect 11796 38548 11848 38554
rect 11796 38490 11848 38496
rect 11704 38344 11756 38350
rect 11704 38286 11756 38292
rect 11428 37732 11480 37738
rect 11428 37674 11480 37680
rect 11612 37664 11664 37670
rect 11612 37606 11664 37612
rect 11336 37324 11388 37330
rect 11336 37266 11388 37272
rect 11428 34740 11480 34746
rect 11428 34682 11480 34688
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 11244 33992 11296 33998
rect 11244 33934 11296 33940
rect 11060 33380 11112 33386
rect 11060 33322 11112 33328
rect 10968 32836 11020 32842
rect 10968 32778 11020 32784
rect 10600 32496 10652 32502
rect 10600 32438 10652 32444
rect 10284 31844 10364 31872
rect 10232 31826 10284 31832
rect 10612 31754 10640 32438
rect 10980 32230 11008 32778
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10980 31754 11008 32166
rect 11072 32008 11100 33322
rect 11152 32020 11204 32026
rect 11072 31980 11152 32008
rect 11152 31962 11204 31968
rect 11256 31754 11284 33934
rect 11440 33862 11468 34682
rect 11520 34672 11572 34678
rect 11520 34614 11572 34620
rect 11532 34202 11560 34614
rect 11520 34196 11572 34202
rect 11520 34138 11572 34144
rect 11532 34066 11560 34138
rect 11520 34060 11572 34066
rect 11520 34002 11572 34008
rect 11428 33856 11480 33862
rect 11428 33798 11480 33804
rect 11440 33522 11468 33798
rect 11428 33516 11480 33522
rect 11428 33458 11480 33464
rect 11428 31884 11480 31890
rect 11428 31826 11480 31832
rect 10612 31748 10744 31754
rect 10612 31726 10692 31748
rect 10692 31690 10744 31696
rect 10796 31726 11008 31754
rect 11164 31726 11284 31754
rect 10704 30666 10732 31690
rect 10692 30660 10744 30666
rect 10692 30602 10744 30608
rect 9956 30116 10008 30122
rect 9956 30058 10008 30064
rect 9864 30048 9916 30054
rect 9864 29990 9916 29996
rect 10324 29504 10376 29510
rect 10324 29446 10376 29452
rect 10336 29170 10364 29446
rect 10324 29164 10376 29170
rect 10324 29106 10376 29112
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9784 28014 9812 28494
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 9312 27464 9364 27470
rect 9312 27406 9364 27412
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9232 25974 9260 26250
rect 9220 25968 9272 25974
rect 9220 25910 9272 25916
rect 9232 24750 9260 25910
rect 9324 24818 9352 27406
rect 9496 27396 9548 27402
rect 9496 27338 9548 27344
rect 9508 25362 9536 27338
rect 9784 26858 9812 27950
rect 10796 26908 10824 31726
rect 11164 30802 11192 31726
rect 11336 31340 11388 31346
rect 11336 31282 11388 31288
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 10876 30660 10928 30666
rect 10876 30602 10928 30608
rect 10888 29510 10916 30602
rect 11164 30274 11192 30738
rect 11072 30258 11192 30274
rect 11060 30252 11192 30258
rect 11112 30246 11192 30252
rect 11060 30194 11112 30200
rect 11256 29714 11284 31078
rect 11348 30598 11376 31282
rect 11440 30802 11468 31826
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 11440 30682 11468 30738
rect 11440 30654 11560 30682
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 11348 30190 11376 30534
rect 11336 30184 11388 30190
rect 11336 30126 11388 30132
rect 11532 29714 11560 30654
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11072 28694 11100 29106
rect 11428 29028 11480 29034
rect 11428 28970 11480 28976
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10612 26880 10824 26908
rect 9772 26852 9824 26858
rect 9772 26794 9824 26800
rect 10048 26308 10100 26314
rect 10048 26250 10100 26256
rect 9680 25764 9732 25770
rect 9680 25706 9732 25712
rect 9496 25356 9548 25362
rect 9496 25298 9548 25304
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 9508 24954 9536 25094
rect 9496 24948 9548 24954
rect 9496 24890 9548 24896
rect 9692 24886 9720 25706
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9324 24206 9352 24754
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9968 23866 9996 24006
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 9680 23248 9732 23254
rect 9680 23190 9732 23196
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8956 20466 8984 20742
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8864 15978 8892 18634
rect 8956 18578 8984 20402
rect 9048 20058 9076 21490
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9140 18970 9168 20334
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 8956 18550 9168 18578
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8956 15858 8984 17478
rect 8864 15830 8984 15858
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8404 13110 8708 13138
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7760 8634 7788 8774
rect 7852 8634 7880 11698
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8312 7954 8340 12242
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8404 6914 8432 13110
rect 8864 13002 8892 15830
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 14074 8984 14214
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8680 12974 8892 13002
rect 8680 12434 8708 12974
rect 8956 12866 8984 13806
rect 8588 12406 8708 12434
rect 8772 12838 8984 12866
rect 8588 7818 8616 12406
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8312 6886 8432 6914
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 8312 4690 8340 6886
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3602 7512 4014
rect 8772 3942 8800 12838
rect 9048 12434 9076 18362
rect 8956 12406 9076 12434
rect 9140 12434 9168 18550
rect 9232 16658 9260 21966
rect 9600 21894 9628 22918
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9324 20942 9352 21082
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9600 20806 9628 21558
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9324 17066 9352 20334
rect 9692 20330 9720 23190
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 21010 9812 23054
rect 9772 21004 9824 21010
rect 9824 20964 9904 20992
rect 9772 20946 9824 20952
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9416 18086 9444 19246
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9508 18290 9536 18634
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9416 17134 9444 18022
rect 9600 17338 9628 19654
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9784 18426 9812 18702
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9876 18222 9904 20964
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9876 17338 9904 18158
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 10060 17202 10088 26250
rect 10232 25288 10284 25294
rect 10232 25230 10284 25236
rect 10244 25158 10272 25230
rect 10232 25152 10284 25158
rect 10230 25120 10232 25129
rect 10284 25120 10286 25129
rect 10230 25055 10286 25064
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10336 23254 10364 24210
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10140 21480 10192 21486
rect 10140 21422 10192 21428
rect 10152 21350 10180 21422
rect 10140 21344 10192 21350
rect 10138 21312 10140 21321
rect 10192 21312 10194 21321
rect 10138 21247 10194 21256
rect 10140 21004 10192 21010
rect 10140 20946 10192 20952
rect 10152 19514 10180 20946
rect 10244 19922 10272 23122
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10520 22778 10548 22918
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10336 20602 10364 21626
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10428 21010 10456 21286
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10612 20346 10640 26880
rect 10888 25362 10916 28358
rect 11072 26450 11100 28630
rect 11152 27396 11204 27402
rect 11152 27338 11204 27344
rect 11164 26926 11192 27338
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11164 26790 11192 26862
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 11164 26194 11192 26386
rect 11256 26382 11284 26862
rect 11440 26518 11468 28970
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11428 26512 11480 26518
rect 11428 26454 11480 26460
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 11164 26166 11284 26194
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10336 20318 10640 20346
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10244 18766 10272 19858
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10336 18630 10364 20318
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10520 19854 10548 20198
rect 10508 19848 10560 19854
rect 10506 19816 10508 19825
rect 10560 19816 10562 19825
rect 10506 19751 10562 19760
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9416 15502 9444 17070
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9508 16590 9536 16662
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 14822 9444 15438
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9416 13802 9444 14758
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9140 12406 9260 12434
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8956 3738 8984 12406
rect 9232 11778 9260 12406
rect 9692 12306 9720 14758
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9876 11898 9904 16390
rect 10060 16114 10088 17138
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10060 15994 10088 16050
rect 9968 15966 10088 15994
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9140 11750 9260 11778
rect 9140 4758 9168 11750
rect 9968 10810 9996 15966
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 14346 10088 15846
rect 10152 14346 10180 18566
rect 10336 17814 10364 18566
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10046 10976 10102 10985
rect 10046 10911 10102 10920
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9218 7984 9274 7993
rect 9218 7919 9274 7928
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9232 3738 9260 7919
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6472 800 6500 2790
rect 6840 800 6868 2994
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1970 7144 2246
rect 7104 1964 7156 1970
rect 7104 1906 7156 1912
rect 7208 800 7236 2382
rect 7576 800 7604 2382
rect 7852 1986 7880 3334
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8312 3058 8340 3538
rect 9416 3534 9444 3878
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8390 3224 8446 3233
rect 8390 3159 8392 3168
rect 8444 3159 8446 3168
rect 8392 3130 8444 3136
rect 8680 3058 8708 3334
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 7852 1958 7972 1986
rect 7944 800 7972 1958
rect 8312 800 8340 2994
rect 8680 800 8708 2994
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8956 2106 8984 2382
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9048 800 9076 2994
rect 9416 800 9444 3470
rect 9508 2990 9536 4966
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9600 3126 9628 3946
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3534 9812 3878
rect 10060 3738 10088 10911
rect 10428 4078 10456 19314
rect 10520 18970 10548 19654
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10520 18222 10548 18770
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10520 17542 10548 18158
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10520 13734 10548 17070
rect 10612 15502 10640 20198
rect 10704 19378 10732 23802
rect 11164 23798 11192 24550
rect 11152 23792 11204 23798
rect 11152 23734 11204 23740
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10796 21962 10824 22442
rect 10784 21956 10836 21962
rect 10784 21898 10836 21904
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10980 20890 11008 21422
rect 10796 20862 11008 20890
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10704 16250 10732 18838
rect 10796 17377 10824 20862
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20398 11008 20742
rect 11072 20602 11100 22918
rect 11256 22094 11284 26166
rect 11440 25498 11468 26454
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 11440 25158 11468 25434
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11348 23186 11376 23666
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11164 22066 11284 22094
rect 11164 21622 11192 22066
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10968 20392 11020 20398
rect 11020 20340 11100 20346
rect 10968 20334 11100 20340
rect 10888 19514 10916 20334
rect 10980 20318 11100 20334
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 11072 18834 11100 20318
rect 11256 19990 11284 20878
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 11256 19310 11284 19926
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11164 18426 11192 18634
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 10782 17368 10838 17377
rect 10782 17303 10838 17312
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10796 15094 10824 17303
rect 10888 16658 10916 18362
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10980 17338 11008 18226
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 11164 17610 11192 18158
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10980 17134 11008 17274
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15638 10916 15982
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10796 14006 10824 15030
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10520 6914 10548 13670
rect 10796 12782 10824 13942
rect 11072 13530 11100 15302
rect 11164 14958 11192 17546
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11164 14482 11192 14894
rect 11256 14618 11284 15302
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11256 14074 11284 14554
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11256 12986 11284 14010
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 11256 12306 11284 12922
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10612 11694 10640 12038
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10520 6886 10640 6914
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9784 800 9812 3470
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10152 800 10180 2382
rect 10520 800 10548 2994
rect 10612 2514 10640 6886
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10888 800 10916 3470
rect 10980 3058 11008 3878
rect 11072 3194 11100 11698
rect 11256 11082 11284 12038
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11256 3058 11284 3334
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11164 1902 11192 2382
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 11256 800 11284 2994
rect 11348 2854 11376 22374
rect 11440 22098 11468 24142
rect 11532 22778 11560 28494
rect 11624 26314 11652 37606
rect 11704 36168 11756 36174
rect 11704 36110 11756 36116
rect 11716 35834 11744 36110
rect 11796 36032 11848 36038
rect 11796 35974 11848 35980
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11808 35018 11836 35974
rect 11796 35012 11848 35018
rect 11796 34954 11848 34960
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11716 34066 11744 34886
rect 11900 34134 11928 39460
rect 11980 39442 12032 39448
rect 11980 38480 12032 38486
rect 11980 38422 12032 38428
rect 11992 37466 12020 38422
rect 11980 37460 12032 37466
rect 11980 37402 12032 37408
rect 11980 37120 12032 37126
rect 11980 37062 12032 37068
rect 11992 34678 12020 37062
rect 12084 36174 12112 40530
rect 12360 39642 12388 43590
rect 12544 40526 12572 43982
rect 12624 43852 12676 43858
rect 12624 43794 12676 43800
rect 12636 42770 12664 43794
rect 12728 43246 12756 44270
rect 12820 43450 12848 44678
rect 13464 44334 13492 45766
rect 13556 45354 13584 49166
rect 14188 46912 14240 46918
rect 14188 46854 14240 46860
rect 14096 46708 14148 46714
rect 14096 46650 14148 46656
rect 13820 46504 13872 46510
rect 13820 46446 13872 46452
rect 13832 45626 13860 46446
rect 13820 45620 13872 45626
rect 13820 45562 13872 45568
rect 13728 45484 13780 45490
rect 13728 45426 13780 45432
rect 13544 45348 13596 45354
rect 13544 45290 13596 45296
rect 13636 45348 13688 45354
rect 13636 45290 13688 45296
rect 13648 44878 13676 45290
rect 13636 44872 13688 44878
rect 13636 44814 13688 44820
rect 13452 44328 13504 44334
rect 13452 44270 13504 44276
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12808 43444 12860 43450
rect 12808 43386 12860 43392
rect 12716 43240 12768 43246
rect 12716 43182 12768 43188
rect 12624 42764 12676 42770
rect 12624 42706 12676 42712
rect 12624 42628 12676 42634
rect 12624 42570 12676 42576
rect 12636 41818 12664 42570
rect 12624 41812 12676 41818
rect 12624 41754 12676 41760
rect 12532 40520 12584 40526
rect 12532 40462 12584 40468
rect 12636 40066 12664 41754
rect 12728 41614 12756 43182
rect 13464 43110 13492 44270
rect 12808 43104 12860 43110
rect 12808 43046 12860 43052
rect 13452 43104 13504 43110
rect 13452 43046 13504 43052
rect 12716 41608 12768 41614
rect 12716 41550 12768 41556
rect 12716 40384 12768 40390
rect 12716 40326 12768 40332
rect 12452 40038 12664 40066
rect 12348 39636 12400 39642
rect 12348 39578 12400 39584
rect 12452 39574 12480 40038
rect 12728 39574 12756 40326
rect 12440 39568 12492 39574
rect 12440 39510 12492 39516
rect 12716 39568 12768 39574
rect 12716 39510 12768 39516
rect 12440 39092 12492 39098
rect 12440 39034 12492 39040
rect 12452 39001 12480 39034
rect 12438 38992 12494 39001
rect 12820 38944 12848 43046
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 13464 42838 13492 43046
rect 13452 42832 13504 42838
rect 13452 42774 13504 42780
rect 13360 42560 13412 42566
rect 13360 42502 13412 42508
rect 13372 42362 13400 42502
rect 13740 42362 13768 45426
rect 13820 45416 13872 45422
rect 13820 45358 13872 45364
rect 13832 43994 13860 45358
rect 13820 43988 13872 43994
rect 13820 43930 13872 43936
rect 13360 42356 13412 42362
rect 13360 42298 13412 42304
rect 13728 42356 13780 42362
rect 13728 42298 13780 42304
rect 13728 42220 13780 42226
rect 13728 42162 13780 42168
rect 13360 42152 13412 42158
rect 13360 42094 13412 42100
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12898 39536 12954 39545
rect 12898 39471 12954 39480
rect 12992 39500 13044 39506
rect 12438 38927 12494 38936
rect 12544 38916 12848 38944
rect 12346 38856 12402 38865
rect 12346 38791 12348 38800
rect 12400 38791 12402 38800
rect 12348 38762 12400 38768
rect 12254 38448 12310 38457
rect 12254 38383 12310 38392
rect 12440 38412 12492 38418
rect 12268 36582 12296 38383
rect 12440 38354 12492 38360
rect 12164 36576 12216 36582
rect 12164 36518 12216 36524
rect 12256 36576 12308 36582
rect 12256 36518 12308 36524
rect 12348 36576 12400 36582
rect 12348 36518 12400 36524
rect 12176 36174 12204 36518
rect 12072 36168 12124 36174
rect 12072 36110 12124 36116
rect 12164 36168 12216 36174
rect 12164 36110 12216 36116
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 12084 34746 12112 35634
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 11980 34672 12032 34678
rect 11980 34614 12032 34620
rect 12176 34524 12204 36110
rect 12268 36038 12296 36518
rect 12256 36032 12308 36038
rect 12256 35974 12308 35980
rect 12360 34626 12388 36518
rect 12452 35494 12480 38354
rect 12544 36242 12572 38916
rect 12912 38876 12940 39471
rect 12992 39442 13044 39448
rect 13004 39409 13032 39442
rect 12990 39400 13046 39409
rect 12990 39335 13046 39344
rect 13268 39296 13320 39302
rect 13268 39238 13320 39244
rect 12820 38848 12940 38876
rect 12624 38820 12676 38826
rect 12624 38762 12676 38768
rect 12636 37262 12664 38762
rect 12820 38282 12848 38848
rect 13280 38758 13308 39238
rect 13268 38752 13320 38758
rect 13268 38694 13320 38700
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12808 38276 12860 38282
rect 12808 38218 12860 38224
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12636 36854 12664 37198
rect 12624 36848 12676 36854
rect 12624 36790 12676 36796
rect 12716 36644 12768 36650
rect 12716 36586 12768 36592
rect 12532 36236 12584 36242
rect 12532 36178 12584 36184
rect 12728 36122 12756 36586
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 13372 36378 13400 42094
rect 13740 41274 13768 42162
rect 13912 42016 13964 42022
rect 13912 41958 13964 41964
rect 13728 41268 13780 41274
rect 13728 41210 13780 41216
rect 13820 41268 13872 41274
rect 13820 41210 13872 41216
rect 13450 41168 13506 41177
rect 13450 41103 13452 41112
rect 13504 41103 13506 41112
rect 13636 41132 13688 41138
rect 13452 41074 13504 41080
rect 13832 41120 13860 41210
rect 13688 41092 13860 41120
rect 13636 41074 13688 41080
rect 13464 40934 13492 41074
rect 13544 40996 13596 41002
rect 13544 40938 13596 40944
rect 13452 40928 13504 40934
rect 13452 40870 13504 40876
rect 13556 40730 13584 40938
rect 13544 40724 13596 40730
rect 13544 40666 13596 40672
rect 13452 40520 13504 40526
rect 13452 40462 13504 40468
rect 13464 40186 13492 40462
rect 13544 40384 13596 40390
rect 13544 40326 13596 40332
rect 13452 40180 13504 40186
rect 13452 40122 13504 40128
rect 13452 39840 13504 39846
rect 13452 39782 13504 39788
rect 13464 39001 13492 39782
rect 13450 38992 13506 39001
rect 13450 38927 13506 38936
rect 13452 38752 13504 38758
rect 13452 38694 13504 38700
rect 13360 36372 13412 36378
rect 13360 36314 13412 36320
rect 12544 36094 12756 36122
rect 12544 35630 12572 36094
rect 12716 36032 12768 36038
rect 12716 35974 12768 35980
rect 12900 36032 12952 36038
rect 12900 35974 12952 35980
rect 12728 35737 12756 35974
rect 12714 35728 12770 35737
rect 12714 35663 12770 35672
rect 12532 35624 12584 35630
rect 12532 35566 12584 35572
rect 12440 35488 12492 35494
rect 12440 35430 12492 35436
rect 12084 34496 12204 34524
rect 12268 34598 12388 34626
rect 11888 34128 11940 34134
rect 11888 34070 11940 34076
rect 11704 34060 11756 34066
rect 11704 34002 11756 34008
rect 11796 33516 11848 33522
rect 11796 33458 11848 33464
rect 11704 32360 11756 32366
rect 11704 32302 11756 32308
rect 11716 32026 11744 32302
rect 11704 32020 11756 32026
rect 11704 31962 11756 31968
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11716 27062 11744 31826
rect 11808 31754 11836 33458
rect 12084 31890 12112 34496
rect 12164 33924 12216 33930
rect 12164 33866 12216 33872
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 11808 31726 12020 31754
rect 11888 30592 11940 30598
rect 11888 30534 11940 30540
rect 11900 30326 11928 30534
rect 11888 30320 11940 30326
rect 11888 30262 11940 30268
rect 11888 30116 11940 30122
rect 11888 30058 11940 30064
rect 11796 30048 11848 30054
rect 11796 29990 11848 29996
rect 11704 27056 11756 27062
rect 11704 26998 11756 27004
rect 11716 26450 11744 26998
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11716 24138 11744 24550
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11532 22681 11560 22714
rect 11518 22672 11574 22681
rect 11518 22607 11574 22616
rect 11428 22092 11480 22098
rect 11808 22094 11836 29990
rect 11900 29850 11928 30058
rect 11888 29844 11940 29850
rect 11888 29786 11940 29792
rect 11992 29730 12020 31726
rect 12072 31136 12124 31142
rect 12072 31078 12124 31084
rect 11900 29702 12020 29730
rect 11900 26994 11928 29702
rect 12084 27538 12112 31078
rect 12176 30938 12204 33866
rect 12268 33658 12296 34598
rect 12348 34536 12400 34542
rect 12348 34478 12400 34484
rect 12256 33652 12308 33658
rect 12256 33594 12308 33600
rect 12360 33454 12388 34478
rect 12452 34134 12480 35430
rect 12544 34542 12572 35566
rect 12912 35476 12940 35974
rect 13464 35766 13492 38694
rect 13452 35760 13504 35766
rect 13452 35702 13504 35708
rect 13452 35624 13504 35630
rect 13452 35566 13504 35572
rect 12820 35448 12940 35476
rect 13360 35488 13412 35494
rect 12624 35284 12676 35290
rect 12624 35226 12676 35232
rect 12532 34536 12584 34542
rect 12532 34478 12584 34484
rect 12440 34128 12492 34134
rect 12440 34070 12492 34076
rect 12348 33448 12400 33454
rect 12348 33390 12400 33396
rect 12636 32026 12664 35226
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12728 34746 12756 34886
rect 12716 34740 12768 34746
rect 12716 34682 12768 34688
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 12360 31346 12388 31826
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12164 30932 12216 30938
rect 12164 30874 12216 30880
rect 12440 30592 12492 30598
rect 12440 30534 12492 30540
rect 12346 30424 12402 30433
rect 12452 30410 12480 30534
rect 12402 30382 12480 30410
rect 12346 30359 12402 30368
rect 12360 30054 12388 30359
rect 12728 30326 12756 33798
rect 12820 32842 12848 35448
rect 13360 35430 13412 35436
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 13372 35290 13400 35430
rect 13360 35284 13412 35290
rect 13360 35226 13412 35232
rect 13464 35154 13492 35566
rect 13452 35148 13504 35154
rect 13452 35090 13504 35096
rect 13452 35012 13504 35018
rect 13452 34954 13504 34960
rect 13464 34542 13492 34954
rect 13452 34536 13504 34542
rect 13452 34478 13504 34484
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 13360 33856 13412 33862
rect 13360 33798 13412 33804
rect 13372 33425 13400 33798
rect 13358 33416 13414 33425
rect 13358 33351 13360 33360
rect 13412 33351 13414 33360
rect 13360 33322 13412 33328
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12808 32836 12860 32842
rect 12808 32778 12860 32784
rect 12820 32570 12848 32778
rect 12808 32564 12860 32570
rect 12808 32506 12860 32512
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12820 31890 12848 32370
rect 13464 32366 13492 34478
rect 13556 33930 13584 40326
rect 13648 40118 13676 41074
rect 13728 40724 13780 40730
rect 13728 40666 13780 40672
rect 13636 40112 13688 40118
rect 13636 40054 13688 40060
rect 13740 37670 13768 40666
rect 13924 39030 13952 41958
rect 14002 40760 14058 40769
rect 14002 40695 14004 40704
rect 14056 40695 14058 40704
rect 14004 40666 14056 40672
rect 14016 40594 14044 40666
rect 14004 40588 14056 40594
rect 14004 40530 14056 40536
rect 14108 39574 14136 46650
rect 14200 46646 14228 46854
rect 14188 46640 14240 46646
rect 14188 46582 14240 46588
rect 14200 46170 14228 46582
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14200 45898 14228 46106
rect 14188 45892 14240 45898
rect 14188 45834 14240 45840
rect 14556 45892 14608 45898
rect 14556 45834 14608 45840
rect 14280 44804 14332 44810
rect 14280 44746 14332 44752
rect 14188 42696 14240 42702
rect 14188 42638 14240 42644
rect 14200 41614 14228 42638
rect 14188 41608 14240 41614
rect 14188 41550 14240 41556
rect 14096 39568 14148 39574
rect 14096 39510 14148 39516
rect 13820 39024 13872 39030
rect 13820 38966 13872 38972
rect 13912 39024 13964 39030
rect 13912 38966 13964 38972
rect 13832 38758 13860 38966
rect 14200 38962 14228 41550
rect 14188 38956 14240 38962
rect 14188 38898 14240 38904
rect 14188 38820 14240 38826
rect 14108 38780 14188 38808
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13832 38400 13860 38694
rect 13832 38372 13952 38400
rect 13820 38276 13872 38282
rect 13820 38218 13872 38224
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 13636 37188 13688 37194
rect 13636 37130 13688 37136
rect 13648 34746 13676 37130
rect 13832 37126 13860 38218
rect 13820 37120 13872 37126
rect 13820 37062 13872 37068
rect 13728 36848 13780 36854
rect 13728 36790 13780 36796
rect 13740 36718 13768 36790
rect 13728 36712 13780 36718
rect 13728 36654 13780 36660
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 13636 34604 13688 34610
rect 13636 34546 13688 34552
rect 13544 33924 13596 33930
rect 13544 33866 13596 33872
rect 13452 32360 13504 32366
rect 13358 32328 13414 32337
rect 13452 32302 13504 32308
rect 13358 32263 13414 32272
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 12808 31884 12860 31890
rect 12808 31826 12860 31832
rect 13372 31822 13400 32263
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13648 31754 13676 34546
rect 13740 32434 13768 36654
rect 13924 35834 13952 38372
rect 14004 37800 14056 37806
rect 14004 37742 14056 37748
rect 14016 37262 14044 37742
rect 14004 37256 14056 37262
rect 14004 37198 14056 37204
rect 13912 35828 13964 35834
rect 13912 35770 13964 35776
rect 14108 33862 14136 38780
rect 14188 38762 14240 38768
rect 14292 37806 14320 44746
rect 14372 44532 14424 44538
rect 14372 44474 14424 44480
rect 14384 42362 14412 44474
rect 14568 44402 14596 45834
rect 14556 44396 14608 44402
rect 14556 44338 14608 44344
rect 14372 42356 14424 42362
rect 14372 42298 14424 42304
rect 14372 41812 14424 41818
rect 14372 41754 14424 41760
rect 14280 37800 14332 37806
rect 14280 37742 14332 37748
rect 14384 37398 14412 41754
rect 14464 40656 14516 40662
rect 14464 40598 14516 40604
rect 14476 37466 14504 40598
rect 14568 40458 14596 44338
rect 14556 40452 14608 40458
rect 14556 40394 14608 40400
rect 14556 38752 14608 38758
rect 14556 38694 14608 38700
rect 14568 37942 14596 38694
rect 14556 37936 14608 37942
rect 14556 37878 14608 37884
rect 14464 37460 14516 37466
rect 14464 37402 14516 37408
rect 14372 37392 14424 37398
rect 14372 37334 14424 37340
rect 14372 36576 14424 36582
rect 14372 36518 14424 36524
rect 14280 36100 14332 36106
rect 14280 36042 14332 36048
rect 14292 34202 14320 36042
rect 14188 34196 14240 34202
rect 14188 34138 14240 34144
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 14200 34105 14228 34138
rect 14186 34096 14242 34105
rect 14186 34031 14242 34040
rect 14096 33856 14148 33862
rect 14096 33798 14148 33804
rect 14108 33318 14136 33798
rect 14280 33516 14332 33522
rect 14280 33458 14332 33464
rect 14096 33312 14148 33318
rect 14094 33280 14096 33289
rect 14148 33280 14150 33289
rect 14094 33215 14150 33224
rect 14188 32768 14240 32774
rect 14188 32710 14240 32716
rect 14200 32502 14228 32710
rect 14188 32496 14240 32502
rect 14188 32438 14240 32444
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 13648 31748 13780 31754
rect 13648 31726 13728 31748
rect 13728 31690 13780 31696
rect 14004 31680 14056 31686
rect 14004 31622 14056 31628
rect 13912 31408 13964 31414
rect 13912 31350 13964 31356
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 13924 30802 13952 31350
rect 13912 30796 13964 30802
rect 13912 30738 13964 30744
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12360 29345 12388 29990
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 12346 29336 12402 29345
rect 12346 29271 12402 29280
rect 12348 29164 12400 29170
rect 12348 29106 12400 29112
rect 12360 28626 12388 29106
rect 12624 29028 12676 29034
rect 12624 28970 12676 28976
rect 12348 28620 12400 28626
rect 12348 28562 12400 28568
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12360 27674 12388 28018
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12348 27668 12400 27674
rect 12348 27610 12400 27616
rect 12256 27600 12308 27606
rect 12256 27542 12308 27548
rect 12072 27532 12124 27538
rect 12072 27474 12124 27480
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11992 27130 12020 27270
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11900 23662 11928 25842
rect 12072 25424 12124 25430
rect 12072 25366 12124 25372
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11992 24614 12020 24754
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 12084 23866 12112 25366
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12268 23730 12296 27542
rect 12360 25906 12388 27610
rect 12452 26926 12480 27950
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 12360 24138 12388 24550
rect 12452 24274 12480 26862
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12544 25294 12572 25774
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 11888 23656 11940 23662
rect 11888 23598 11940 23604
rect 12530 23216 12586 23225
rect 12530 23151 12586 23160
rect 12544 23050 12572 23151
rect 12532 23044 12584 23050
rect 12532 22986 12584 22992
rect 12544 22778 12572 22986
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12544 22166 12572 22374
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 11428 22034 11480 22040
rect 11716 22066 11836 22094
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11440 18970 11468 21354
rect 11624 21350 11652 21490
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11624 21146 11652 21286
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11716 20806 11744 22066
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 11808 21690 11836 21898
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11808 21350 11836 21626
rect 12452 21622 12480 21830
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11716 20602 11744 20742
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11716 20058 11744 20538
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11440 11762 11468 17274
rect 11624 17270 11652 19110
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 16454 11560 16526
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11532 15026 11560 16390
rect 11716 16114 11744 18022
rect 11808 17678 11836 21286
rect 12452 21010 12480 21286
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12636 20942 12664 28970
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12808 28620 12860 28626
rect 12808 28562 12860 28568
rect 12820 28218 12848 28562
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13464 28218 13492 28358
rect 12808 28212 12860 28218
rect 12808 28154 12860 28160
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 13360 28144 13412 28150
rect 13360 28086 13412 28092
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12728 22438 12756 27270
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 12992 26512 13044 26518
rect 13372 26466 13400 28086
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 12992 26454 13044 26460
rect 13004 26042 13032 26454
rect 13280 26438 13400 26466
rect 13280 26042 13308 26438
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 13280 25702 13308 25978
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 12820 25362 12848 25638
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13372 25498 13400 26182
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 22710 13400 23462
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12820 22098 12848 22510
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12808 22092 12860 22098
rect 13464 22094 13492 27270
rect 13556 25974 13584 28358
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 13648 27062 13676 27474
rect 13740 27130 13768 30534
rect 13924 29850 13952 30738
rect 13912 29844 13964 29850
rect 13912 29786 13964 29792
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13544 25968 13596 25974
rect 13544 25910 13596 25916
rect 13636 25696 13688 25702
rect 13636 25638 13688 25644
rect 13464 22066 13584 22094
rect 12808 22034 12860 22040
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 11992 19446 12020 20470
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 16040 11664 16046
rect 11664 15988 11744 15994
rect 11612 15982 11744 15988
rect 11624 15966 11744 15982
rect 11716 15570 11744 15966
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 15366 11744 15506
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11532 8430 11560 14962
rect 11716 13802 11744 15302
rect 11808 14074 11836 16118
rect 11900 15162 11928 18566
rect 12084 18426 12112 18634
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 17066 12020 18022
rect 12084 17882 12112 18226
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 12268 17814 12296 19654
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12360 18834 12388 19246
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11900 8430 11928 14214
rect 11992 11898 12020 17002
rect 12360 16114 12388 18770
rect 12544 18698 12572 20742
rect 12728 19854 12756 21830
rect 12820 21010 12848 22034
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13268 21616 13320 21622
rect 13268 21558 13320 21564
rect 13280 21418 13308 21558
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 13372 21350 13400 21830
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 13556 19786 13584 22066
rect 13648 21962 13676 25638
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13740 24834 13768 25094
rect 13740 24806 13952 24834
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23730 13860 24006
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13740 23118 13768 23598
rect 13832 23186 13860 23666
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13924 22778 13952 24806
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 13728 22160 13780 22166
rect 13728 22102 13780 22108
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 12728 19446 12756 19654
rect 13464 19446 13492 19654
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12452 17377 12480 17682
rect 12438 17368 12494 17377
rect 12438 17303 12494 17312
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12452 15450 12480 15506
rect 12360 15422 12480 15450
rect 12360 14958 12388 15422
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12162 13016 12218 13025
rect 12162 12951 12164 12960
rect 12216 12951 12218 12960
rect 12164 12922 12216 12928
rect 12360 12434 12388 14894
rect 12176 12406 12388 12434
rect 12176 12306 12204 12406
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12176 11694 12204 12242
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11218 12204 11630
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12268 11082 12296 12174
rect 12452 11778 12480 15030
rect 12544 12434 12572 18634
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17134 12664 17478
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 14618 12664 16594
rect 12728 15094 12756 19382
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12820 16454 12848 17274
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13372 16658 13400 18634
rect 13464 17082 13492 19382
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13648 18222 13676 18838
rect 13740 18442 13768 22102
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13832 21350 13860 21830
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 13924 21418 13952 21558
rect 13912 21412 13964 21418
rect 13912 21354 13964 21360
rect 14016 21350 14044 31622
rect 14096 31136 14148 31142
rect 14096 31078 14148 31084
rect 14108 29102 14136 31078
rect 14200 29238 14228 32438
rect 14292 30938 14320 33458
rect 14384 32502 14412 36518
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 14372 32496 14424 32502
rect 14372 32438 14424 32444
rect 14476 31142 14504 33458
rect 14660 32586 14688 53382
rect 14924 45824 14976 45830
rect 14924 45766 14976 45772
rect 14740 45484 14792 45490
rect 14740 45426 14792 45432
rect 14752 44198 14780 45426
rect 14936 44402 14964 45766
rect 14924 44396 14976 44402
rect 14924 44338 14976 44344
rect 14740 44192 14792 44198
rect 14740 44134 14792 44140
rect 14752 43858 14780 44134
rect 14740 43852 14792 43858
rect 14740 43794 14792 43800
rect 14752 42294 14780 43794
rect 14924 43648 14976 43654
rect 14924 43590 14976 43596
rect 14832 43308 14884 43314
rect 14832 43250 14884 43256
rect 14844 42566 14872 43250
rect 14936 42906 14964 43590
rect 14924 42900 14976 42906
rect 14924 42842 14976 42848
rect 14832 42560 14884 42566
rect 14832 42502 14884 42508
rect 14844 42378 14872 42502
rect 14844 42350 14964 42378
rect 14740 42288 14792 42294
rect 14740 42230 14792 42236
rect 14740 42084 14792 42090
rect 14740 42026 14792 42032
rect 14752 40730 14780 42026
rect 14844 41274 14872 42350
rect 14936 42294 14964 42350
rect 14924 42288 14976 42294
rect 14924 42230 14976 42236
rect 14832 41268 14884 41274
rect 14832 41210 14884 41216
rect 14740 40724 14792 40730
rect 14740 40666 14792 40672
rect 14844 40594 14872 41210
rect 14832 40588 14884 40594
rect 14832 40530 14884 40536
rect 14924 40452 14976 40458
rect 14924 40394 14976 40400
rect 14832 39976 14884 39982
rect 14832 39918 14884 39924
rect 14844 39846 14872 39918
rect 14936 39846 14964 40394
rect 14832 39840 14884 39846
rect 14832 39782 14884 39788
rect 14924 39840 14976 39846
rect 14924 39782 14976 39788
rect 14924 38344 14976 38350
rect 14924 38286 14976 38292
rect 14740 38208 14792 38214
rect 14740 38150 14792 38156
rect 14752 38010 14780 38150
rect 14740 38004 14792 38010
rect 14740 37946 14792 37952
rect 14832 37324 14884 37330
rect 14832 37266 14884 37272
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 14752 34746 14780 37062
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 14844 32774 14872 37266
rect 14936 36242 14964 38286
rect 14924 36236 14976 36242
rect 14924 36178 14976 36184
rect 14832 32768 14884 32774
rect 14832 32710 14884 32716
rect 14660 32558 14780 32586
rect 14648 32496 14700 32502
rect 14648 32438 14700 32444
rect 14660 31686 14688 32438
rect 14648 31680 14700 31686
rect 14648 31622 14700 31628
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14280 30932 14332 30938
rect 14280 30874 14332 30880
rect 14660 30802 14688 31078
rect 14648 30796 14700 30802
rect 14648 30738 14700 30744
rect 14752 30326 14780 32558
rect 14832 32224 14884 32230
rect 14832 32166 14884 32172
rect 14924 32224 14976 32230
rect 14924 32166 14976 32172
rect 14740 30320 14792 30326
rect 14740 30262 14792 30268
rect 14372 30048 14424 30054
rect 14372 29990 14424 29996
rect 14188 29232 14240 29238
rect 14188 29174 14240 29180
rect 14096 29096 14148 29102
rect 14096 29038 14148 29044
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 14108 27674 14136 28562
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14096 27668 14148 27674
rect 14096 27610 14148 27616
rect 14108 26466 14136 27610
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14200 27334 14228 27406
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14200 26586 14228 27270
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 14292 26518 14320 27814
rect 14280 26512 14332 26518
rect 14108 26438 14228 26466
rect 14280 26454 14332 26460
rect 14096 25220 14148 25226
rect 14096 25162 14148 25168
rect 13820 21344 13872 21350
rect 14004 21344 14056 21350
rect 13820 21286 13872 21292
rect 14002 21312 14004 21321
rect 14056 21312 14058 21321
rect 13832 20806 13860 21286
rect 14002 21247 14058 21256
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 14108 20534 14136 25162
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14200 19904 14228 26438
rect 14384 25430 14412 29990
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14752 28422 14780 28562
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 14476 27334 14504 28086
rect 14844 27334 14872 32166
rect 14936 31278 14964 32166
rect 14924 31272 14976 31278
rect 14924 31214 14976 31220
rect 15028 30682 15056 53926
rect 15488 53582 15516 56200
rect 15856 55214 15884 56200
rect 15856 55186 15976 55214
rect 15752 53984 15804 53990
rect 15752 53926 15804 53932
rect 15476 53576 15528 53582
rect 15476 53518 15528 53524
rect 15568 52964 15620 52970
rect 15568 52906 15620 52912
rect 15476 47116 15528 47122
rect 15476 47058 15528 47064
rect 15292 46640 15344 46646
rect 15344 46600 15424 46628
rect 15292 46582 15344 46588
rect 15396 45898 15424 46600
rect 15384 45892 15436 45898
rect 15384 45834 15436 45840
rect 15488 45778 15516 47058
rect 15396 45750 15516 45778
rect 15396 45286 15424 45750
rect 15580 45554 15608 52906
rect 15488 45526 15608 45554
rect 15384 45280 15436 45286
rect 15384 45222 15436 45228
rect 15200 44192 15252 44198
rect 15200 44134 15252 44140
rect 15108 43104 15160 43110
rect 15108 43046 15160 43052
rect 15120 36854 15148 43046
rect 15212 41682 15240 44134
rect 15488 43450 15516 45526
rect 15568 45280 15620 45286
rect 15568 45222 15620 45228
rect 15580 44810 15608 45222
rect 15568 44804 15620 44810
rect 15568 44746 15620 44752
rect 15580 43994 15608 44746
rect 15568 43988 15620 43994
rect 15568 43930 15620 43936
rect 15476 43444 15528 43450
rect 15476 43386 15528 43392
rect 15580 43330 15608 43930
rect 15396 43302 15608 43330
rect 15292 43172 15344 43178
rect 15292 43114 15344 43120
rect 15200 41676 15252 41682
rect 15200 41618 15252 41624
rect 15304 41138 15332 43114
rect 15292 41132 15344 41138
rect 15292 41074 15344 41080
rect 15292 40928 15344 40934
rect 15292 40870 15344 40876
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 15108 36848 15160 36854
rect 15108 36790 15160 36796
rect 15212 36038 15240 37810
rect 15304 37126 15332 40870
rect 15396 40050 15424 43302
rect 15476 43240 15528 43246
rect 15476 43182 15528 43188
rect 15568 43240 15620 43246
rect 15568 43182 15620 43188
rect 15488 42106 15516 43182
rect 15580 42226 15608 43182
rect 15660 42628 15712 42634
rect 15660 42570 15712 42576
rect 15568 42220 15620 42226
rect 15568 42162 15620 42168
rect 15488 42078 15608 42106
rect 15476 42016 15528 42022
rect 15476 41958 15528 41964
rect 15488 41070 15516 41958
rect 15580 41414 15608 42078
rect 15672 41614 15700 42570
rect 15660 41608 15712 41614
rect 15660 41550 15712 41556
rect 15580 41386 15700 41414
rect 15476 41064 15528 41070
rect 15476 41006 15528 41012
rect 15568 41064 15620 41070
rect 15568 41006 15620 41012
rect 15384 40044 15436 40050
rect 15384 39986 15436 39992
rect 15580 39642 15608 41006
rect 15568 39636 15620 39642
rect 15568 39578 15620 39584
rect 15580 39438 15608 39578
rect 15568 39432 15620 39438
rect 15568 39374 15620 39380
rect 15476 39296 15528 39302
rect 15476 39238 15528 39244
rect 15568 39296 15620 39302
rect 15568 39238 15620 39244
rect 15382 38856 15438 38865
rect 15382 38791 15384 38800
rect 15436 38791 15438 38800
rect 15384 38762 15436 38768
rect 15382 38448 15438 38457
rect 15382 38383 15384 38392
rect 15436 38383 15438 38392
rect 15384 38354 15436 38360
rect 15384 38208 15436 38214
rect 15384 38150 15436 38156
rect 15396 38010 15424 38150
rect 15384 38004 15436 38010
rect 15384 37946 15436 37952
rect 15384 37800 15436 37806
rect 15384 37742 15436 37748
rect 15292 37120 15344 37126
rect 15292 37062 15344 37068
rect 15292 36916 15344 36922
rect 15292 36858 15344 36864
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 15120 33658 15148 33866
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 15120 32298 15148 32710
rect 15108 32292 15160 32298
rect 15108 32234 15160 32240
rect 15120 31686 15148 32234
rect 15108 31680 15160 31686
rect 15108 31622 15160 31628
rect 15212 30734 15240 33390
rect 15200 30728 15252 30734
rect 15028 30654 15148 30682
rect 15200 30670 15252 30676
rect 15120 30598 15148 30654
rect 15108 30592 15160 30598
rect 15108 30534 15160 30540
rect 15016 27872 15068 27878
rect 15016 27814 15068 27820
rect 14924 27532 14976 27538
rect 14924 27474 14976 27480
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14476 26994 14504 27270
rect 14936 27062 14964 27474
rect 14924 27056 14976 27062
rect 14924 26998 14976 27004
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14476 26790 14504 26930
rect 15028 26926 15056 27814
rect 15120 27402 15148 30534
rect 15304 29850 15332 36858
rect 15396 36174 15424 37742
rect 15488 36378 15516 39238
rect 15580 37942 15608 39238
rect 15672 38962 15700 41386
rect 15660 38956 15712 38962
rect 15660 38898 15712 38904
rect 15672 38865 15700 38898
rect 15658 38856 15714 38865
rect 15658 38791 15714 38800
rect 15660 38412 15712 38418
rect 15660 38354 15712 38360
rect 15568 37936 15620 37942
rect 15568 37878 15620 37884
rect 15672 37874 15700 38354
rect 15660 37868 15712 37874
rect 15660 37810 15712 37816
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 15384 36168 15436 36174
rect 15384 36110 15436 36116
rect 15384 36032 15436 36038
rect 15384 35974 15436 35980
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15108 27396 15160 27402
rect 15108 27338 15160 27344
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 14464 26784 14516 26790
rect 14464 26726 14516 26732
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 14372 25424 14424 25430
rect 14372 25366 14424 25372
rect 14476 22710 14504 26726
rect 14556 26512 14608 26518
rect 14556 26454 14608 26460
rect 14568 23186 14596 26454
rect 14752 26382 14780 26726
rect 15028 26518 15056 26726
rect 15016 26512 15068 26518
rect 14922 26480 14978 26489
rect 14832 26444 14884 26450
rect 15016 26454 15068 26460
rect 14922 26415 14978 26424
rect 14832 26386 14884 26392
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14648 26240 14700 26246
rect 14648 26182 14700 26188
rect 14660 25294 14688 26182
rect 14752 25362 14780 26318
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14844 24818 14872 26386
rect 14936 26314 14964 26415
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 13924 19876 14228 19904
rect 13740 18426 13860 18442
rect 13740 18420 13872 18426
rect 13740 18414 13820 18420
rect 13636 18216 13688 18222
rect 13556 18176 13636 18204
rect 13556 17270 13584 18176
rect 13636 18158 13688 18164
rect 13634 17640 13690 17649
rect 13634 17575 13636 17584
rect 13688 17575 13690 17584
rect 13636 17546 13688 17552
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13464 17054 13584 17082
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12820 14074 12848 15914
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13464 15570 13492 16526
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13556 15450 13584 17054
rect 13372 15422 13584 15450
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14226 13400 15422
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13464 14482 13492 15030
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 14362 13492 14418
rect 13464 14334 13584 14362
rect 13372 14198 13492 14226
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12898 13424 12954 13433
rect 12716 13388 12768 13394
rect 12898 13359 12900 13368
rect 12716 13330 12768 13336
rect 12952 13359 12954 13368
rect 12900 13330 12952 13336
rect 12544 12406 12664 12434
rect 12452 11750 12572 11778
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12452 11354 12480 11630
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12544 11286 12572 11750
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11992 4146 12020 10542
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11624 800 11652 4014
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11992 800 12020 2450
rect 12084 2446 12112 10406
rect 12636 9654 12664 12406
rect 12728 11218 12756 13330
rect 13372 12986 13400 13874
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13464 12866 13492 14198
rect 13372 12838 13492 12866
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 2038 12296 2246
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 12360 800 12388 1838
rect 12728 800 12756 3402
rect 12820 2446 12848 12650
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13004 11082 13032 11290
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 13004 10810 13032 11018
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13372 5030 13400 12838
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 9738 13492 12582
rect 13556 11665 13584 14334
rect 13542 11656 13598 11665
rect 13542 11591 13598 11600
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 10538 13584 11494
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13464 9710 13584 9738
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13464 4690 13492 9522
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13556 4146 13584 9710
rect 13648 6914 13676 17546
rect 13740 17134 13768 18414
rect 13820 18362 13872 18368
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13832 17338 13860 18226
rect 13924 18086 13952 19876
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 14016 17338 14044 18566
rect 14200 18222 14228 19246
rect 14292 18358 14320 21286
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13740 14550 13768 17070
rect 13832 16658 13860 17070
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12646 13768 13330
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11558 13768 12174
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13726 11384 13782 11393
rect 13726 11319 13782 11328
rect 13740 9586 13768 11319
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13648 6886 13768 6914
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 13096 870 13216 898
rect 13096 800 13124 870
rect 3252 734 3464 762
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13188 762 13216 870
rect 13372 762 13400 2926
rect 13464 800 13492 4014
rect 13648 2582 13676 4626
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13740 1970 13768 6886
rect 13832 2802 13860 16594
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14108 15162 14136 15914
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14016 14346 14044 14962
rect 14200 14958 14228 18158
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14384 13938 14412 21966
rect 14476 21554 14504 22374
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14476 20874 14504 21490
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14476 19378 14504 20538
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13924 11354 13952 11630
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14016 6914 14044 13262
rect 13924 6886 14044 6914
rect 13924 2922 13952 6886
rect 14200 3534 14228 13806
rect 14292 11898 14320 13874
rect 14384 13530 14412 13874
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14384 12850 14412 13330
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14292 3058 14320 11018
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13832 2774 13952 2802
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13728 1964 13780 1970
rect 13728 1906 13780 1912
rect 13832 800 13860 2314
rect 13924 2106 13952 2774
rect 13912 2100 13964 2106
rect 13912 2042 13964 2048
rect 14200 800 14228 2926
rect 14476 2650 14504 17682
rect 14568 17134 14596 20402
rect 14660 20058 14688 22034
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14752 21321 14780 21422
rect 14738 21312 14794 21321
rect 14738 21247 14794 21256
rect 14844 20754 14872 24550
rect 14936 24410 14964 26250
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14752 20726 14872 20754
rect 14752 20602 14780 20726
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14660 18834 14688 19994
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14752 18766 14780 20198
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14738 18456 14794 18465
rect 14648 18420 14700 18426
rect 14738 18391 14740 18400
rect 14648 18362 14700 18368
rect 14792 18391 14794 18400
rect 14740 18362 14792 18368
rect 14660 17814 14688 18362
rect 14648 17808 14700 17814
rect 14648 17750 14700 17756
rect 14752 17746 14780 18362
rect 14936 17898 14964 24346
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 15028 22166 15056 22646
rect 15120 22438 15148 26794
rect 15198 26616 15254 26625
rect 15198 26551 15254 26560
rect 15212 26246 15240 26551
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 15212 22710 15240 23258
rect 15200 22704 15252 22710
rect 15200 22646 15252 22652
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 15016 22160 15068 22166
rect 15016 22102 15068 22108
rect 15028 20482 15056 22102
rect 15212 22094 15240 22170
rect 15304 22094 15332 29786
rect 15396 29238 15424 35974
rect 15672 35290 15700 37810
rect 15660 35284 15712 35290
rect 15660 35226 15712 35232
rect 15660 35148 15712 35154
rect 15660 35090 15712 35096
rect 15568 33992 15620 33998
rect 15672 33980 15700 35090
rect 15620 33952 15700 33980
rect 15568 33934 15620 33940
rect 15568 33312 15620 33318
rect 15568 33254 15620 33260
rect 15476 31272 15528 31278
rect 15476 31214 15528 31220
rect 15488 30394 15516 31214
rect 15476 30388 15528 30394
rect 15476 30330 15528 30336
rect 15580 29306 15608 33254
rect 15672 32978 15700 33952
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15660 32836 15712 32842
rect 15660 32778 15712 32784
rect 15672 32570 15700 32778
rect 15660 32564 15712 32570
rect 15660 32506 15712 32512
rect 15672 32026 15700 32506
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 15660 31748 15712 31754
rect 15660 31690 15712 31696
rect 15672 31482 15700 31690
rect 15660 31476 15712 31482
rect 15660 31418 15712 31424
rect 15568 29300 15620 29306
rect 15568 29242 15620 29248
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15660 29232 15712 29238
rect 15660 29174 15712 29180
rect 15568 29164 15620 29170
rect 15568 29106 15620 29112
rect 15384 29028 15436 29034
rect 15384 28970 15436 28976
rect 15396 25226 15424 28970
rect 15580 28422 15608 29106
rect 15672 29034 15700 29174
rect 15660 29028 15712 29034
rect 15660 28970 15712 28976
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15672 28370 15700 28970
rect 15764 28490 15792 53926
rect 15844 53440 15896 53446
rect 15844 53382 15896 53388
rect 15856 45554 15884 53382
rect 15948 53106 15976 55186
rect 16224 54330 16252 56200
rect 16212 54324 16264 54330
rect 16212 54266 16264 54272
rect 16592 53786 16620 56200
rect 16960 54194 16988 56200
rect 16948 54188 17000 54194
rect 16948 54130 17000 54136
rect 16764 54052 16816 54058
rect 16764 53994 16816 54000
rect 16580 53780 16632 53786
rect 16580 53722 16632 53728
rect 16592 53582 16620 53722
rect 16580 53576 16632 53582
rect 16580 53518 16632 53524
rect 15936 53100 15988 53106
rect 15936 53042 15988 53048
rect 16120 52896 16172 52902
rect 16120 52838 16172 52844
rect 16132 47802 16160 52838
rect 16304 52488 16356 52494
rect 16304 52430 16356 52436
rect 16120 47796 16172 47802
rect 16120 47738 16172 47744
rect 16120 46640 16172 46646
rect 16120 46582 16172 46588
rect 16132 45830 16160 46582
rect 16212 46164 16264 46170
rect 16212 46106 16264 46112
rect 16224 46034 16252 46106
rect 16212 46028 16264 46034
rect 16212 45970 16264 45976
rect 16120 45824 16172 45830
rect 16120 45766 16172 45772
rect 15856 45526 15976 45554
rect 15844 43648 15896 43654
rect 15844 43590 15896 43596
rect 15856 42566 15884 43590
rect 15844 42560 15896 42566
rect 15844 42502 15896 42508
rect 15844 42016 15896 42022
rect 15844 41958 15896 41964
rect 15856 41274 15884 41958
rect 15948 41414 15976 45526
rect 16224 44742 16252 45970
rect 16212 44736 16264 44742
rect 16212 44678 16264 44684
rect 16120 43920 16172 43926
rect 16120 43862 16172 43868
rect 16132 42242 16160 43862
rect 16212 42288 16264 42294
rect 16132 42236 16212 42242
rect 16132 42230 16264 42236
rect 16132 42214 16252 42230
rect 15948 41386 16068 41414
rect 15844 41268 15896 41274
rect 15844 41210 15896 41216
rect 15856 39545 15884 41210
rect 15936 41132 15988 41138
rect 15936 41074 15988 41080
rect 15948 40186 15976 41074
rect 15936 40180 15988 40186
rect 15936 40122 15988 40128
rect 15936 39976 15988 39982
rect 15936 39918 15988 39924
rect 15842 39536 15898 39545
rect 15842 39471 15898 39480
rect 15844 38888 15896 38894
rect 15844 38830 15896 38836
rect 15856 38418 15884 38830
rect 15844 38412 15896 38418
rect 15844 38354 15896 38360
rect 15948 38298 15976 39918
rect 15856 38270 15976 38298
rect 15856 36802 15884 38270
rect 15936 37324 15988 37330
rect 15936 37266 15988 37272
rect 15948 37126 15976 37266
rect 15936 37120 15988 37126
rect 15936 37062 15988 37068
rect 15948 36922 15976 37062
rect 15936 36916 15988 36922
rect 15936 36858 15988 36864
rect 15856 36786 15976 36802
rect 15856 36780 15988 36786
rect 15856 36774 15936 36780
rect 15936 36722 15988 36728
rect 15948 36582 15976 36722
rect 15936 36576 15988 36582
rect 15936 36518 15988 36524
rect 15948 33318 15976 36518
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15948 31142 15976 31622
rect 16040 31414 16068 41386
rect 16132 38486 16160 42214
rect 16316 41414 16344 52430
rect 16580 47116 16632 47122
rect 16500 47076 16580 47104
rect 16500 46170 16528 47076
rect 16580 47058 16632 47064
rect 16672 46504 16724 46510
rect 16672 46446 16724 46452
rect 16684 46170 16712 46446
rect 16488 46164 16540 46170
rect 16488 46106 16540 46112
rect 16672 46164 16724 46170
rect 16672 46106 16724 46112
rect 16580 45824 16632 45830
rect 16580 45766 16632 45772
rect 16592 45082 16620 45766
rect 16776 45554 16804 53994
rect 17040 53984 17092 53990
rect 17038 53952 17040 53961
rect 17092 53952 17094 53961
rect 17038 53887 17094 53896
rect 17328 53582 17356 56200
rect 17696 55214 17724 56200
rect 18064 56114 18092 56200
rect 18156 56114 18184 56222
rect 18064 56086 18184 56114
rect 17696 55186 17908 55214
rect 17880 54312 17908 55186
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17880 54284 18000 54312
rect 17972 54194 18000 54284
rect 17960 54188 18012 54194
rect 17960 54130 18012 54136
rect 18340 53582 18368 56222
rect 18418 56200 18474 57000
rect 18786 56200 18842 57000
rect 19154 56200 19210 57000
rect 19522 56200 19578 57000
rect 19890 56200 19946 57000
rect 20258 56200 20314 57000
rect 20626 56200 20682 57000
rect 20994 56200 21050 57000
rect 21362 56200 21418 57000
rect 21730 56200 21786 57000
rect 22098 56200 22154 57000
rect 22466 56200 22522 57000
rect 22834 56200 22890 57000
rect 23202 56200 23258 57000
rect 23570 56200 23626 57000
rect 24490 56264 24546 56273
rect 18432 55214 18460 56200
rect 18432 55186 18644 55214
rect 18616 54194 18644 55186
rect 18512 54188 18564 54194
rect 18512 54130 18564 54136
rect 18604 54188 18656 54194
rect 18604 54130 18656 54136
rect 18420 53984 18472 53990
rect 18420 53926 18472 53932
rect 17316 53576 17368 53582
rect 17316 53518 17368 53524
rect 18328 53576 18380 53582
rect 18328 53518 18380 53524
rect 17040 53440 17092 53446
rect 17040 53382 17092 53388
rect 16948 47456 17000 47462
rect 16948 47398 17000 47404
rect 16856 46912 16908 46918
rect 16856 46854 16908 46860
rect 16868 46646 16896 46854
rect 16856 46640 16908 46646
rect 16856 46582 16908 46588
rect 16856 45892 16908 45898
rect 16856 45834 16908 45840
rect 16868 45558 16896 45834
rect 16684 45526 16804 45554
rect 16856 45552 16908 45558
rect 16580 45076 16632 45082
rect 16580 45018 16632 45024
rect 16684 44962 16712 45526
rect 16856 45494 16908 45500
rect 16592 44934 16712 44962
rect 16488 44736 16540 44742
rect 16488 44678 16540 44684
rect 16500 44334 16528 44678
rect 16488 44328 16540 44334
rect 16488 44270 16540 44276
rect 16396 41472 16448 41478
rect 16396 41414 16448 41420
rect 16224 41386 16344 41414
rect 16120 38480 16172 38486
rect 16120 38422 16172 38428
rect 16132 37874 16160 38422
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 16120 37732 16172 37738
rect 16120 37674 16172 37680
rect 16132 37466 16160 37674
rect 16120 37460 16172 37466
rect 16120 37402 16172 37408
rect 16120 33448 16172 33454
rect 16120 33390 16172 33396
rect 16132 32434 16160 33390
rect 16224 33114 16252 41386
rect 16304 40928 16356 40934
rect 16304 40870 16356 40876
rect 16316 40594 16344 40870
rect 16304 40588 16356 40594
rect 16304 40530 16356 40536
rect 16304 39296 16356 39302
rect 16304 39238 16356 39244
rect 16316 38758 16344 39238
rect 16304 38752 16356 38758
rect 16304 38694 16356 38700
rect 16408 38418 16436 41414
rect 16500 41206 16528 44270
rect 16592 43450 16620 44934
rect 16672 44396 16724 44402
rect 16672 44338 16724 44344
rect 16580 43444 16632 43450
rect 16580 43386 16632 43392
rect 16580 42220 16632 42226
rect 16580 42162 16632 42168
rect 16592 41682 16620 42162
rect 16684 41818 16712 44338
rect 16856 43716 16908 43722
rect 16856 43658 16908 43664
rect 16764 42696 16816 42702
rect 16764 42638 16816 42644
rect 16672 41812 16724 41818
rect 16672 41754 16724 41760
rect 16580 41676 16632 41682
rect 16580 41618 16632 41624
rect 16488 41200 16540 41206
rect 16488 41142 16540 41148
rect 16488 39500 16540 39506
rect 16488 39442 16540 39448
rect 16396 38412 16448 38418
rect 16396 38354 16448 38360
rect 16500 38010 16528 39442
rect 16592 38486 16620 41618
rect 16776 40662 16804 42638
rect 16764 40656 16816 40662
rect 16764 40598 16816 40604
rect 16868 40186 16896 43658
rect 16960 41682 16988 47398
rect 17052 46050 17080 53382
rect 17328 53242 17356 53518
rect 17592 53440 17644 53446
rect 17592 53382 17644 53388
rect 18328 53440 18380 53446
rect 18328 53382 18380 53388
rect 17316 53236 17368 53242
rect 17316 53178 17368 53184
rect 17316 48204 17368 48210
rect 17316 48146 17368 48152
rect 17132 46980 17184 46986
rect 17132 46922 17184 46928
rect 17144 46170 17172 46922
rect 17328 46374 17356 48146
rect 17604 48142 17632 53382
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 18340 48278 18368 53382
rect 18328 48272 18380 48278
rect 18328 48214 18380 48220
rect 17592 48136 17644 48142
rect 17592 48078 17644 48084
rect 17684 48000 17736 48006
rect 17684 47942 17736 47948
rect 17408 47592 17460 47598
rect 17408 47534 17460 47540
rect 17420 46714 17448 47534
rect 17500 47184 17552 47190
rect 17500 47126 17552 47132
rect 17408 46708 17460 46714
rect 17408 46650 17460 46656
rect 17316 46368 17368 46374
rect 17316 46310 17368 46316
rect 17132 46164 17184 46170
rect 17132 46106 17184 46112
rect 17052 46022 17264 46050
rect 17040 45960 17092 45966
rect 17040 45902 17092 45908
rect 17052 44742 17080 45902
rect 17040 44736 17092 44742
rect 17040 44678 17092 44684
rect 16948 41676 17000 41682
rect 16948 41618 17000 41624
rect 17052 41070 17080 44678
rect 17132 44328 17184 44334
rect 17132 44270 17184 44276
rect 17144 43246 17172 44270
rect 17236 43738 17264 46022
rect 17420 45490 17448 46650
rect 17408 45484 17460 45490
rect 17408 45426 17460 45432
rect 17236 43710 17448 43738
rect 17224 43648 17276 43654
rect 17224 43590 17276 43596
rect 17132 43240 17184 43246
rect 17132 43182 17184 43188
rect 17040 41064 17092 41070
rect 17040 41006 17092 41012
rect 16856 40180 16908 40186
rect 16856 40122 16908 40128
rect 16764 40112 16816 40118
rect 16764 40054 16816 40060
rect 16672 39568 16724 39574
rect 16672 39510 16724 39516
rect 16684 39137 16712 39510
rect 16670 39128 16726 39137
rect 16670 39063 16726 39072
rect 16672 38752 16724 38758
rect 16672 38694 16724 38700
rect 16580 38480 16632 38486
rect 16580 38422 16632 38428
rect 16488 38004 16540 38010
rect 16488 37946 16540 37952
rect 16580 37120 16632 37126
rect 16394 37088 16450 37097
rect 16580 37062 16632 37068
rect 16394 37023 16450 37032
rect 16408 36922 16436 37023
rect 16396 36916 16448 36922
rect 16396 36858 16448 36864
rect 16592 36378 16620 37062
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 16304 35488 16356 35494
rect 16304 35430 16356 35436
rect 16212 33108 16264 33114
rect 16212 33050 16264 33056
rect 16120 32428 16172 32434
rect 16120 32370 16172 32376
rect 16028 31408 16080 31414
rect 16026 31376 16028 31385
rect 16080 31376 16082 31385
rect 16026 31311 16082 31320
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 15844 30864 15896 30870
rect 15844 30806 15896 30812
rect 15856 29306 15884 30806
rect 16028 30796 16080 30802
rect 16028 30738 16080 30744
rect 15844 29300 15896 29306
rect 15844 29242 15896 29248
rect 15936 29096 15988 29102
rect 15936 29038 15988 29044
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15476 27396 15528 27402
rect 15476 27338 15528 27344
rect 15488 26586 15516 27338
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15384 25220 15436 25226
rect 15384 25162 15436 25168
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15212 22066 15332 22094
rect 15212 21690 15240 22066
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15304 21554 15332 21898
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15028 20454 15148 20482
rect 15016 20392 15068 20398
rect 15014 20360 15016 20369
rect 15068 20360 15070 20369
rect 15014 20295 15070 20304
rect 15120 19922 15148 20454
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15120 19786 15148 19858
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15120 19446 15148 19722
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 15212 18970 15240 19450
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14844 17870 14964 17898
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14568 15706 14596 17070
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15366 14596 15438
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14568 12434 14596 15302
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 13954 14688 14350
rect 14752 14074 14780 15302
rect 14844 15042 14872 17870
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14936 17542 14964 17750
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 15120 15434 15148 16118
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15028 15337 15056 15370
rect 15014 15328 15070 15337
rect 15014 15263 15070 15272
rect 15028 15094 15056 15263
rect 15016 15088 15068 15094
rect 14844 15014 14964 15042
rect 15016 15030 15068 15036
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14660 13926 14780 13954
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13326 14688 13738
rect 14752 13734 14780 13926
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12918 14688 13262
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14568 12406 14688 12434
rect 14660 3602 14688 12406
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14844 3126 14872 14826
rect 14936 13394 14964 15014
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 15212 12986 15240 17478
rect 15304 14090 15332 21082
rect 15488 17678 15516 25094
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15580 14822 15608 28358
rect 15672 28342 15792 28370
rect 15660 28212 15712 28218
rect 15660 28154 15712 28160
rect 15672 28121 15700 28154
rect 15658 28112 15714 28121
rect 15658 28047 15714 28056
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 15672 26450 15700 26998
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15764 24698 15792 28342
rect 15948 28082 15976 29038
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 16040 26926 16068 30738
rect 16120 27532 16172 27538
rect 16120 27474 16172 27480
rect 16028 26920 16080 26926
rect 16028 26862 16080 26868
rect 15936 26036 15988 26042
rect 16040 26024 16068 26862
rect 15988 25996 16068 26024
rect 15936 25978 15988 25984
rect 16132 25974 16160 27474
rect 16120 25968 16172 25974
rect 16120 25910 16172 25916
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 16040 25498 16068 25774
rect 16028 25492 16080 25498
rect 16028 25434 16080 25440
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15856 24818 15884 25094
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15764 24670 15884 24698
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15764 23662 15792 24346
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15856 22982 15884 24670
rect 16040 24070 16068 25230
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 16040 23662 16068 24006
rect 16132 23866 16160 24754
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 16224 23236 16252 33050
rect 16316 31482 16344 35430
rect 16684 34048 16712 38694
rect 16776 38214 16804 40054
rect 16948 39840 17000 39846
rect 16948 39782 17000 39788
rect 16764 38208 16816 38214
rect 16764 38150 16816 38156
rect 16776 34116 16804 38150
rect 16856 38004 16908 38010
rect 16856 37946 16908 37952
rect 16868 36174 16896 37946
rect 16960 37874 16988 39782
rect 17144 39506 17172 43182
rect 17236 41274 17264 43590
rect 17316 42764 17368 42770
rect 17316 42706 17368 42712
rect 17328 41614 17356 42706
rect 17316 41608 17368 41614
rect 17316 41550 17368 41556
rect 17224 41268 17276 41274
rect 17224 41210 17276 41216
rect 17420 40769 17448 43710
rect 17512 43450 17540 47126
rect 17592 46368 17644 46374
rect 17592 46310 17644 46316
rect 17604 45966 17632 46310
rect 17592 45960 17644 45966
rect 17592 45902 17644 45908
rect 17592 44804 17644 44810
rect 17592 44746 17644 44752
rect 17604 44470 17632 44746
rect 17592 44464 17644 44470
rect 17592 44406 17644 44412
rect 17696 43858 17724 47942
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 18236 47796 18288 47802
rect 18432 47784 18460 53926
rect 18524 53786 18552 54130
rect 18512 53780 18564 53786
rect 18512 53722 18564 53728
rect 18800 53106 18828 56200
rect 19168 53582 19196 56200
rect 19536 54262 19564 56200
rect 19524 54256 19576 54262
rect 19524 54198 19576 54204
rect 19708 54188 19760 54194
rect 19708 54130 19760 54136
rect 19340 53984 19392 53990
rect 19340 53926 19392 53932
rect 19156 53576 19208 53582
rect 19156 53518 19208 53524
rect 19168 53242 19196 53518
rect 19156 53236 19208 53242
rect 19156 53178 19208 53184
rect 18788 53100 18840 53106
rect 18788 53042 18840 53048
rect 18880 52896 18932 52902
rect 18880 52838 18932 52844
rect 18696 48272 18748 48278
rect 18696 48214 18748 48220
rect 18288 47756 18460 47784
rect 18236 47738 18288 47744
rect 17776 47456 17828 47462
rect 17776 47398 17828 47404
rect 17788 44334 17816 47398
rect 18248 47258 18276 47738
rect 18236 47252 18288 47258
rect 18236 47194 18288 47200
rect 18512 47252 18564 47258
rect 18512 47194 18564 47200
rect 18248 47161 18276 47194
rect 18234 47152 18290 47161
rect 18234 47087 18290 47096
rect 18524 46986 18552 47194
rect 18604 47048 18656 47054
rect 18604 46990 18656 46996
rect 18512 46980 18564 46986
rect 18512 46922 18564 46928
rect 17868 46912 17920 46918
rect 17868 46854 17920 46860
rect 17880 46646 17908 46854
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17868 46640 17920 46646
rect 17868 46582 17920 46588
rect 18616 46578 18644 46990
rect 18604 46572 18656 46578
rect 18604 46514 18656 46520
rect 18328 46504 18380 46510
rect 18328 46446 18380 46452
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18340 45626 18368 46446
rect 18328 45620 18380 45626
rect 18328 45562 18380 45568
rect 18328 45484 18380 45490
rect 18328 45426 18380 45432
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17776 44328 17828 44334
rect 17776 44270 17828 44276
rect 18340 44198 18368 45426
rect 18328 44192 18380 44198
rect 18328 44134 18380 44140
rect 17684 43852 17736 43858
rect 17684 43794 17736 43800
rect 17776 43648 17828 43654
rect 17776 43590 17828 43596
rect 17500 43444 17552 43450
rect 17500 43386 17552 43392
rect 17788 43314 17816 43590
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17776 43308 17828 43314
rect 17776 43250 17828 43256
rect 17500 42900 17552 42906
rect 17500 42842 17552 42848
rect 17406 40760 17462 40769
rect 17316 40724 17368 40730
rect 17406 40695 17462 40704
rect 17316 40666 17368 40672
rect 17328 40050 17356 40666
rect 17408 40588 17460 40594
rect 17408 40530 17460 40536
rect 17316 40044 17368 40050
rect 17316 39986 17368 39992
rect 17132 39500 17184 39506
rect 17132 39442 17184 39448
rect 17328 39030 17356 39986
rect 17420 39438 17448 40530
rect 17408 39432 17460 39438
rect 17408 39374 17460 39380
rect 17316 39024 17368 39030
rect 17316 38966 17368 38972
rect 17420 38350 17448 39374
rect 17408 38344 17460 38350
rect 17408 38286 17460 38292
rect 17224 38208 17276 38214
rect 17224 38150 17276 38156
rect 16948 37868 17000 37874
rect 16948 37810 17000 37816
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16856 34128 16908 34134
rect 16776 34088 16856 34116
rect 16856 34070 16908 34076
rect 16684 34020 16804 34048
rect 16396 33312 16448 33318
rect 16396 33254 16448 33260
rect 16408 31754 16436 33254
rect 16672 32904 16724 32910
rect 16672 32846 16724 32852
rect 16580 32768 16632 32774
rect 16580 32710 16632 32716
rect 16408 31726 16528 31754
rect 16304 31476 16356 31482
rect 16304 31418 16356 31424
rect 16316 31210 16344 31418
rect 16304 31204 16356 31210
rect 16304 31146 16356 31152
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16316 30394 16344 30534
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16394 28112 16450 28121
rect 16394 28047 16450 28056
rect 16304 27940 16356 27946
rect 16304 27882 16356 27888
rect 15948 23208 16252 23236
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15948 22794 15976 23208
rect 16316 23066 16344 27882
rect 16408 27878 16436 28047
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16394 26616 16450 26625
rect 16394 26551 16396 26560
rect 16448 26551 16450 26560
rect 16396 26522 16448 26528
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16408 24138 16436 24754
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 15672 22766 15976 22794
rect 16132 23038 16344 23066
rect 15672 22030 15700 22766
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15856 22166 15884 22578
rect 15844 22160 15896 22166
rect 15844 22102 15896 22108
rect 16132 22094 16160 23038
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 15948 22066 16160 22094
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15764 21146 15792 21422
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15948 21078 15976 22066
rect 15936 21072 15988 21078
rect 15936 21014 15988 21020
rect 15750 20360 15806 20369
rect 15750 20295 15752 20304
rect 15804 20295 15806 20304
rect 15752 20266 15804 20272
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15672 15026 15700 17070
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14414 15608 14758
rect 15672 14618 15700 14962
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15304 14062 15516 14090
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15304 12434 15332 13942
rect 15488 13682 15516 14062
rect 15580 13870 15608 14350
rect 15764 14006 15792 20266
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15948 18290 15976 18566
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15488 13654 15608 13682
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15212 12406 15332 12434
rect 15212 11642 15240 12406
rect 15212 11614 15332 11642
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 10742 15240 11494
rect 15304 11354 15332 11614
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15396 10606 15424 13398
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15488 7478 15516 12922
rect 15580 12918 15608 13654
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 11642 15608 12718
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15672 11830 15700 12174
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15580 11614 15700 11642
rect 15672 11218 15700 11614
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10810 15608 10950
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15856 4078 15884 13806
rect 15948 7818 15976 18226
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16040 13297 16068 14418
rect 16132 13734 16160 19246
rect 16224 18902 16252 22918
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16408 18766 16436 23462
rect 16500 21962 16528 31726
rect 16592 31686 16620 32710
rect 16684 31754 16712 32846
rect 16672 31748 16724 31754
rect 16672 31690 16724 31696
rect 16580 31680 16632 31686
rect 16580 31622 16632 31628
rect 16672 31204 16724 31210
rect 16672 31146 16724 31152
rect 16684 30938 16712 31146
rect 16672 30932 16724 30938
rect 16672 30874 16724 30880
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16592 28626 16620 29786
rect 16776 29696 16804 34020
rect 16856 33992 16908 33998
rect 16856 33934 16908 33940
rect 16868 32298 16896 33934
rect 16960 33522 16988 37810
rect 17236 37330 17264 38150
rect 17316 37664 17368 37670
rect 17420 37618 17448 38286
rect 17368 37612 17448 37618
rect 17316 37606 17448 37612
rect 17328 37590 17448 37606
rect 17224 37324 17276 37330
rect 17224 37266 17276 37272
rect 17316 37256 17368 37262
rect 17316 37198 17368 37204
rect 17224 37120 17276 37126
rect 17224 37062 17276 37068
rect 17236 36922 17264 37062
rect 17224 36916 17276 36922
rect 17224 36858 17276 36864
rect 17328 36310 17356 37198
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 17316 36304 17368 36310
rect 17316 36246 17368 36252
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 17236 35154 17264 35634
rect 17224 35148 17276 35154
rect 17224 35090 17276 35096
rect 17224 35012 17276 35018
rect 17224 34954 17276 34960
rect 17236 34746 17264 34954
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 17040 34672 17092 34678
rect 17040 34614 17092 34620
rect 16948 33516 17000 33522
rect 16948 33458 17000 33464
rect 16948 32428 17000 32434
rect 16948 32370 17000 32376
rect 16856 32292 16908 32298
rect 16856 32234 16908 32240
rect 16960 31754 16988 32370
rect 16684 29668 16804 29696
rect 16868 31726 16988 31754
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16592 27470 16620 28154
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 16592 26042 16620 27406
rect 16684 26518 16712 29668
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16776 29073 16804 29514
rect 16868 29170 16896 31726
rect 16948 31476 17000 31482
rect 16948 31418 17000 31424
rect 16960 30802 16988 31418
rect 16948 30796 17000 30802
rect 16948 30738 17000 30744
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16960 29510 16988 30194
rect 16948 29504 17000 29510
rect 16948 29446 17000 29452
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16762 29064 16818 29073
rect 16762 28999 16764 29008
rect 16816 28999 16818 29008
rect 16764 28970 16816 28976
rect 16854 27704 16910 27713
rect 16854 27639 16856 27648
rect 16908 27639 16910 27648
rect 16856 27610 16908 27616
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16672 26512 16724 26518
rect 16672 26454 16724 26460
rect 16776 26314 16804 26862
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 16764 26308 16816 26314
rect 16764 26250 16816 26256
rect 16776 26217 16804 26250
rect 16762 26208 16818 26217
rect 16762 26143 16818 26152
rect 16580 26036 16632 26042
rect 16580 25978 16632 25984
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16776 24954 16804 25162
rect 16764 24948 16816 24954
rect 16764 24890 16816 24896
rect 16580 24608 16632 24614
rect 16580 24550 16632 24556
rect 16592 23866 16620 24550
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16580 23588 16632 23594
rect 16580 23530 16632 23536
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16500 19990 16528 20538
rect 16488 19984 16540 19990
rect 16486 19952 16488 19961
rect 16540 19952 16542 19961
rect 16486 19887 16542 19896
rect 16592 19854 16620 23530
rect 16776 23322 16804 24890
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16684 21894 16712 22374
rect 16776 22030 16804 22918
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16868 21690 16896 26726
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16868 20874 16896 21286
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16960 20806 16988 29446
rect 17052 29238 17080 34614
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17236 32774 17264 33050
rect 17224 32768 17276 32774
rect 17224 32710 17276 32716
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 17144 30938 17172 32302
rect 17236 31754 17264 32710
rect 17328 32570 17356 36246
rect 17420 33658 17448 37062
rect 17512 36718 17540 42842
rect 17592 41812 17644 41818
rect 17592 41754 17644 41760
rect 17604 41478 17632 41754
rect 17592 41472 17644 41478
rect 17592 41414 17644 41420
rect 17788 41414 17816 43250
rect 17868 43240 17920 43246
rect 17868 43182 17920 43188
rect 17880 41682 17908 43182
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17868 41676 17920 41682
rect 17868 41618 17920 41624
rect 17696 41386 17816 41414
rect 17592 40928 17644 40934
rect 17592 40870 17644 40876
rect 17500 36712 17552 36718
rect 17500 36654 17552 36660
rect 17500 35760 17552 35766
rect 17500 35702 17552 35708
rect 17512 35290 17540 35702
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17498 34504 17554 34513
rect 17498 34439 17554 34448
rect 17408 33652 17460 33658
rect 17408 33594 17460 33600
rect 17408 33040 17460 33046
rect 17408 32982 17460 32988
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 17420 32434 17448 32982
rect 17512 32978 17540 34439
rect 17500 32972 17552 32978
rect 17500 32914 17552 32920
rect 17604 32910 17632 40870
rect 17696 39914 17724 41386
rect 17880 40458 17908 41618
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 18340 41070 18368 44134
rect 18420 43172 18472 43178
rect 18420 43114 18472 43120
rect 18432 41274 18460 43114
rect 18512 41472 18564 41478
rect 18512 41414 18564 41420
rect 18420 41268 18472 41274
rect 18420 41210 18472 41216
rect 18328 41064 18380 41070
rect 18328 41006 18380 41012
rect 18524 40594 18552 41414
rect 18708 41274 18736 48214
rect 18788 48136 18840 48142
rect 18788 48078 18840 48084
rect 18800 47122 18828 48078
rect 18788 47116 18840 47122
rect 18788 47058 18840 47064
rect 18800 46714 18828 47058
rect 18892 46986 18920 52838
rect 18972 49088 19024 49094
rect 18972 49030 19024 49036
rect 18880 46980 18932 46986
rect 18880 46922 18932 46928
rect 18788 46708 18840 46714
rect 18788 46650 18840 46656
rect 18984 45554 19012 49030
rect 19064 47728 19116 47734
rect 19116 47676 19196 47682
rect 19064 47670 19196 47676
rect 19076 47654 19196 47670
rect 19168 46714 19196 47654
rect 19352 47258 19380 53926
rect 19616 53440 19668 53446
rect 19616 53382 19668 53388
rect 19524 48000 19576 48006
rect 19524 47942 19576 47948
rect 19536 47734 19564 47942
rect 19524 47728 19576 47734
rect 19524 47670 19576 47676
rect 19524 47456 19576 47462
rect 19524 47398 19576 47404
rect 19340 47252 19392 47258
rect 19340 47194 19392 47200
rect 19246 47152 19302 47161
rect 19352 47138 19380 47194
rect 19302 47110 19380 47138
rect 19246 47087 19302 47096
rect 19156 46708 19208 46714
rect 19156 46650 19208 46656
rect 19536 46458 19564 47398
rect 19628 47054 19656 53382
rect 19720 53242 19748 54130
rect 19904 53582 19932 56200
rect 19892 53576 19944 53582
rect 19892 53518 19944 53524
rect 19708 53236 19760 53242
rect 19708 53178 19760 53184
rect 20272 53106 20300 56200
rect 20640 55214 20668 56200
rect 20640 55186 20760 55214
rect 20732 54194 20760 55186
rect 20720 54188 20772 54194
rect 20720 54130 20772 54136
rect 20444 53984 20496 53990
rect 20444 53926 20496 53932
rect 20260 53100 20312 53106
rect 20260 53042 20312 53048
rect 20076 52896 20128 52902
rect 20076 52838 20128 52844
rect 19800 49768 19852 49774
rect 19800 49710 19852 49716
rect 19616 47048 19668 47054
rect 19614 47016 19616 47025
rect 19668 47016 19670 47025
rect 19614 46951 19670 46960
rect 19444 46430 19564 46458
rect 19248 45892 19300 45898
rect 19248 45834 19300 45840
rect 18800 45526 19012 45554
rect 18800 42362 18828 45526
rect 19156 45280 19208 45286
rect 19156 45222 19208 45228
rect 18880 44872 18932 44878
rect 18880 44814 18932 44820
rect 18892 43110 18920 44814
rect 19168 44402 19196 45222
rect 19156 44396 19208 44402
rect 19156 44338 19208 44344
rect 18880 43104 18932 43110
rect 18880 43046 18932 43052
rect 18788 42356 18840 42362
rect 18788 42298 18840 42304
rect 18696 41268 18748 41274
rect 18696 41210 18748 41216
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18512 40588 18564 40594
rect 18512 40530 18564 40536
rect 17868 40452 17920 40458
rect 17868 40394 17920 40400
rect 18512 40452 18564 40458
rect 18512 40394 18564 40400
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17776 40112 17828 40118
rect 17776 40054 17828 40060
rect 18328 40112 18380 40118
rect 18328 40054 18380 40060
rect 17684 39908 17736 39914
rect 17684 39850 17736 39856
rect 17696 38758 17724 39850
rect 17684 38752 17736 38758
rect 17684 38694 17736 38700
rect 17682 38584 17738 38593
rect 17682 38519 17738 38528
rect 17696 33386 17724 38519
rect 17788 38350 17816 40054
rect 17868 39568 17920 39574
rect 17868 39510 17920 39516
rect 17880 39098 17908 39510
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17868 39092 17920 39098
rect 17868 39034 17920 39040
rect 18340 38554 18368 40054
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18328 38548 18380 38554
rect 18328 38490 18380 38496
rect 17776 38344 17828 38350
rect 17776 38286 17828 38292
rect 18328 38344 18380 38350
rect 18328 38286 18380 38292
rect 17960 38208 18012 38214
rect 17788 38168 17960 38196
rect 17788 37806 17816 38168
rect 17960 38150 18012 38156
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17776 37800 17828 37806
rect 17776 37742 17828 37748
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 17788 35630 17816 36314
rect 17776 35624 17828 35630
rect 17776 35566 17828 35572
rect 17788 34542 17816 35566
rect 17776 34536 17828 34542
rect 17776 34478 17828 34484
rect 17776 33856 17828 33862
rect 17776 33798 17828 33804
rect 17684 33380 17736 33386
rect 17684 33322 17736 33328
rect 17682 33280 17738 33289
rect 17682 33215 17738 33224
rect 17696 33114 17724 33215
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17500 32768 17552 32774
rect 17500 32710 17552 32716
rect 17512 32570 17540 32710
rect 17500 32564 17552 32570
rect 17500 32506 17552 32512
rect 17788 32502 17816 33798
rect 17776 32496 17828 32502
rect 17776 32438 17828 32444
rect 17408 32428 17460 32434
rect 17408 32370 17460 32376
rect 17500 32292 17552 32298
rect 17500 32234 17552 32240
rect 17408 31952 17460 31958
rect 17408 31894 17460 31900
rect 17236 31726 17356 31754
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17132 30932 17184 30938
rect 17132 30874 17184 30880
rect 17144 30326 17172 30874
rect 17132 30320 17184 30326
rect 17132 30262 17184 30268
rect 17132 30116 17184 30122
rect 17132 30058 17184 30064
rect 17040 29232 17092 29238
rect 17040 29174 17092 29180
rect 17040 28416 17092 28422
rect 17040 28358 17092 28364
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16960 20346 16988 20742
rect 17052 20466 17080 28358
rect 17144 26489 17172 30058
rect 17236 29714 17264 31282
rect 17224 29708 17276 29714
rect 17224 29650 17276 29656
rect 17130 26480 17186 26489
rect 17130 26415 17186 26424
rect 17144 26246 17172 26415
rect 17132 26240 17184 26246
rect 17132 26182 17184 26188
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17144 24682 17172 25842
rect 17236 25362 17264 29650
rect 17328 27033 17356 31726
rect 17420 30394 17448 31894
rect 17512 31686 17540 32234
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 17512 30870 17540 31622
rect 17500 30864 17552 30870
rect 17500 30806 17552 30812
rect 17408 30388 17460 30394
rect 17408 30330 17460 30336
rect 17420 30161 17448 30330
rect 17500 30184 17552 30190
rect 17406 30152 17462 30161
rect 17500 30126 17552 30132
rect 17406 30087 17462 30096
rect 17512 29170 17540 30126
rect 17500 29164 17552 29170
rect 17420 29124 17500 29152
rect 17420 27606 17448 29124
rect 17500 29106 17552 29112
rect 17500 28960 17552 28966
rect 17500 28902 17552 28908
rect 17512 28558 17540 28902
rect 17604 28626 17632 32166
rect 17684 31816 17736 31822
rect 17684 31758 17736 31764
rect 17696 29850 17724 31758
rect 17776 31680 17828 31686
rect 17776 31622 17828 31628
rect 17788 31210 17816 31622
rect 17776 31204 17828 31210
rect 17776 31146 17828 31152
rect 17880 30938 17908 37266
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 18340 35494 18368 38286
rect 18432 37942 18460 39238
rect 18420 37936 18472 37942
rect 18420 37878 18472 37884
rect 18420 36032 18472 36038
rect 18420 35974 18472 35980
rect 18432 35766 18460 35974
rect 18420 35760 18472 35766
rect 18420 35702 18472 35708
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 18420 35148 18472 35154
rect 18420 35090 18472 35096
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 18340 33318 18368 34546
rect 18432 34202 18460 35090
rect 18420 34196 18472 34202
rect 18420 34138 18472 34144
rect 18328 33312 18380 33318
rect 18524 33266 18552 40394
rect 18616 39642 18644 41074
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18604 39636 18656 39642
rect 18604 39578 18656 39584
rect 18604 39296 18656 39302
rect 18604 39238 18656 39244
rect 18616 39030 18644 39238
rect 18604 39024 18656 39030
rect 18604 38966 18656 38972
rect 18604 38480 18656 38486
rect 18604 38422 18656 38428
rect 18616 37194 18644 38422
rect 18604 37188 18656 37194
rect 18604 37130 18656 37136
rect 18616 34746 18644 37130
rect 18604 34740 18656 34746
rect 18604 34682 18656 34688
rect 18708 34592 18736 40870
rect 18800 37262 18828 42298
rect 18892 39982 18920 43046
rect 18972 42016 19024 42022
rect 18972 41958 19024 41964
rect 18984 41206 19012 41958
rect 19064 41268 19116 41274
rect 19064 41210 19116 41216
rect 18972 41200 19024 41206
rect 18972 41142 19024 41148
rect 18984 40594 19012 41142
rect 18972 40588 19024 40594
rect 18972 40530 19024 40536
rect 18972 40384 19024 40390
rect 18972 40326 19024 40332
rect 18880 39976 18932 39982
rect 18880 39918 18932 39924
rect 18880 38820 18932 38826
rect 18880 38762 18932 38768
rect 18892 38350 18920 38762
rect 18880 38344 18932 38350
rect 18880 38286 18932 38292
rect 18892 37942 18920 38286
rect 18880 37936 18932 37942
rect 18880 37878 18932 37884
rect 18880 37460 18932 37466
rect 18880 37402 18932 37408
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 18892 37126 18920 37402
rect 18880 37120 18932 37126
rect 18880 37062 18932 37068
rect 18708 34564 18828 34592
rect 18604 34468 18656 34474
rect 18604 34410 18656 34416
rect 18696 34468 18748 34474
rect 18696 34410 18748 34416
rect 18328 33254 18380 33260
rect 18432 33238 18552 33266
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18328 32020 18380 32026
rect 18328 31962 18380 31968
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 17868 30796 17920 30802
rect 17868 30738 17920 30744
rect 17880 30666 17908 30738
rect 18340 30682 18368 31962
rect 18432 31958 18460 33238
rect 18512 33108 18564 33114
rect 18512 33050 18564 33056
rect 18420 31952 18472 31958
rect 18420 31894 18472 31900
rect 17868 30660 17920 30666
rect 18340 30654 18460 30682
rect 17868 30602 17920 30608
rect 17776 30388 17828 30394
rect 17776 30330 17828 30336
rect 17684 29844 17736 29850
rect 17684 29786 17736 29792
rect 17788 29102 17816 30330
rect 17880 29578 17908 30602
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18340 30394 18368 30534
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18432 30138 18460 30654
rect 18340 30110 18460 30138
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 18064 29714 18092 29786
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 17868 29572 17920 29578
rect 17868 29514 17920 29520
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17776 29096 17828 29102
rect 17776 29038 17828 29044
rect 18340 29034 18368 30110
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18432 29714 18460 29990
rect 18420 29708 18472 29714
rect 18420 29650 18472 29656
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 18328 29028 18380 29034
rect 18328 28970 18380 28976
rect 17592 28620 17644 28626
rect 17592 28562 17644 28568
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 18248 28422 18276 28562
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17684 28416 17736 28422
rect 17684 28358 17736 28364
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 17500 28144 17552 28150
rect 17500 28086 17552 28092
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 17512 27418 17540 28086
rect 17604 27538 17632 28358
rect 17696 28218 17724 28358
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17684 28212 17736 28218
rect 17684 28154 17736 28160
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 17866 28112 17922 28121
rect 17866 28047 17868 28056
rect 17920 28047 17922 28056
rect 17868 28018 17920 28024
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 17592 27532 17644 27538
rect 17592 27474 17644 27480
rect 17420 27390 17540 27418
rect 17314 27024 17370 27033
rect 17314 26959 17370 26968
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 17328 26790 17356 26862
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 17316 26512 17368 26518
rect 17316 26454 17368 26460
rect 17224 25356 17276 25362
rect 17224 25298 17276 25304
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17144 24274 17172 24618
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 17144 22642 17172 24210
rect 17132 22636 17184 22642
rect 17132 22578 17184 22584
rect 17328 22094 17356 26454
rect 17420 23746 17448 27390
rect 17500 27328 17552 27334
rect 17500 27270 17552 27276
rect 17512 23866 17540 27270
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17604 26450 17632 26930
rect 17696 26926 17724 27542
rect 18248 27538 18276 28154
rect 18340 27962 18368 28970
rect 18432 28966 18460 29514
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18420 28756 18472 28762
rect 18420 28698 18472 28704
rect 18432 28626 18460 28698
rect 18420 28620 18472 28626
rect 18420 28562 18472 28568
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 28218 18460 28358
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18340 27934 18460 27962
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 18236 27532 18288 27538
rect 18236 27474 18288 27480
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17682 26752 17738 26761
rect 17682 26687 17738 26696
rect 17592 26444 17644 26450
rect 17592 26386 17644 26392
rect 17696 24834 17724 26687
rect 17788 26353 17816 26930
rect 17774 26344 17830 26353
rect 17774 26279 17830 26288
rect 17788 26246 17816 26279
rect 17776 26240 17828 26246
rect 17776 26182 17828 26188
rect 17788 25226 17816 26182
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 17604 24806 17724 24834
rect 17604 24596 17632 24806
rect 17684 24744 17736 24750
rect 17880 24698 17908 27406
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26042 18368 27814
rect 18432 27130 18460 27934
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 17736 24692 17908 24698
rect 17684 24686 17908 24692
rect 17696 24670 17908 24686
rect 17604 24568 17816 24596
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17420 23718 17724 23746
rect 17408 23248 17460 23254
rect 17408 23190 17460 23196
rect 17236 22066 17356 22094
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16960 20318 17080 20346
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16500 18970 16528 19110
rect 16684 18970 16712 19314
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16684 18766 16712 18906
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16960 17762 16988 20198
rect 16776 17734 16988 17762
rect 16776 17678 16804 17734
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16408 16833 16436 17070
rect 16394 16824 16450 16833
rect 16394 16759 16396 16768
rect 16448 16759 16450 16768
rect 16396 16730 16448 16736
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16500 15910 16528 16458
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 16224 15162 16252 15370
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16224 14618 16344 14634
rect 16224 14612 16356 14618
rect 16224 14606 16304 14612
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16026 13288 16082 13297
rect 16026 13223 16082 13232
rect 16040 12442 16068 13223
rect 16028 12436 16080 12442
rect 16224 12434 16252 14606
rect 16304 14554 16356 14560
rect 16500 14346 16528 15846
rect 16684 14958 16712 17478
rect 16868 17338 16896 17614
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 12850 16436 14214
rect 16500 13190 16528 14282
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16028 12378 16080 12384
rect 16132 12406 16252 12434
rect 16132 11082 16160 12406
rect 16500 12238 16528 13126
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10742 16436 10950
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16316 4146 16344 7210
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 16132 3670 16160 4082
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14568 800 14596 2450
rect 14936 800 14964 3402
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15304 800 15332 2450
rect 15672 800 15700 2926
rect 16040 800 16068 3538
rect 16408 800 16436 3946
rect 16500 3058 16528 11562
rect 16592 3534 16620 14826
rect 16960 13954 16988 17734
rect 17052 17524 17080 20318
rect 17144 19786 17172 20742
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 17236 18834 17264 22066
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17144 17678 17172 18770
rect 17328 17678 17356 21830
rect 17420 19378 17448 23190
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17512 21622 17540 22986
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17512 21350 17540 21558
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17696 21162 17724 23718
rect 17788 23186 17816 24568
rect 17880 24206 17908 24670
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17512 21134 17724 21162
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17052 17496 17356 17524
rect 17224 15700 17276 15706
rect 16776 13926 16988 13954
rect 17052 15660 17224 15688
rect 16776 8974 16804 13926
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16868 3534 16896 12650
rect 17052 12434 17080 15660
rect 17224 15642 17276 15648
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17144 12986 17172 13806
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 16960 12406 17080 12434
rect 16960 11830 16988 12406
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 800 16804 2790
rect 17052 2446 17080 9930
rect 17236 6798 17264 14894
rect 17328 13394 17356 17496
rect 17512 16182 17540 21134
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17604 15910 17632 16594
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15502 17632 15846
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17498 15192 17554 15201
rect 17498 15127 17500 15136
rect 17552 15127 17554 15136
rect 17500 15098 17552 15104
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17420 13462 17448 14418
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17328 11694 17356 12106
rect 17420 11744 17448 13398
rect 17500 13320 17552 13326
rect 17498 13288 17500 13297
rect 17552 13288 17554 13297
rect 17498 13223 17554 13232
rect 17500 11756 17552 11762
rect 17420 11716 17500 11744
rect 17500 11698 17552 11704
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17144 800 17172 2858
rect 17328 2038 17356 11630
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17316 2032 17368 2038
rect 17316 1974 17368 1980
rect 17512 800 17540 4014
rect 17696 3058 17724 20198
rect 17788 16538 17816 23122
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17972 22166 18000 22714
rect 18340 22166 18368 25638
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 18328 22160 18380 22166
rect 18328 22102 18380 22108
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18340 21554 18368 21830
rect 18432 21690 18460 22034
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17880 19786 17908 21286
rect 17972 21010 18000 21422
rect 18524 21146 18552 33050
rect 18616 31482 18644 34410
rect 18708 31482 18736 34410
rect 18800 32570 18828 34564
rect 18892 33114 18920 37062
rect 18984 36650 19012 40326
rect 19076 37466 19104 41210
rect 19168 41070 19196 44338
rect 19156 41064 19208 41070
rect 19156 41006 19208 41012
rect 19168 38282 19196 41006
rect 19156 38276 19208 38282
rect 19156 38218 19208 38224
rect 19064 37460 19116 37466
rect 19064 37402 19116 37408
rect 18972 36644 19024 36650
rect 18972 36586 19024 36592
rect 19260 36564 19288 45834
rect 19340 43920 19392 43926
rect 19340 43862 19392 43868
rect 19352 38554 19380 43862
rect 19444 43450 19472 46430
rect 19524 46368 19576 46374
rect 19524 46310 19576 46316
rect 19536 45014 19564 46310
rect 19524 45008 19576 45014
rect 19524 44950 19576 44956
rect 19616 44192 19668 44198
rect 19616 44134 19668 44140
rect 19432 43444 19484 43450
rect 19432 43386 19484 43392
rect 19444 42022 19472 43386
rect 19628 43246 19656 44134
rect 19708 43648 19760 43654
rect 19708 43590 19760 43596
rect 19720 43450 19748 43590
rect 19708 43444 19760 43450
rect 19708 43386 19760 43392
rect 19524 43240 19576 43246
rect 19524 43182 19576 43188
rect 19616 43240 19668 43246
rect 19616 43182 19668 43188
rect 19536 43110 19564 43182
rect 19524 43104 19576 43110
rect 19524 43046 19576 43052
rect 19720 42906 19748 43386
rect 19708 42900 19760 42906
rect 19708 42842 19760 42848
rect 19616 42832 19668 42838
rect 19616 42774 19668 42780
rect 19432 42016 19484 42022
rect 19432 41958 19484 41964
rect 19444 41682 19472 41958
rect 19432 41676 19484 41682
rect 19432 41618 19484 41624
rect 19432 40928 19484 40934
rect 19432 40870 19484 40876
rect 19444 40186 19472 40870
rect 19524 40384 19576 40390
rect 19524 40326 19576 40332
rect 19432 40180 19484 40186
rect 19432 40122 19484 40128
rect 19432 39500 19484 39506
rect 19432 39442 19484 39448
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 19444 37890 19472 39442
rect 19536 38010 19564 40326
rect 19628 38418 19656 42774
rect 19812 42634 19840 49710
rect 19892 47184 19944 47190
rect 19892 47126 19944 47132
rect 19800 42628 19852 42634
rect 19800 42570 19852 42576
rect 19800 42356 19852 42362
rect 19800 42298 19852 42304
rect 19708 38956 19760 38962
rect 19708 38898 19760 38904
rect 19616 38412 19668 38418
rect 19616 38354 19668 38360
rect 19524 38004 19576 38010
rect 19524 37946 19576 37952
rect 19444 37862 19564 37890
rect 19432 37732 19484 37738
rect 19432 37674 19484 37680
rect 19340 37188 19392 37194
rect 19340 37130 19392 37136
rect 19076 36536 19288 36564
rect 18972 33312 19024 33318
rect 18972 33254 19024 33260
rect 18880 33108 18932 33114
rect 18880 33050 18932 33056
rect 18788 32564 18840 32570
rect 18788 32506 18840 32512
rect 18880 32292 18932 32298
rect 18880 32234 18932 32240
rect 18892 32042 18920 32234
rect 18800 32014 18920 32042
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18696 31476 18748 31482
rect 18696 31418 18748 31424
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18616 23202 18644 27950
rect 18708 25770 18736 31282
rect 18800 28778 18828 32014
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 18892 30734 18920 31690
rect 18984 31278 19012 33254
rect 18972 31272 19024 31278
rect 18972 31214 19024 31220
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 18892 29714 18920 30670
rect 18970 30424 19026 30433
rect 18970 30359 19026 30368
rect 18880 29708 18932 29714
rect 18880 29650 18932 29656
rect 18800 28750 18920 28778
rect 18984 28762 19012 30359
rect 19076 29510 19104 36536
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19260 35290 19288 35634
rect 19156 35284 19208 35290
rect 19156 35226 19208 35232
rect 19248 35284 19300 35290
rect 19248 35226 19300 35232
rect 19168 32434 19196 35226
rect 19260 34950 19288 35226
rect 19352 35086 19380 37130
rect 19444 35834 19472 37674
rect 19536 36718 19564 37862
rect 19616 37120 19668 37126
rect 19616 37062 19668 37068
rect 19628 36854 19656 37062
rect 19720 36922 19748 38898
rect 19708 36916 19760 36922
rect 19708 36858 19760 36864
rect 19616 36848 19668 36854
rect 19616 36790 19668 36796
rect 19524 36712 19576 36718
rect 19524 36654 19576 36660
rect 19524 36576 19576 36582
rect 19524 36518 19576 36524
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19248 34944 19300 34950
rect 19248 34886 19300 34892
rect 19260 34066 19288 34886
rect 19248 34060 19300 34066
rect 19248 34002 19300 34008
rect 19260 33590 19288 34002
rect 19248 33584 19300 33590
rect 19248 33526 19300 33532
rect 19352 33436 19380 35022
rect 19430 34640 19486 34649
rect 19430 34575 19432 34584
rect 19484 34575 19486 34584
rect 19432 34546 19484 34552
rect 19432 33448 19484 33454
rect 19352 33408 19432 33436
rect 19352 33130 19380 33408
rect 19432 33390 19484 33396
rect 19260 33102 19380 33130
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19156 32224 19208 32230
rect 19156 32166 19208 32172
rect 19064 29504 19116 29510
rect 19064 29446 19116 29452
rect 19064 29164 19116 29170
rect 19064 29106 19116 29112
rect 18788 28688 18840 28694
rect 18788 28630 18840 28636
rect 18696 25764 18748 25770
rect 18696 25706 18748 25712
rect 18696 25356 18748 25362
rect 18696 25298 18748 25304
rect 18708 24750 18736 25298
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18708 24410 18736 24686
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18708 23322 18736 24346
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18616 23174 18736 23202
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18616 22098 18644 23054
rect 18708 22982 18736 23174
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18708 22574 18736 22918
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18708 21672 18736 22102
rect 18616 21644 18736 21672
rect 18616 21486 18644 21644
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18800 21298 18828 28630
rect 18892 28014 18920 28750
rect 18972 28756 19024 28762
rect 18972 28698 19024 28704
rect 19076 28626 19104 29106
rect 19064 28620 19116 28626
rect 19064 28562 19116 28568
rect 18972 28212 19024 28218
rect 18972 28154 19024 28160
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18880 27872 18932 27878
rect 18878 27840 18880 27849
rect 18932 27840 18934 27849
rect 18878 27775 18934 27784
rect 18880 27464 18932 27470
rect 18880 27406 18932 27412
rect 18892 25362 18920 27406
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22094 18920 22918
rect 18984 22522 19012 28154
rect 19076 26042 19104 28562
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 19076 23730 19104 25978
rect 19168 25974 19196 32166
rect 19260 31754 19288 33102
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19352 32366 19380 32710
rect 19536 32502 19564 36518
rect 19812 36242 19840 42298
rect 19904 41274 19932 47126
rect 20088 47122 20116 52838
rect 20168 47660 20220 47666
rect 20168 47602 20220 47608
rect 20180 47122 20208 47602
rect 20076 47116 20128 47122
rect 20076 47058 20128 47064
rect 20168 47116 20220 47122
rect 20168 47058 20220 47064
rect 20180 45082 20208 47058
rect 20456 45898 20484 53926
rect 20628 53712 20680 53718
rect 20628 53654 20680 53660
rect 20536 53440 20588 53446
rect 20536 53382 20588 53388
rect 20548 47258 20576 53382
rect 20536 47252 20588 47258
rect 20536 47194 20588 47200
rect 20444 45892 20496 45898
rect 20444 45834 20496 45840
rect 20260 45824 20312 45830
rect 20260 45766 20312 45772
rect 20168 45076 20220 45082
rect 20168 45018 20220 45024
rect 20168 44396 20220 44402
rect 20168 44338 20220 44344
rect 19984 42560 20036 42566
rect 19984 42502 20036 42508
rect 19996 41274 20024 42502
rect 20076 42084 20128 42090
rect 20076 42026 20128 42032
rect 19892 41268 19944 41274
rect 19892 41210 19944 41216
rect 19984 41268 20036 41274
rect 19984 41210 20036 41216
rect 19982 41168 20038 41177
rect 19892 41132 19944 41138
rect 19982 41103 20038 41112
rect 19892 41074 19944 41080
rect 19904 40458 19932 41074
rect 19892 40452 19944 40458
rect 19892 40394 19944 40400
rect 19996 40338 20024 41103
rect 19904 40310 20024 40338
rect 19800 36236 19852 36242
rect 19800 36178 19852 36184
rect 19616 36032 19668 36038
rect 19616 35974 19668 35980
rect 19628 33658 19656 35974
rect 19708 34128 19760 34134
rect 19708 34070 19760 34076
rect 19720 33658 19748 34070
rect 19904 33946 19932 40310
rect 19984 40180 20036 40186
rect 19984 40122 20036 40128
rect 19996 40089 20024 40122
rect 19982 40080 20038 40089
rect 19982 40015 20038 40024
rect 20088 38418 20116 42026
rect 20180 42022 20208 44338
rect 20272 42770 20300 45766
rect 20548 45554 20576 47194
rect 20640 46034 20668 53654
rect 21008 53582 21036 56200
rect 21376 54194 21404 56200
rect 21180 54188 21232 54194
rect 21180 54130 21232 54136
rect 21364 54188 21416 54194
rect 21364 54130 21416 54136
rect 20996 53576 21048 53582
rect 20996 53518 21048 53524
rect 21008 53242 21036 53518
rect 21192 53242 21220 54130
rect 21640 53984 21692 53990
rect 21640 53926 21692 53932
rect 21272 53440 21324 53446
rect 21272 53382 21324 53388
rect 20996 53236 21048 53242
rect 20996 53178 21048 53184
rect 21180 53236 21232 53242
rect 21180 53178 21232 53184
rect 20720 47456 20772 47462
rect 20720 47398 20772 47404
rect 20628 46028 20680 46034
rect 20628 45970 20680 45976
rect 20732 45558 20760 47398
rect 21180 46504 21232 46510
rect 21180 46446 21232 46452
rect 20456 45526 20576 45554
rect 20628 45552 20680 45558
rect 20260 42764 20312 42770
rect 20260 42706 20312 42712
rect 20352 42560 20404 42566
rect 20352 42502 20404 42508
rect 20168 42016 20220 42022
rect 20168 41958 20220 41964
rect 20180 38894 20208 41958
rect 20260 39840 20312 39846
rect 20258 39808 20260 39817
rect 20312 39808 20314 39817
rect 20258 39743 20314 39752
rect 20272 39642 20300 39743
rect 20260 39636 20312 39642
rect 20260 39578 20312 39584
rect 20260 39500 20312 39506
rect 20260 39442 20312 39448
rect 20168 38888 20220 38894
rect 20168 38830 20220 38836
rect 20076 38412 20128 38418
rect 20128 38372 20208 38400
rect 20076 38354 20128 38360
rect 20076 38276 20128 38282
rect 20076 38218 20128 38224
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 19812 33918 19932 33946
rect 19616 33652 19668 33658
rect 19616 33594 19668 33600
rect 19708 33652 19760 33658
rect 19708 33594 19760 33600
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19524 32496 19576 32502
rect 19524 32438 19576 32444
rect 19340 32360 19392 32366
rect 19392 32320 19472 32348
rect 19340 32302 19392 32308
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19248 31748 19300 31754
rect 19248 31690 19300 31696
rect 19248 30184 19300 30190
rect 19248 30126 19300 30132
rect 19260 28422 19288 30126
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 19260 27878 19288 28018
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19352 27334 19380 32166
rect 19444 31890 19472 32320
rect 19628 32026 19656 32914
rect 19812 32774 19840 33918
rect 19892 33856 19944 33862
rect 19892 33798 19944 33804
rect 19904 33046 19932 33798
rect 19892 33040 19944 33046
rect 19892 32982 19944 32988
rect 19800 32768 19852 32774
rect 19800 32710 19852 32716
rect 19800 32428 19852 32434
rect 19800 32370 19852 32376
rect 19812 32298 19840 32370
rect 19800 32292 19852 32298
rect 19800 32234 19852 32240
rect 19812 32026 19840 32234
rect 19616 32020 19668 32026
rect 19616 31962 19668 31968
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19524 31952 19576 31958
rect 19524 31894 19576 31900
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19536 31754 19564 31894
rect 19444 31726 19564 31754
rect 19444 30190 19472 31726
rect 19628 31226 19656 31962
rect 19536 31198 19656 31226
rect 19536 30598 19564 31198
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 19524 30592 19576 30598
rect 19524 30534 19576 30540
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19432 29708 19484 29714
rect 19432 29650 19484 29656
rect 19444 29102 19472 29650
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19444 28422 19472 29038
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19444 27146 19472 28358
rect 19352 27118 19472 27146
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19260 26382 19288 26794
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 19064 23044 19116 23050
rect 19064 22986 19116 22992
rect 19076 22642 19104 22986
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18984 22494 19104 22522
rect 18892 22066 19012 22094
rect 18708 21270 18828 21298
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18524 20534 18552 21082
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18340 18358 18368 19858
rect 18616 19417 18644 20266
rect 18602 19408 18658 19417
rect 18602 19343 18658 19352
rect 18708 19174 18736 21270
rect 18786 21176 18842 21185
rect 18786 21111 18842 21120
rect 18800 21010 18828 21111
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18800 20466 18828 20946
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18694 18864 18750 18873
rect 18694 18799 18750 18808
rect 18708 18766 18736 18799
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17972 17882 18000 18158
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18340 17678 18368 18294
rect 18418 18048 18474 18057
rect 18418 17983 18474 17992
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17270 17908 17478
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17880 16658 17908 17206
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17788 16510 17908 16538
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17788 13530 17816 14350
rect 17880 14006 17908 16510
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18340 15502 18368 17614
rect 18432 17338 18460 17983
rect 18800 17814 18828 19654
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18340 15026 18368 15438
rect 18432 15162 18460 15982
rect 18524 15706 18552 16526
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18524 15094 18552 15642
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18340 14482 18368 14962
rect 18616 14958 18644 16934
rect 18708 16794 18736 17206
rect 18800 17066 18828 17750
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18708 15502 18736 15846
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18708 14890 18736 15302
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18708 14550 18736 14826
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 18800 13938 18828 15506
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 12782 17816 13466
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18064 12306 18092 12650
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17788 2514 17816 8774
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17880 800 17908 3538
rect 18340 3534 18368 13806
rect 18800 12986 18828 13874
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18892 12434 18920 19926
rect 18984 19514 19012 22066
rect 19076 21894 19104 22494
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 19076 19530 19104 21830
rect 19168 19854 19196 24618
rect 19260 22166 19288 26318
rect 19352 25838 19380 27118
rect 19536 27010 19564 30534
rect 19444 26982 19564 27010
rect 19444 26926 19472 26982
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19524 26920 19576 26926
rect 19524 26862 19576 26868
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19444 25906 19472 26726
rect 19536 26042 19564 26862
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19352 24206 19380 24550
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 19352 23730 19380 24142
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19352 22710 19380 23666
rect 19444 22778 19472 25638
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19248 22160 19300 22166
rect 19248 22102 19300 22108
rect 19444 22030 19472 22170
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21690 19472 21830
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 18972 19508 19024 19514
rect 19076 19502 19196 19530
rect 18972 19450 19024 19456
rect 19064 19440 19116 19446
rect 19064 19382 19116 19388
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18984 15042 19012 17274
rect 19076 15162 19104 19382
rect 19168 17082 19196 19502
rect 19260 17202 19288 21286
rect 19536 21162 19564 25638
rect 19628 23746 19656 31078
rect 19798 30696 19854 30705
rect 19708 30660 19760 30666
rect 19798 30631 19800 30640
rect 19708 30602 19760 30608
rect 19852 30631 19854 30640
rect 19800 30602 19852 30608
rect 19720 30326 19748 30602
rect 19708 30320 19760 30326
rect 19708 30262 19760 30268
rect 19892 30252 19944 30258
rect 19892 30194 19944 30200
rect 19800 30116 19852 30122
rect 19800 30058 19852 30064
rect 19812 29714 19840 30058
rect 19800 29708 19852 29714
rect 19800 29650 19852 29656
rect 19800 29572 19852 29578
rect 19800 29514 19852 29520
rect 19812 29170 19840 29514
rect 19800 29164 19852 29170
rect 19800 29106 19852 29112
rect 19904 29034 19932 30194
rect 19996 30054 20024 36722
rect 20088 32858 20116 38218
rect 20180 36922 20208 38372
rect 20168 36916 20220 36922
rect 20168 36858 20220 36864
rect 20272 35154 20300 39442
rect 20364 39098 20392 42502
rect 20456 40526 20484 45526
rect 20628 45494 20680 45500
rect 20720 45552 20772 45558
rect 20720 45494 20772 45500
rect 20640 44810 20668 45494
rect 21192 45422 21220 46446
rect 21180 45416 21232 45422
rect 21180 45358 21232 45364
rect 21192 44878 21220 45358
rect 21180 44872 21232 44878
rect 21180 44814 21232 44820
rect 20628 44804 20680 44810
rect 20628 44746 20680 44752
rect 20640 43722 20668 44746
rect 21284 44742 21312 53382
rect 21548 50176 21600 50182
rect 21548 50118 21600 50124
rect 21560 47818 21588 50118
rect 21652 49722 21680 53926
rect 21744 53582 21772 56200
rect 22112 53582 22140 56200
rect 22480 54194 22508 56200
rect 22468 54188 22520 54194
rect 22468 54130 22520 54136
rect 22192 53984 22244 53990
rect 22284 53984 22336 53990
rect 22192 53926 22244 53932
rect 22282 53952 22284 53961
rect 22336 53952 22338 53961
rect 21732 53576 21784 53582
rect 21732 53518 21784 53524
rect 22100 53576 22152 53582
rect 22100 53518 22152 53524
rect 21744 53242 21772 53518
rect 21916 53440 21968 53446
rect 21916 53382 21968 53388
rect 21732 53236 21784 53242
rect 21732 53178 21784 53184
rect 21652 49694 21772 49722
rect 21560 47790 21680 47818
rect 21548 47116 21600 47122
rect 21548 47058 21600 47064
rect 21560 44810 21588 47058
rect 21364 44804 21416 44810
rect 21364 44746 21416 44752
rect 21548 44804 21600 44810
rect 21548 44746 21600 44752
rect 21272 44736 21324 44742
rect 21272 44678 21324 44684
rect 21376 44538 21404 44746
rect 21364 44532 21416 44538
rect 21364 44474 21416 44480
rect 21088 43852 21140 43858
rect 21088 43794 21140 43800
rect 20628 43716 20680 43722
rect 20628 43658 20680 43664
rect 20640 43110 20668 43658
rect 20628 43104 20680 43110
rect 20628 43046 20680 43052
rect 20996 43104 21048 43110
rect 20996 43046 21048 43052
rect 20640 42634 20668 43046
rect 20536 42628 20588 42634
rect 20536 42570 20588 42576
rect 20628 42628 20680 42634
rect 20628 42570 20680 42576
rect 20444 40520 20496 40526
rect 20444 40462 20496 40468
rect 20352 39092 20404 39098
rect 20352 39034 20404 39040
rect 20352 37868 20404 37874
rect 20352 37810 20404 37816
rect 20260 35148 20312 35154
rect 20260 35090 20312 35096
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20272 32978 20300 34546
rect 20364 33454 20392 37810
rect 20548 36854 20576 42570
rect 20640 42294 20668 42570
rect 20628 42288 20680 42294
rect 20628 42230 20680 42236
rect 21008 42158 21036 43046
rect 20996 42152 21048 42158
rect 20996 42094 21048 42100
rect 20904 42016 20956 42022
rect 20904 41958 20956 41964
rect 20720 41608 20772 41614
rect 20720 41550 20772 41556
rect 20812 41608 20864 41614
rect 20812 41550 20864 41556
rect 20732 40594 20760 41550
rect 20824 41274 20852 41550
rect 20916 41546 20944 41958
rect 20904 41540 20956 41546
rect 20904 41482 20956 41488
rect 20996 41472 21048 41478
rect 20996 41414 21048 41420
rect 20812 41268 20864 41274
rect 20812 41210 20864 41216
rect 20720 40588 20772 40594
rect 20720 40530 20772 40536
rect 21008 40372 21036 41414
rect 21100 41070 21128 43794
rect 21272 43648 21324 43654
rect 21272 43590 21324 43596
rect 21284 42770 21312 43590
rect 21364 43308 21416 43314
rect 21364 43250 21416 43256
rect 21376 43110 21404 43250
rect 21364 43104 21416 43110
rect 21362 43072 21364 43081
rect 21456 43104 21508 43110
rect 21416 43072 21418 43081
rect 21456 43046 21508 43052
rect 21362 43007 21418 43016
rect 21272 42764 21324 42770
rect 21272 42706 21324 42712
rect 21284 42362 21312 42706
rect 21468 42702 21496 43046
rect 21560 42838 21588 44746
rect 21548 42832 21600 42838
rect 21548 42774 21600 42780
rect 21456 42696 21508 42702
rect 21456 42638 21508 42644
rect 21272 42356 21324 42362
rect 21272 42298 21324 42304
rect 21272 41540 21324 41546
rect 21272 41482 21324 41488
rect 21180 41200 21232 41206
rect 21178 41168 21180 41177
rect 21232 41168 21234 41177
rect 21178 41103 21234 41112
rect 21088 41064 21140 41070
rect 21088 41006 21140 41012
rect 21100 40934 21128 41006
rect 21088 40928 21140 40934
rect 21088 40870 21140 40876
rect 21180 40520 21232 40526
rect 21180 40462 21232 40468
rect 21088 40384 21140 40390
rect 21008 40344 21088 40372
rect 21088 40326 21140 40332
rect 20996 40112 21048 40118
rect 20996 40054 21048 40060
rect 20904 39296 20956 39302
rect 20904 39238 20956 39244
rect 20720 38888 20772 38894
rect 20720 38830 20772 38836
rect 20732 38758 20760 38830
rect 20720 38752 20772 38758
rect 20720 38694 20772 38700
rect 20812 38752 20864 38758
rect 20812 38694 20864 38700
rect 20628 38208 20680 38214
rect 20628 38150 20680 38156
rect 20640 38010 20668 38150
rect 20628 38004 20680 38010
rect 20628 37946 20680 37952
rect 20640 37369 20668 37946
rect 20626 37360 20682 37369
rect 20626 37295 20682 37304
rect 20628 37120 20680 37126
rect 20628 37062 20680 37068
rect 20536 36848 20588 36854
rect 20536 36790 20588 36796
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20352 33448 20404 33454
rect 20352 33390 20404 33396
rect 20260 32972 20312 32978
rect 20260 32914 20312 32920
rect 20456 32858 20484 36654
rect 20088 32830 20300 32858
rect 20364 32842 20484 32858
rect 20076 30796 20128 30802
rect 20076 30738 20128 30744
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19892 29028 19944 29034
rect 19892 28970 19944 28976
rect 19706 28248 19762 28257
rect 19904 28218 19932 28970
rect 19706 28183 19708 28192
rect 19760 28183 19762 28192
rect 19892 28212 19944 28218
rect 19708 28154 19760 28160
rect 19892 28154 19944 28160
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 19720 27878 19748 27950
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 19800 27668 19852 27674
rect 19800 27610 19852 27616
rect 19812 27470 19840 27610
rect 19800 27464 19852 27470
rect 19800 27406 19852 27412
rect 19708 27328 19760 27334
rect 19706 27296 19708 27305
rect 19760 27296 19762 27305
rect 19706 27231 19762 27240
rect 19720 26790 19748 27231
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19708 26512 19760 26518
rect 19708 26454 19760 26460
rect 19720 25702 19748 26454
rect 19708 25696 19760 25702
rect 19708 25638 19760 25644
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19708 25152 19760 25158
rect 19760 25112 19840 25140
rect 19708 25094 19760 25100
rect 19628 23718 19748 23746
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19628 23322 19656 23598
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19720 22094 19748 23718
rect 19812 23610 19840 25112
rect 19904 24954 19932 25638
rect 19892 24948 19944 24954
rect 19892 24890 19944 24896
rect 19996 24818 20024 29446
rect 20088 27538 20116 30738
rect 20272 30122 20300 32830
rect 20352 32836 20484 32842
rect 20404 32830 20484 32836
rect 20352 32778 20404 32784
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 20364 31686 20392 32438
rect 20352 31680 20404 31686
rect 20352 31622 20404 31628
rect 20456 30258 20484 32830
rect 20640 32570 20668 37062
rect 20824 34610 20852 38694
rect 20916 36242 20944 39238
rect 21008 39030 21036 40054
rect 20996 39024 21048 39030
rect 20996 38966 21048 38972
rect 20996 38752 21048 38758
rect 20996 38694 21048 38700
rect 21008 36650 21036 38694
rect 20996 36644 21048 36650
rect 20996 36586 21048 36592
rect 20904 36236 20956 36242
rect 20904 36178 20956 36184
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20720 34536 20772 34542
rect 20720 34478 20772 34484
rect 20732 33862 20760 34478
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20812 33856 20864 33862
rect 20812 33798 20864 33804
rect 20720 33312 20772 33318
rect 20720 33254 20772 33260
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20536 32360 20588 32366
rect 20536 32302 20588 32308
rect 20548 31958 20576 32302
rect 20640 32026 20668 32506
rect 20628 32020 20680 32026
rect 20628 31962 20680 31968
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 20732 31482 20760 33254
rect 20720 31476 20772 31482
rect 20720 31418 20772 31424
rect 20720 31136 20772 31142
rect 20720 31078 20772 31084
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 20260 30116 20312 30122
rect 20260 30058 20312 30064
rect 20536 30116 20588 30122
rect 20536 30058 20588 30064
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20260 27600 20312 27606
rect 20260 27542 20312 27548
rect 20076 27532 20128 27538
rect 20076 27474 20128 27480
rect 20088 26926 20116 27474
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 20180 25294 20208 27270
rect 20168 25288 20220 25294
rect 20168 25230 20220 25236
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19812 23582 20024 23610
rect 19720 22066 19840 22094
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19444 21134 19564 21162
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20398 19380 20742
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19444 18970 19472 21134
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19536 20602 19564 21014
rect 19720 20874 19748 21626
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19444 18630 19472 18906
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19168 17054 19288 17082
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19168 15502 19196 15982
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19260 15314 19288 17054
rect 19352 16538 19380 18362
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 17542 19472 18226
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19352 16510 19472 16538
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19352 15434 19380 16390
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19168 15286 19288 15314
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 18984 15014 19104 15042
rect 18892 12406 19012 12434
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11830 18920 12174
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18984 10062 19012 12406
rect 19076 11354 19104 15014
rect 19168 13258 19196 15286
rect 19444 15042 19472 16510
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19352 15014 19472 15042
rect 19352 13802 19380 15014
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19444 14074 19472 14894
rect 19536 14074 19564 15302
rect 19628 14414 19656 20198
rect 19812 19922 19840 22066
rect 19996 20534 20024 23582
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 20088 21554 20116 22646
rect 20272 21622 20300 27542
rect 20352 27056 20404 27062
rect 20352 26998 20404 27004
rect 20364 26586 20392 26998
rect 20456 26994 20484 29990
rect 20548 29306 20576 30058
rect 20536 29300 20588 29306
rect 20536 29242 20588 29248
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20548 28626 20576 28902
rect 20536 28620 20588 28626
rect 20536 28562 20588 28568
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20364 24750 20392 26522
rect 20444 25968 20496 25974
rect 20444 25910 20496 25916
rect 20456 25158 20484 25910
rect 20444 25152 20496 25158
rect 20444 25094 20496 25100
rect 20352 24744 20404 24750
rect 20352 24686 20404 24692
rect 20548 24274 20576 27338
rect 20640 26586 20668 27814
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20732 25226 20760 31078
rect 20824 29646 20852 33798
rect 20916 31414 20944 35974
rect 21008 35086 21036 36586
rect 21100 36174 21128 40326
rect 21192 39438 21220 40462
rect 21180 39432 21232 39438
rect 21180 39374 21232 39380
rect 21284 38010 21312 41482
rect 21468 41414 21496 42638
rect 21548 41540 21600 41546
rect 21548 41482 21600 41488
rect 21376 41386 21496 41414
rect 21376 40186 21404 41386
rect 21456 40928 21508 40934
rect 21456 40870 21508 40876
rect 21364 40180 21416 40186
rect 21364 40122 21416 40128
rect 21468 39817 21496 40870
rect 21454 39808 21510 39817
rect 21454 39743 21510 39752
rect 21560 38826 21588 41482
rect 21652 40526 21680 47790
rect 21744 43314 21772 49694
rect 21928 46986 21956 53382
rect 22112 53242 22140 53518
rect 22100 53236 22152 53242
rect 22100 53178 22152 53184
rect 21916 46980 21968 46986
rect 21916 46922 21968 46928
rect 22204 46646 22232 53926
rect 22282 53887 22338 53896
rect 22284 53712 22336 53718
rect 22284 53654 22336 53660
rect 22192 46640 22244 46646
rect 22192 46582 22244 46588
rect 21916 46028 21968 46034
rect 21916 45970 21968 45976
rect 21928 45286 21956 45970
rect 21916 45280 21968 45286
rect 21916 45222 21968 45228
rect 21824 44736 21876 44742
rect 21822 44704 21824 44713
rect 21876 44704 21878 44713
rect 21822 44639 21878 44648
rect 21836 44538 21864 44639
rect 21824 44532 21876 44538
rect 21824 44474 21876 44480
rect 21928 44470 21956 45222
rect 22008 44872 22060 44878
rect 22008 44814 22060 44820
rect 21916 44464 21968 44470
rect 21916 44406 21968 44412
rect 21732 43308 21784 43314
rect 21732 43250 21784 43256
rect 21732 42832 21784 42838
rect 21732 42774 21784 42780
rect 21744 40662 21772 42774
rect 21824 42220 21876 42226
rect 21824 42162 21876 42168
rect 21732 40656 21784 40662
rect 21732 40598 21784 40604
rect 21640 40520 21692 40526
rect 21640 40462 21692 40468
rect 21732 40452 21784 40458
rect 21732 40394 21784 40400
rect 21640 39976 21692 39982
rect 21640 39918 21692 39924
rect 21652 39438 21680 39918
rect 21640 39432 21692 39438
rect 21640 39374 21692 39380
rect 21548 38820 21600 38826
rect 21548 38762 21600 38768
rect 21548 38480 21600 38486
rect 21548 38422 21600 38428
rect 21364 38344 21416 38350
rect 21364 38286 21416 38292
rect 21272 38004 21324 38010
rect 21272 37946 21324 37952
rect 21284 37466 21312 37946
rect 21272 37460 21324 37466
rect 21272 37402 21324 37408
rect 21284 37262 21312 37402
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 21376 36922 21404 38286
rect 21560 37806 21588 38422
rect 21548 37800 21600 37806
rect 21652 37788 21680 39374
rect 21744 37942 21772 40394
rect 21836 39137 21864 42162
rect 21928 41070 21956 44406
rect 22020 43722 22048 44814
rect 22100 44192 22152 44198
rect 22100 44134 22152 44140
rect 22008 43716 22060 43722
rect 22008 43658 22060 43664
rect 22020 42770 22048 43658
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 22020 41682 22048 42706
rect 22008 41676 22060 41682
rect 22008 41618 22060 41624
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 21916 41064 21968 41070
rect 21916 41006 21968 41012
rect 22020 41002 22048 41210
rect 22008 40996 22060 41002
rect 22008 40938 22060 40944
rect 22008 40656 22060 40662
rect 22008 40598 22060 40604
rect 21916 40588 21968 40594
rect 21916 40530 21968 40536
rect 21928 40118 21956 40530
rect 21916 40112 21968 40118
rect 21916 40054 21968 40060
rect 22020 39982 22048 40598
rect 22008 39976 22060 39982
rect 22008 39918 22060 39924
rect 21914 39808 21970 39817
rect 21914 39743 21970 39752
rect 21822 39128 21878 39137
rect 21822 39063 21878 39072
rect 21824 38888 21876 38894
rect 21824 38830 21876 38836
rect 21732 37936 21784 37942
rect 21732 37878 21784 37884
rect 21652 37760 21772 37788
rect 21548 37742 21600 37748
rect 21548 37664 21600 37670
rect 21548 37606 21600 37612
rect 21364 36916 21416 36922
rect 21364 36858 21416 36864
rect 21376 36650 21404 36858
rect 21364 36644 21416 36650
rect 21364 36586 21416 36592
rect 21180 36304 21232 36310
rect 21180 36246 21232 36252
rect 21088 36168 21140 36174
rect 21088 36110 21140 36116
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 21088 35012 21140 35018
rect 21088 34954 21140 34960
rect 21100 34202 21128 34954
rect 21192 34950 21220 36246
rect 21180 34944 21232 34950
rect 21180 34886 21232 34892
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 20996 33992 21048 33998
rect 20996 33934 21048 33940
rect 21008 31482 21036 33934
rect 21192 33522 21220 34886
rect 21364 34196 21416 34202
rect 21364 34138 21416 34144
rect 21376 34066 21404 34138
rect 21364 34060 21416 34066
rect 21364 34002 21416 34008
rect 21456 34060 21508 34066
rect 21456 34002 21508 34008
rect 21180 33516 21232 33522
rect 21180 33458 21232 33464
rect 21088 32972 21140 32978
rect 21088 32914 21140 32920
rect 21100 31890 21128 32914
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 21180 31884 21232 31890
rect 21180 31826 21232 31832
rect 21192 31754 21220 31826
rect 21100 31726 21220 31754
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 20904 31408 20956 31414
rect 20904 31350 20956 31356
rect 21100 30682 21128 31726
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21178 31512 21234 31521
rect 21178 31447 21180 31456
rect 21232 31447 21234 31456
rect 21180 31418 21232 31424
rect 21192 30938 21220 31418
rect 21272 31272 21324 31278
rect 21272 31214 21324 31220
rect 21180 30932 21232 30938
rect 21180 30874 21232 30880
rect 21100 30654 21220 30682
rect 21088 30592 21140 30598
rect 21088 30534 21140 30540
rect 20904 30184 20956 30190
rect 20904 30126 20956 30132
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20916 29238 20944 30126
rect 20996 29776 21048 29782
rect 20996 29718 21048 29724
rect 20904 29232 20956 29238
rect 20904 29174 20956 29180
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20916 27130 20944 27270
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20824 26518 20852 26862
rect 20812 26512 20864 26518
rect 20812 26454 20864 26460
rect 20904 25764 20956 25770
rect 20904 25706 20956 25712
rect 20916 25226 20944 25706
rect 20720 25220 20772 25226
rect 20720 25162 20772 25168
rect 20904 25220 20956 25226
rect 20904 25162 20956 25168
rect 21008 24818 21036 29718
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20548 23644 20576 24210
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 20628 23656 20680 23662
rect 20548 23616 20628 23644
rect 20628 23598 20680 23604
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20364 22710 20392 22918
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20364 22234 20392 22646
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 20180 19446 20208 20810
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 20364 18970 20392 22170
rect 20548 21554 20576 22714
rect 20628 22500 20680 22506
rect 20628 22442 20680 22448
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19720 17542 19748 18770
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19812 18086 19840 18702
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17270 19748 17478
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19812 16046 19840 18022
rect 19904 16250 19932 18838
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18426 20024 18566
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 16250 20024 16390
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 20088 15586 20116 18634
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20180 16250 20208 18566
rect 20364 18358 20392 18906
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20456 17524 20484 19110
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20548 17592 20576 18226
rect 20640 18154 20668 22442
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 20890 20760 21898
rect 20824 21010 20852 23054
rect 20916 21894 20944 23734
rect 21008 22642 21036 23802
rect 21100 23798 21128 30534
rect 21192 28150 21220 30654
rect 21180 28144 21232 28150
rect 21180 28086 21232 28092
rect 21180 28008 21232 28014
rect 21180 27950 21232 27956
rect 21192 24818 21220 27950
rect 21284 27402 21312 31214
rect 21376 30598 21404 31622
rect 21364 30592 21416 30598
rect 21364 30534 21416 30540
rect 21376 28082 21404 30534
rect 21468 29510 21496 34002
rect 21560 32502 21588 37606
rect 21640 36916 21692 36922
rect 21640 36858 21692 36864
rect 21548 32496 21600 32502
rect 21548 32438 21600 32444
rect 21548 32360 21600 32366
rect 21548 32302 21600 32308
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21560 28608 21588 32302
rect 21652 31686 21680 36858
rect 21744 33930 21772 37760
rect 21836 34678 21864 38830
rect 21824 34672 21876 34678
rect 21824 34614 21876 34620
rect 21836 33998 21864 34614
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21732 33924 21784 33930
rect 21732 33866 21784 33872
rect 21824 33380 21876 33386
rect 21824 33322 21876 33328
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21640 31680 21692 31686
rect 21640 31622 21692 31628
rect 21640 29504 21692 29510
rect 21640 29446 21692 29452
rect 21652 29306 21680 29446
rect 21640 29300 21692 29306
rect 21640 29242 21692 29248
rect 21468 28580 21588 28608
rect 21364 28076 21416 28082
rect 21364 28018 21416 28024
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 21272 27396 21324 27402
rect 21272 27338 21324 27344
rect 21376 27130 21404 27406
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 21468 26926 21496 28580
rect 21548 28484 21600 28490
rect 21548 28426 21600 28432
rect 21456 26920 21508 26926
rect 21456 26862 21508 26868
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21088 23792 21140 23798
rect 21088 23734 21140 23740
rect 21284 23730 21312 25298
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21088 23248 21140 23254
rect 21088 23190 21140 23196
rect 21100 22642 21128 23190
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21690 20944 21830
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20732 20862 20852 20890
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20628 17604 20680 17610
rect 20548 17564 20628 17592
rect 20628 17546 20680 17552
rect 20456 17496 20576 17524
rect 20260 17060 20312 17066
rect 20260 17002 20312 17008
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 19996 15558 20116 15586
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 19812 14958 19840 15030
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19536 12918 19564 13670
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19444 11354 19472 11630
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19076 11150 19104 11290
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19536 10810 19564 12038
rect 19720 11898 19748 14214
rect 19812 13734 19840 14894
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18800 4049 18828 4082
rect 18786 4040 18842 4049
rect 18786 3975 18842 3984
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18340 1170 18368 2926
rect 18524 2650 18552 2994
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18248 1142 18368 1170
rect 18248 800 18276 1142
rect 18616 800 18644 3062
rect 18984 800 19012 3402
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19352 800 19380 3130
rect 19444 2446 19472 9318
rect 19628 4622 19656 11018
rect 19720 6390 19748 11834
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19904 11558 19932 11698
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19904 10674 19932 11494
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 9586 19932 10406
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19996 5574 20024 15558
rect 20272 12434 20300 17002
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20364 12889 20392 13194
rect 20350 12880 20406 12889
rect 20350 12815 20406 12824
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20272 12406 20392 12434
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 20088 11150 20116 12310
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20364 8974 20392 12406
rect 20456 10674 20484 12582
rect 20548 11830 20576 17496
rect 20640 16794 20668 17546
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20732 15162 20760 17138
rect 20824 16590 20852 20862
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20824 16114 20852 16390
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20824 15570 20852 16050
rect 20916 15706 20944 18362
rect 21008 16590 21036 19994
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21100 18834 21128 19246
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21100 18222 21128 18770
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 21100 17746 21128 18158
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 17134 21128 17682
rect 21192 17610 21220 18566
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21284 17134 21312 20266
rect 21468 19700 21496 24550
rect 21560 23866 21588 28426
rect 21744 26994 21772 32846
rect 21836 32842 21864 33322
rect 21824 32836 21876 32842
rect 21824 32778 21876 32784
rect 21928 32366 21956 39743
rect 22008 38752 22060 38758
rect 22008 38694 22060 38700
rect 22020 38350 22048 38694
rect 22112 38418 22140 44134
rect 22192 43784 22244 43790
rect 22192 43726 22244 43732
rect 22204 42566 22232 43726
rect 22296 43450 22324 53654
rect 22480 53242 22508 54130
rect 22848 53582 22876 56200
rect 23216 55214 23244 56200
rect 23216 55186 23336 55214
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 22836 53576 22888 53582
rect 22836 53518 22888 53524
rect 23308 53242 23336 55186
rect 22468 53236 22520 53242
rect 22468 53178 22520 53184
rect 23296 53236 23348 53242
rect 23296 53178 23348 53184
rect 23584 53106 23612 56200
rect 24490 56199 24546 56208
rect 24504 54330 24532 56199
rect 24674 55448 24730 55457
rect 24674 55383 24730 55392
rect 24688 54330 24716 55383
rect 24766 54632 24822 54641
rect 24766 54567 24822 54576
rect 24492 54324 24544 54330
rect 24492 54266 24544 54272
rect 24676 54324 24728 54330
rect 24676 54266 24728 54272
rect 24504 53582 24532 54266
rect 24584 53984 24636 53990
rect 24584 53926 24636 53932
rect 24492 53576 24544 53582
rect 24492 53518 24544 53524
rect 23848 53440 23900 53446
rect 23848 53382 23900 53388
rect 23572 53100 23624 53106
rect 23572 53042 23624 53048
rect 23296 52896 23348 52902
rect 23296 52838 23348 52844
rect 23388 52896 23440 52902
rect 23388 52838 23440 52844
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22468 47184 22520 47190
rect 22468 47126 22520 47132
rect 22376 46028 22428 46034
rect 22376 45970 22428 45976
rect 22388 45830 22416 45970
rect 22376 45824 22428 45830
rect 22376 45766 22428 45772
rect 22388 43450 22416 45766
rect 22480 43654 22508 47126
rect 22744 46572 22796 46578
rect 22744 46514 22796 46520
rect 22560 46504 22612 46510
rect 22560 46446 22612 46452
rect 22468 43648 22520 43654
rect 22468 43590 22520 43596
rect 22284 43444 22336 43450
rect 22284 43386 22336 43392
rect 22376 43444 22428 43450
rect 22376 43386 22428 43392
rect 22572 43330 22600 46446
rect 22756 46322 22784 46514
rect 22664 46294 22784 46322
rect 22664 43994 22692 46294
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22744 44736 22796 44742
rect 22744 44678 22796 44684
rect 22652 43988 22704 43994
rect 22652 43930 22704 43936
rect 22756 43858 22784 44678
rect 23308 44538 23336 52838
rect 23400 46714 23428 52838
rect 23860 52601 23888 53382
rect 23846 52592 23902 52601
rect 23846 52527 23902 52536
rect 24124 47116 24176 47122
rect 24124 47058 24176 47064
rect 23388 46708 23440 46714
rect 23388 46650 23440 46656
rect 23664 46504 23716 46510
rect 23664 46446 23716 46452
rect 23676 45898 23704 46446
rect 24032 45960 24084 45966
rect 24032 45902 24084 45908
rect 23664 45892 23716 45898
rect 23664 45834 23716 45840
rect 23480 45824 23532 45830
rect 23480 45766 23532 45772
rect 23492 45558 23520 45766
rect 23388 45552 23440 45558
rect 23388 45494 23440 45500
rect 23480 45552 23532 45558
rect 23480 45494 23532 45500
rect 23296 44532 23348 44538
rect 23296 44474 23348 44480
rect 22836 44192 22888 44198
rect 22836 44134 22888 44140
rect 22848 43926 22876 44134
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22836 43920 22888 43926
rect 22836 43862 22888 43868
rect 22744 43852 22796 43858
rect 22744 43794 22796 43800
rect 22652 43648 22704 43654
rect 22652 43590 22704 43596
rect 22296 43302 22600 43330
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 22190 41576 22246 41585
rect 22190 41511 22246 41520
rect 22204 40526 22232 41511
rect 22192 40520 22244 40526
rect 22192 40462 22244 40468
rect 22204 40050 22232 40462
rect 22192 40044 22244 40050
rect 22192 39986 22244 39992
rect 22192 39908 22244 39914
rect 22296 39896 22324 43302
rect 22468 43240 22520 43246
rect 22468 43182 22520 43188
rect 22376 43172 22428 43178
rect 22376 43114 22428 43120
rect 22244 39868 22324 39896
rect 22192 39850 22244 39856
rect 22296 39574 22324 39868
rect 22284 39568 22336 39574
rect 22284 39510 22336 39516
rect 22192 39296 22244 39302
rect 22192 39238 22244 39244
rect 22284 39296 22336 39302
rect 22284 39238 22336 39244
rect 22204 38962 22232 39238
rect 22192 38956 22244 38962
rect 22192 38898 22244 38904
rect 22100 38412 22152 38418
rect 22100 38354 22152 38360
rect 22008 38344 22060 38350
rect 22204 38321 22232 38898
rect 22008 38286 22060 38292
rect 22190 38312 22246 38321
rect 22100 38276 22152 38282
rect 22296 38282 22324 39238
rect 22388 38298 22416 43114
rect 22480 41478 22508 43182
rect 22560 42356 22612 42362
rect 22560 42298 22612 42304
rect 22572 42226 22600 42298
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 22560 42016 22612 42022
rect 22560 41958 22612 41964
rect 22572 41818 22600 41958
rect 22560 41812 22612 41818
rect 22560 41754 22612 41760
rect 22468 41472 22520 41478
rect 22468 41414 22520 41420
rect 22466 41168 22522 41177
rect 22466 41103 22468 41112
rect 22520 41103 22522 41112
rect 22468 41074 22520 41080
rect 22468 40928 22520 40934
rect 22468 40870 22520 40876
rect 22480 40730 22508 40870
rect 22468 40724 22520 40730
rect 22468 40666 22520 40672
rect 22480 40474 22508 40666
rect 22572 40594 22600 41754
rect 22664 41274 22692 43590
rect 22756 41682 22784 43794
rect 23400 43450 23428 45494
rect 23676 45370 23704 45834
rect 24044 45490 24072 45902
rect 24032 45484 24084 45490
rect 24032 45426 24084 45432
rect 23492 45342 23704 45370
rect 23492 44810 23520 45342
rect 24044 44946 24072 45426
rect 24032 44940 24084 44946
rect 24032 44882 24084 44888
rect 23480 44804 23532 44810
rect 23480 44746 23532 44752
rect 23492 43994 23520 44746
rect 23572 44328 23624 44334
rect 23572 44270 23624 44276
rect 23480 43988 23532 43994
rect 23480 43930 23532 43936
rect 23480 43648 23532 43654
rect 23480 43590 23532 43596
rect 23388 43444 23440 43450
rect 23388 43386 23440 43392
rect 23388 43172 23440 43178
rect 23388 43114 23440 43120
rect 23296 43104 23348 43110
rect 23296 43046 23348 43052
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 23308 42378 23336 43046
rect 23216 42350 23336 42378
rect 22836 42152 22888 42158
rect 22836 42094 22888 42100
rect 22744 41676 22796 41682
rect 22744 41618 22796 41624
rect 22848 41614 22876 42094
rect 23216 42022 23244 42350
rect 23204 42016 23256 42022
rect 23204 41958 23256 41964
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22836 41608 22888 41614
rect 22836 41550 22888 41556
rect 22744 41472 22796 41478
rect 22744 41414 22796 41420
rect 22836 41472 22888 41478
rect 22836 41414 22888 41420
rect 22652 41268 22704 41274
rect 22652 41210 22704 41216
rect 22756 41070 22784 41414
rect 22848 41274 22876 41414
rect 22836 41268 22888 41274
rect 22836 41210 22888 41216
rect 22834 41168 22890 41177
rect 22834 41103 22890 41112
rect 22744 41064 22796 41070
rect 22744 41006 22796 41012
rect 22560 40588 22612 40594
rect 22560 40530 22612 40536
rect 22480 40446 22600 40474
rect 22468 40384 22520 40390
rect 22468 40326 22520 40332
rect 22480 40089 22508 40326
rect 22466 40080 22522 40089
rect 22466 40015 22522 40024
rect 22572 39930 22600 40446
rect 22480 39902 22600 39930
rect 22480 39030 22508 39902
rect 22560 39840 22612 39846
rect 22558 39808 22560 39817
rect 22612 39808 22614 39817
rect 22558 39743 22614 39752
rect 22468 39024 22520 39030
rect 22468 38966 22520 38972
rect 22480 38758 22508 38966
rect 22572 38894 22600 39743
rect 22652 39568 22704 39574
rect 22652 39510 22704 39516
rect 22560 38888 22612 38894
rect 22560 38830 22612 38836
rect 22468 38752 22520 38758
rect 22466 38720 22468 38729
rect 22520 38720 22522 38729
rect 22466 38655 22522 38664
rect 22664 38486 22692 39510
rect 22652 38480 22704 38486
rect 22652 38422 22704 38428
rect 22190 38247 22246 38256
rect 22284 38276 22336 38282
rect 22100 38218 22152 38224
rect 22388 38270 22508 38298
rect 22284 38218 22336 38224
rect 22112 37262 22140 38218
rect 22376 38208 22428 38214
rect 22376 38150 22428 38156
rect 22190 38040 22246 38049
rect 22190 37975 22192 37984
rect 22244 37975 22246 37984
rect 22192 37946 22244 37952
rect 22388 37874 22416 38150
rect 22376 37868 22428 37874
rect 22376 37810 22428 37816
rect 22284 37800 22336 37806
rect 22284 37742 22336 37748
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 22020 33998 22048 35430
rect 22112 34474 22140 37198
rect 22296 37194 22324 37742
rect 22284 37188 22336 37194
rect 22284 37130 22336 37136
rect 22190 36952 22246 36961
rect 22190 36887 22192 36896
rect 22244 36887 22246 36896
rect 22192 36858 22244 36864
rect 22190 36680 22246 36689
rect 22190 36615 22192 36624
rect 22244 36615 22246 36624
rect 22192 36586 22244 36592
rect 22296 36242 22324 37130
rect 22284 36236 22336 36242
rect 22284 36178 22336 36184
rect 22282 36136 22338 36145
rect 22282 36071 22338 36080
rect 22192 35148 22244 35154
rect 22192 35090 22244 35096
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 22020 32978 22048 33934
rect 22100 33040 22152 33046
rect 22100 32982 22152 32988
rect 22008 32972 22060 32978
rect 22008 32914 22060 32920
rect 21916 32360 21968 32366
rect 21916 32302 21968 32308
rect 21914 32056 21970 32065
rect 21914 31991 21970 32000
rect 21928 31958 21956 31991
rect 21916 31952 21968 31958
rect 21916 31894 21968 31900
rect 22112 31686 22140 32982
rect 22204 32570 22232 35090
rect 22296 33318 22324 36071
rect 22388 35873 22416 37810
rect 22480 37738 22508 38270
rect 22560 38208 22612 38214
rect 22560 38150 22612 38156
rect 22468 37732 22520 37738
rect 22468 37674 22520 37680
rect 22480 36854 22508 37674
rect 22468 36848 22520 36854
rect 22468 36790 22520 36796
rect 22374 35864 22430 35873
rect 22374 35799 22430 35808
rect 22480 35494 22508 36790
rect 22468 35488 22520 35494
rect 22468 35430 22520 35436
rect 22376 34604 22428 34610
rect 22376 34546 22428 34552
rect 22284 33312 22336 33318
rect 22284 33254 22336 33260
rect 22284 33040 22336 33046
rect 22284 32982 22336 32988
rect 22192 32564 22244 32570
rect 22192 32506 22244 32512
rect 22192 32360 22244 32366
rect 22192 32302 22244 32308
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21916 30048 21968 30054
rect 21916 29990 21968 29996
rect 21824 29844 21876 29850
rect 21824 29786 21876 29792
rect 21836 29578 21864 29786
rect 21824 29572 21876 29578
rect 21824 29514 21876 29520
rect 21928 29510 21956 29990
rect 21916 29504 21968 29510
rect 21916 29446 21968 29452
rect 22112 29186 22140 31214
rect 22204 29714 22232 32302
rect 22192 29708 22244 29714
rect 22192 29650 22244 29656
rect 22020 29158 22140 29186
rect 22020 27946 22048 29158
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22008 27940 22060 27946
rect 22008 27882 22060 27888
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 21744 26450 21772 26930
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 21916 25424 21968 25430
rect 21916 25366 21968 25372
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21652 24342 21680 25230
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 21640 24336 21692 24342
rect 21640 24278 21692 24284
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21652 23202 21680 24278
rect 21560 23174 21680 23202
rect 21744 23186 21772 25094
rect 21732 23180 21784 23186
rect 21560 23118 21588 23174
rect 21732 23122 21784 23128
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21560 20602 21588 21898
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21468 19672 21588 19700
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21468 17338 21496 19178
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 21008 15450 21036 16118
rect 20824 15422 21036 15450
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20548 11150 20576 11766
rect 20640 11286 20668 14758
rect 20732 13802 20760 15098
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20640 7410 20668 11222
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19720 800 19748 5102
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19904 2514 19932 2790
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 20088 800 20116 4422
rect 20272 4146 20300 7142
rect 20364 5710 20392 7142
rect 20732 6914 20760 13262
rect 20824 11218 20852 15422
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 14618 21036 15302
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21100 14414 21128 17070
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21192 15570 21220 16458
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20916 12170 20944 13262
rect 21008 13258 21036 13466
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21008 12850 21036 13194
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21100 12782 21128 14350
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 21008 11898 21036 12650
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21192 11762 21220 14826
rect 21376 14482 21404 15846
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21468 14226 21496 15982
rect 21560 15502 21588 19672
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21652 15026 21680 21286
rect 21928 19854 21956 25366
rect 22020 25362 22048 27882
rect 22204 27334 22232 28494
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 22112 25226 22140 26862
rect 22204 26382 22232 27270
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22204 23662 22232 26318
rect 22296 25974 22324 32982
rect 22388 32910 22416 34546
rect 22480 34134 22508 35430
rect 22572 34746 22600 38150
rect 22742 38040 22798 38049
rect 22742 37975 22798 37984
rect 22652 37120 22704 37126
rect 22652 37062 22704 37068
rect 22664 36106 22692 37062
rect 22756 36145 22784 37975
rect 22742 36136 22798 36145
rect 22652 36100 22704 36106
rect 22742 36071 22798 36080
rect 22652 36042 22704 36048
rect 22848 35986 22876 41103
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23296 40384 23348 40390
rect 23296 40326 23348 40332
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 23308 39098 23336 40326
rect 23296 39092 23348 39098
rect 23296 39034 23348 39040
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 23294 38448 23350 38457
rect 23400 38418 23428 43114
rect 23294 38383 23350 38392
rect 23388 38412 23440 38418
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23308 37398 23336 38383
rect 23388 38354 23440 38360
rect 23388 38208 23440 38214
rect 23388 38150 23440 38156
rect 23296 37392 23348 37398
rect 23296 37334 23348 37340
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23308 35986 23336 37334
rect 23400 36922 23428 38150
rect 23388 36916 23440 36922
rect 23388 36858 23440 36864
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 22756 35958 22876 35986
rect 22940 35958 23336 35986
rect 22756 35894 22784 35958
rect 22940 35894 22968 35958
rect 22756 35866 22876 35894
rect 22940 35866 23336 35894
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22664 35086 22692 35566
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22652 34944 22704 34950
rect 22652 34886 22704 34892
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22664 34746 22692 34886
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22468 34128 22520 34134
rect 22468 34070 22520 34076
rect 22468 33924 22520 33930
rect 22468 33866 22520 33872
rect 22480 33454 22508 33866
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 22468 33448 22520 33454
rect 22468 33390 22520 33396
rect 22560 33312 22612 33318
rect 22560 33254 22612 33260
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22376 32768 22428 32774
rect 22428 32716 22508 32722
rect 22376 32710 22508 32716
rect 22388 32694 22508 32710
rect 22480 32570 22508 32694
rect 22376 32564 22428 32570
rect 22376 32506 22428 32512
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22388 32450 22416 32506
rect 22388 32422 22508 32450
rect 22376 32360 22428 32366
rect 22376 32302 22428 32308
rect 22388 32026 22416 32302
rect 22376 32020 22428 32026
rect 22376 31962 22428 31968
rect 22376 29096 22428 29102
rect 22376 29038 22428 29044
rect 22388 26314 22416 29038
rect 22480 28490 22508 32422
rect 22572 28762 22600 33254
rect 22664 32026 22692 33798
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22560 28756 22612 28762
rect 22560 28698 22612 28704
rect 22468 28484 22520 28490
rect 22468 28426 22520 28432
rect 22480 28234 22508 28426
rect 22480 28206 22600 28234
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22480 27418 22508 28018
rect 22572 27538 22600 28206
rect 22560 27532 22612 27538
rect 22560 27474 22612 27480
rect 22480 27402 22600 27418
rect 22480 27396 22612 27402
rect 22480 27390 22560 27396
rect 22560 27338 22612 27344
rect 22468 26852 22520 26858
rect 22468 26794 22520 26800
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22284 25968 22336 25974
rect 22284 25910 22336 25916
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 22296 24954 22324 25094
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22388 23882 22416 25638
rect 22480 25362 22508 26794
rect 22572 26382 22600 27338
rect 22664 26874 22692 31078
rect 22756 29646 22784 34886
rect 22848 34746 22876 35866
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 22836 34740 22888 34746
rect 22836 34682 22888 34688
rect 22834 34640 22890 34649
rect 22834 34575 22890 34584
rect 22848 32910 22876 34575
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 23112 33856 23164 33862
rect 23112 33798 23164 33804
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 23124 33658 23152 33798
rect 23112 33652 23164 33658
rect 23112 33594 23164 33600
rect 23216 33386 23244 33798
rect 23308 33538 23336 35866
rect 23400 33674 23428 36518
rect 23492 33862 23520 43590
rect 23584 43110 23612 44270
rect 24032 43784 24084 43790
rect 24032 43726 24084 43732
rect 23664 43716 23716 43722
rect 23664 43658 23716 43664
rect 23572 43104 23624 43110
rect 23572 43046 23624 43052
rect 23572 42832 23624 42838
rect 23572 42774 23624 42780
rect 23584 39846 23612 42774
rect 23572 39840 23624 39846
rect 23572 39782 23624 39788
rect 23676 39098 23704 43658
rect 23848 43308 23900 43314
rect 23848 43250 23900 43256
rect 23860 42634 23888 43250
rect 24044 42702 24072 43726
rect 24032 42696 24084 42702
rect 24032 42638 24084 42644
rect 23848 42628 23900 42634
rect 23848 42570 23900 42576
rect 23860 42294 23888 42570
rect 23848 42288 23900 42294
rect 23848 42230 23900 42236
rect 23860 41682 23888 42230
rect 23848 41676 23900 41682
rect 23848 41618 23900 41624
rect 23940 41268 23992 41274
rect 23940 41210 23992 41216
rect 23756 41064 23808 41070
rect 23756 41006 23808 41012
rect 23768 40526 23796 41006
rect 23756 40520 23808 40526
rect 23756 40462 23808 40468
rect 23756 39500 23808 39506
rect 23756 39442 23808 39448
rect 23664 39092 23716 39098
rect 23664 39034 23716 39040
rect 23572 38752 23624 38758
rect 23572 38694 23624 38700
rect 23584 38554 23612 38694
rect 23572 38548 23624 38554
rect 23572 38490 23624 38496
rect 23676 37942 23704 39034
rect 23768 38010 23796 39442
rect 23848 38208 23900 38214
rect 23848 38150 23900 38156
rect 23756 38004 23808 38010
rect 23756 37946 23808 37952
rect 23664 37936 23716 37942
rect 23664 37878 23716 37884
rect 23676 37806 23704 37878
rect 23664 37800 23716 37806
rect 23664 37742 23716 37748
rect 23676 37466 23704 37742
rect 23664 37460 23716 37466
rect 23664 37402 23716 37408
rect 23676 36854 23704 37402
rect 23664 36848 23716 36854
rect 23664 36790 23716 36796
rect 23860 36174 23888 38150
rect 23952 37346 23980 41210
rect 24044 38894 24072 42638
rect 24032 38888 24084 38894
rect 24032 38830 24084 38836
rect 24136 37466 24164 47058
rect 24492 46980 24544 46986
rect 24492 46922 24544 46928
rect 24504 45665 24532 46922
rect 24490 45656 24546 45665
rect 24490 45591 24546 45600
rect 24492 45416 24544 45422
rect 24492 45358 24544 45364
rect 24504 44033 24532 45358
rect 24490 44024 24546 44033
rect 24490 43959 24546 43968
rect 24596 43654 24624 53926
rect 24780 53582 24808 54567
rect 25320 54188 25372 54194
rect 25320 54130 25372 54136
rect 25332 53825 25360 54130
rect 25964 53984 26016 53990
rect 25964 53926 26016 53932
rect 25318 53816 25374 53825
rect 25240 53774 25318 53802
rect 24768 53576 24820 53582
rect 24768 53518 24820 53524
rect 24780 52698 24808 53518
rect 25136 53440 25188 53446
rect 25136 53382 25188 53388
rect 24768 52692 24820 52698
rect 24768 52634 24820 52640
rect 24860 51264 24912 51270
rect 24860 51206 24912 51212
rect 24768 45416 24820 45422
rect 24768 45358 24820 45364
rect 24780 44441 24808 45358
rect 24766 44432 24822 44441
rect 24766 44367 24822 44376
rect 24676 44328 24728 44334
rect 24768 44328 24820 44334
rect 24676 44270 24728 44276
rect 24766 44296 24768 44305
rect 24820 44296 24822 44305
rect 24688 43858 24716 44270
rect 24766 44231 24822 44240
rect 24676 43852 24728 43858
rect 24676 43794 24728 43800
rect 24584 43648 24636 43654
rect 24584 43590 24636 43596
rect 24688 43217 24716 43794
rect 24674 43208 24730 43217
rect 24674 43143 24730 43152
rect 24308 43104 24360 43110
rect 24308 43046 24360 43052
rect 24216 41472 24268 41478
rect 24216 41414 24268 41420
rect 24228 40526 24256 41414
rect 24216 40520 24268 40526
rect 24216 40462 24268 40468
rect 24320 40458 24348 43046
rect 24490 42392 24546 42401
rect 24490 42327 24546 42336
rect 24400 42288 24452 42294
rect 24400 42230 24452 42236
rect 24308 40452 24360 40458
rect 24308 40394 24360 40400
rect 24320 38962 24348 40394
rect 24308 38956 24360 38962
rect 24308 38898 24360 38904
rect 24308 38752 24360 38758
rect 24308 38694 24360 38700
rect 24216 37868 24268 37874
rect 24216 37810 24268 37816
rect 24228 37466 24256 37810
rect 24124 37460 24176 37466
rect 24124 37402 24176 37408
rect 24216 37460 24268 37466
rect 24216 37402 24268 37408
rect 23952 37318 24256 37346
rect 24032 37256 24084 37262
rect 24032 37198 24084 37204
rect 24124 37256 24176 37262
rect 24124 37198 24176 37204
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 23572 36100 23624 36106
rect 23572 36042 23624 36048
rect 23940 36100 23992 36106
rect 23940 36042 23992 36048
rect 23584 35894 23612 36042
rect 23584 35866 23704 35894
rect 23584 35222 23612 35866
rect 23676 35834 23704 35866
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 23952 35290 23980 36042
rect 24044 35630 24072 37198
rect 24032 35624 24084 35630
rect 24032 35566 24084 35572
rect 23940 35284 23992 35290
rect 23940 35226 23992 35232
rect 23572 35216 23624 35222
rect 23572 35158 23624 35164
rect 24136 35154 24164 37198
rect 24124 35148 24176 35154
rect 24124 35090 24176 35096
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23480 33856 23532 33862
rect 23480 33798 23532 33804
rect 23400 33646 23520 33674
rect 23308 33510 23428 33538
rect 23296 33448 23348 33454
rect 23296 33390 23348 33396
rect 23204 33380 23256 33386
rect 23204 33322 23256 33328
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22848 30734 22876 32166
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23308 31890 23336 33390
rect 23296 31884 23348 31890
rect 23296 31826 23348 31832
rect 23308 31482 23336 31826
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 23400 31414 23428 33510
rect 23492 33114 23520 33646
rect 23480 33108 23532 33114
rect 23480 33050 23532 33056
rect 23572 32496 23624 32502
rect 23572 32438 23624 32444
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 23388 31408 23440 31414
rect 23388 31350 23440 31356
rect 23492 31278 23520 32370
rect 23480 31272 23532 31278
rect 23480 31214 23532 31220
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22928 30864 22980 30870
rect 22928 30806 22980 30812
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 22940 30036 22968 30806
rect 23492 30802 23520 31214
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 23296 30592 23348 30598
rect 23296 30534 23348 30540
rect 22848 30008 22968 30036
rect 22848 29832 22876 30008
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23308 29850 23336 30534
rect 23296 29844 23348 29850
rect 22848 29804 22968 29832
rect 22940 29714 22968 29804
rect 23296 29786 23348 29792
rect 22928 29708 22980 29714
rect 22928 29650 22980 29656
rect 23480 29708 23532 29714
rect 23480 29650 23532 29656
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22744 28756 22796 28762
rect 22744 28698 22796 28704
rect 22756 26994 22784 28698
rect 23020 28484 23072 28490
rect 23020 28426 23072 28432
rect 23032 28014 23060 28426
rect 23308 28218 23336 28970
rect 23492 28422 23520 29650
rect 23584 29050 23612 32438
rect 23676 30258 23704 34478
rect 24044 34406 24072 35022
rect 24228 34610 24256 37318
rect 24320 34610 24348 38694
rect 24412 38554 24440 42230
rect 24504 41750 24532 42327
rect 24872 42090 24900 51206
rect 25044 47592 25096 47598
rect 25044 47534 25096 47540
rect 25056 47025 25084 47534
rect 25042 47016 25098 47025
rect 25042 46951 25098 46960
rect 25044 46368 25096 46374
rect 25044 46310 25096 46316
rect 24952 45892 25004 45898
rect 24952 45834 25004 45840
rect 24964 45082 24992 45834
rect 24952 45076 25004 45082
rect 24952 45018 25004 45024
rect 24952 43648 25004 43654
rect 24952 43590 25004 43596
rect 24964 43382 24992 43590
rect 24952 43376 25004 43382
rect 24952 43318 25004 43324
rect 24860 42084 24912 42090
rect 24860 42026 24912 42032
rect 24492 41744 24544 41750
rect 24492 41686 24544 41692
rect 24504 41138 24532 41686
rect 25056 41682 25084 46310
rect 24768 41676 24820 41682
rect 24768 41618 24820 41624
rect 25044 41676 25096 41682
rect 25044 41618 25096 41624
rect 24584 41472 24636 41478
rect 24584 41414 24636 41420
rect 24492 41132 24544 41138
rect 24492 41074 24544 41080
rect 24492 40520 24544 40526
rect 24492 40462 24544 40468
rect 24400 38548 24452 38554
rect 24400 38490 24452 38496
rect 24400 38344 24452 38350
rect 24400 38286 24452 38292
rect 24412 38010 24440 38286
rect 24400 38004 24452 38010
rect 24400 37946 24452 37952
rect 24412 37262 24440 37946
rect 24504 37505 24532 40462
rect 24596 39030 24624 41414
rect 24780 40118 24808 41618
rect 25044 41540 25096 41546
rect 25044 41482 25096 41488
rect 24952 41472 25004 41478
rect 24952 41414 25004 41420
rect 24860 40928 24912 40934
rect 24860 40870 24912 40876
rect 24872 40769 24900 40870
rect 24858 40760 24914 40769
rect 24858 40695 24914 40704
rect 24964 40186 24992 41414
rect 24952 40180 25004 40186
rect 24952 40122 25004 40128
rect 24768 40112 24820 40118
rect 25056 40066 25084 41482
rect 25148 40730 25176 53382
rect 25240 52154 25268 53774
rect 25318 53751 25374 53760
rect 25320 53100 25372 53106
rect 25320 53042 25372 53048
rect 25332 53009 25360 53042
rect 25318 53000 25374 53009
rect 25318 52935 25374 52944
rect 25688 52896 25740 52902
rect 25688 52838 25740 52844
rect 25320 52488 25372 52494
rect 25320 52430 25372 52436
rect 25332 52193 25360 52430
rect 25318 52184 25374 52193
rect 25228 52148 25280 52154
rect 25318 52119 25374 52128
rect 25228 52090 25280 52096
rect 25320 51808 25372 51814
rect 25320 51750 25372 51756
rect 25332 51406 25360 51750
rect 25320 51400 25372 51406
rect 25318 51368 25320 51377
rect 25372 51368 25374 51377
rect 25318 51303 25374 51312
rect 25700 51074 25728 52838
rect 25780 52624 25832 52630
rect 25780 52566 25832 52572
rect 25608 51046 25728 51074
rect 25320 50924 25372 50930
rect 25320 50866 25372 50872
rect 25332 50561 25360 50866
rect 25504 50720 25556 50726
rect 25504 50662 25556 50668
rect 25318 50552 25374 50561
rect 25318 50487 25374 50496
rect 25412 50380 25464 50386
rect 25412 50322 25464 50328
rect 25320 50312 25372 50318
rect 25320 50254 25372 50260
rect 25332 49745 25360 50254
rect 25424 49774 25452 50322
rect 25412 49768 25464 49774
rect 25318 49736 25374 49745
rect 25412 49710 25464 49716
rect 25318 49671 25374 49680
rect 25320 49224 25372 49230
rect 25320 49166 25372 49172
rect 25332 48929 25360 49166
rect 25318 48920 25374 48929
rect 25318 48855 25374 48864
rect 25228 48680 25280 48686
rect 25228 48622 25280 48628
rect 25240 48006 25268 48622
rect 25424 48113 25452 49710
rect 25410 48104 25466 48113
rect 25410 48039 25466 48048
rect 25228 48000 25280 48006
rect 25228 47942 25280 47948
rect 25320 48000 25372 48006
rect 25320 47942 25372 47948
rect 25240 46481 25268 47942
rect 25332 47598 25360 47942
rect 25320 47592 25372 47598
rect 25320 47534 25372 47540
rect 25332 47297 25360 47534
rect 25318 47288 25374 47297
rect 25318 47223 25374 47232
rect 25320 46912 25372 46918
rect 25320 46854 25372 46860
rect 25332 46510 25360 46854
rect 25320 46504 25372 46510
rect 25226 46472 25282 46481
rect 25320 46446 25372 46452
rect 25226 46407 25282 46416
rect 25332 44849 25360 46446
rect 25318 44840 25374 44849
rect 25318 44775 25374 44784
rect 25320 43240 25372 43246
rect 25320 43182 25372 43188
rect 25332 42770 25360 43182
rect 25320 42764 25372 42770
rect 25320 42706 25372 42712
rect 25228 42696 25280 42702
rect 25228 42638 25280 42644
rect 25240 41818 25268 42638
rect 25332 42090 25360 42706
rect 25320 42084 25372 42090
rect 25320 42026 25372 42032
rect 25228 41812 25280 41818
rect 25228 41754 25280 41760
rect 25136 40724 25188 40730
rect 25136 40666 25188 40672
rect 25228 40384 25280 40390
rect 25228 40326 25280 40332
rect 24768 40054 24820 40060
rect 24676 39432 24728 39438
rect 24676 39374 24728 39380
rect 24584 39024 24636 39030
rect 24584 38966 24636 38972
rect 24490 37496 24546 37505
rect 24490 37431 24546 37440
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24688 36922 24716 39374
rect 24780 39302 24808 40054
rect 24872 40038 25084 40066
rect 24768 39296 24820 39302
rect 24768 39238 24820 39244
rect 24780 38894 24808 39238
rect 24768 38888 24820 38894
rect 24768 38830 24820 38836
rect 24768 37868 24820 37874
rect 24768 37810 24820 37816
rect 24676 36916 24728 36922
rect 24676 36858 24728 36864
rect 24688 36310 24716 36858
rect 24676 36304 24728 36310
rect 24676 36246 24728 36252
rect 24492 36032 24544 36038
rect 24492 35974 24544 35980
rect 24584 36032 24636 36038
rect 24584 35974 24636 35980
rect 24400 35760 24452 35766
rect 24400 35702 24452 35708
rect 24412 34898 24440 35702
rect 24504 35086 24532 35974
rect 24492 35080 24544 35086
rect 24492 35022 24544 35028
rect 24412 34870 24532 34898
rect 24400 34740 24452 34746
rect 24400 34682 24452 34688
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 24032 34400 24084 34406
rect 24032 34342 24084 34348
rect 23848 33584 23900 33590
rect 23848 33526 23900 33532
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23768 32570 23796 33390
rect 23860 33114 23888 33526
rect 23848 33108 23900 33114
rect 23848 33050 23900 33056
rect 24124 32836 24176 32842
rect 24124 32778 24176 32784
rect 23756 32564 23808 32570
rect 23756 32506 23808 32512
rect 24032 32292 24084 32298
rect 24032 32234 24084 32240
rect 24044 32026 24072 32234
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 23756 29232 23808 29238
rect 23756 29174 23808 29180
rect 23584 29022 23704 29050
rect 23480 28416 23532 28422
rect 23480 28358 23532 28364
rect 23296 28212 23348 28218
rect 23296 28154 23348 28160
rect 23020 28008 23072 28014
rect 23020 27950 23072 27956
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23294 27568 23350 27577
rect 23294 27503 23350 27512
rect 23308 27130 23336 27503
rect 23400 27470 23428 27814
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 23386 27024 23442 27033
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 23296 26988 23348 26994
rect 23386 26959 23442 26968
rect 23296 26930 23348 26936
rect 22664 26846 22784 26874
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22560 26376 22612 26382
rect 22560 26318 22612 26324
rect 22560 26240 22612 26246
rect 22560 26182 22612 26188
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22468 25220 22520 25226
rect 22468 25162 22520 25168
rect 22296 23854 22416 23882
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 22020 21962 22048 22646
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 22020 21146 22048 21898
rect 22204 21690 22232 22918
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22296 20466 22324 23854
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22388 21894 22416 23666
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22480 20210 22508 25162
rect 22572 21690 22600 26182
rect 22664 21706 22692 26726
rect 22756 26382 22784 26846
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23112 26444 23164 26450
rect 23112 26386 23164 26392
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 23124 25786 23152 26386
rect 23202 26072 23258 26081
rect 23202 26007 23204 26016
rect 23256 26007 23258 26016
rect 23204 25978 23256 25984
rect 23308 25922 23336 26930
rect 23400 26858 23428 26959
rect 23388 26852 23440 26858
rect 23388 26794 23440 26800
rect 23388 26308 23440 26314
rect 23388 26250 23440 26256
rect 23216 25906 23336 25922
rect 23400 25906 23428 26250
rect 23204 25900 23336 25906
rect 23256 25894 23336 25900
rect 23388 25900 23440 25906
rect 23204 25842 23256 25848
rect 23388 25842 23440 25848
rect 22848 24682 22876 25774
rect 23124 25758 23336 25786
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22756 23254 22784 24006
rect 22744 23248 22796 23254
rect 22744 23190 22796 23196
rect 22848 22817 22876 24074
rect 23308 24070 23336 25758
rect 23400 24410 23428 25842
rect 23492 25294 23520 27270
rect 23584 27062 23612 27950
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 23676 26382 23704 29022
rect 23768 26432 23796 29174
rect 23860 29050 23888 31622
rect 23940 30592 23992 30598
rect 23940 30534 23992 30540
rect 23952 29170 23980 30534
rect 24032 30048 24084 30054
rect 24032 29990 24084 29996
rect 23940 29164 23992 29170
rect 23940 29106 23992 29112
rect 23860 29022 23980 29050
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23860 27130 23888 27474
rect 23848 27124 23900 27130
rect 23848 27066 23900 27072
rect 23768 26404 23888 26432
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23756 26308 23808 26314
rect 23756 26250 23808 26256
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23400 24070 23428 24346
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23308 23746 23336 24006
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23308 23718 23520 23746
rect 23308 23662 23336 23718
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23386 23624 23442 23633
rect 23386 23559 23442 23568
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22834 22808 22890 22817
rect 22834 22743 22890 22752
rect 23308 22438 23336 23462
rect 23400 23118 23428 23559
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23204 22094 23256 22098
rect 23308 22094 23336 22374
rect 23204 22092 23336 22094
rect 23256 22066 23336 22092
rect 23204 22034 23256 22040
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22560 21684 22612 21690
rect 22664 21678 22784 21706
rect 22560 21626 22612 21632
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22664 21010 22692 21490
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22296 20182 22508 20210
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 22296 19310 22324 20182
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22296 18970 22324 19246
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22112 17338 22140 17546
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21468 14198 21680 14226
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21376 12306 21404 12650
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21468 12170 21496 13806
rect 21652 12322 21680 14198
rect 21744 12986 21772 15302
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21836 14958 21864 15098
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21652 12294 21772 12322
rect 21744 12238 21772 12294
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20732 6886 20852 6914
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20364 3126 20392 4490
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 20456 800 20484 4014
rect 20824 3534 20852 6886
rect 21008 5234 21036 8298
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21284 4622 21312 11018
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21468 7886 21496 10406
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21468 6322 21496 6598
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21560 5710 21588 11018
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21652 6458 21680 7822
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20732 2514 20760 2994
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 20824 800 20852 2790
rect 21192 800 21220 2926
rect 21376 2922 21404 5578
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 3126 21496 5510
rect 21744 4622 21772 7686
rect 21836 5234 21864 8842
rect 21928 8566 21956 15302
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22020 10062 22048 14010
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22112 12782 22140 13874
rect 22204 13326 22232 16594
rect 22296 15706 22324 18906
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22388 15094 22416 19722
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 16794 22508 17478
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22480 16522 22508 16730
rect 22664 16574 22692 19654
rect 22756 18290 22784 21678
rect 22848 21622 22876 21898
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 23216 21554 23244 22034
rect 23492 21622 23520 23718
rect 23584 22094 23612 23802
rect 23584 22066 23704 22094
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23584 21622 23612 21830
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23584 21146 23612 21558
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23584 20058 23612 21082
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23584 19446 23612 19994
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23584 18714 23612 19382
rect 23492 18698 23612 18714
rect 23480 18692 23612 18698
rect 23532 18686 23612 18692
rect 23480 18634 23532 18640
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22664 16546 22784 16574
rect 22468 16516 22520 16522
rect 22468 16458 22520 16464
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22376 14340 22428 14346
rect 22480 14328 22508 16458
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22428 14300 22508 14328
rect 22376 14282 22428 14288
rect 22388 13394 22416 14282
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22388 12306 22416 12786
rect 22664 12306 22692 15846
rect 22756 15502 22784 16546
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22848 14414 22876 16934
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 13938 22876 14214
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 12850 23336 18022
rect 23388 17060 23440 17066
rect 23388 17002 23440 17008
rect 23400 12850 23428 17002
rect 23492 13938 23520 18090
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23584 15978 23612 17818
rect 23676 17202 23704 22066
rect 23768 19854 23796 26250
rect 23860 24818 23888 26404
rect 23952 25294 23980 29022
rect 24044 26382 24072 29990
rect 24136 28150 24164 32778
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24124 28144 24176 28150
rect 24124 28086 24176 28092
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 24124 26308 24176 26314
rect 24124 26250 24176 26256
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 23940 25152 23992 25158
rect 23940 25094 23992 25100
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23860 22234 23888 22510
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23768 18358 23796 19110
rect 23756 18352 23808 18358
rect 23756 18294 23808 18300
rect 23768 17678 23796 18294
rect 23952 18290 23980 25094
rect 24044 24206 24072 25094
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 24136 23118 24164 26250
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 24124 22704 24176 22710
rect 24124 22646 24176 22652
rect 24136 21894 24164 22646
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 24044 16726 24072 18770
rect 24136 17814 24164 19382
rect 24124 17808 24176 17814
rect 24124 17750 24176 17756
rect 24032 16720 24084 16726
rect 24032 16662 24084 16668
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23848 14884 23900 14890
rect 23848 14826 23900 14832
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 22836 12708 22888 12714
rect 22836 12650 22888 12656
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22098 11928 22154 11937
rect 22098 11863 22154 11872
rect 22112 11830 22140 11863
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22560 11620 22612 11626
rect 22560 11562 22612 11568
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21928 5930 21956 6666
rect 22020 6322 22048 7754
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 21928 5902 22048 5930
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21824 5092 21876 5098
rect 21824 5034 21876 5040
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21560 800 21588 3946
rect 21836 2417 21864 5034
rect 21822 2408 21878 2417
rect 21822 2343 21878 2352
rect 21928 800 21956 5714
rect 22020 3398 22048 5902
rect 22204 5710 22232 9862
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22112 3233 22140 4694
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22204 4049 22232 4082
rect 22190 4040 22246 4049
rect 22190 3975 22246 3984
rect 22098 3224 22154 3233
rect 22098 3159 22154 3168
rect 22296 800 22324 6190
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22480 2990 22508 5102
rect 22572 3058 22600 11562
rect 22848 10146 22876 12650
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22848 10118 22968 10146
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22848 9722 22876 9998
rect 22940 9994 22968 10118
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 23216 9466 23244 9862
rect 23308 9586 23336 12582
rect 23860 11762 23888 14826
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23216 9438 23336 9466
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23308 8650 23336 9438
rect 23400 8974 23428 11562
rect 23952 10674 23980 14282
rect 24228 12918 24256 32370
rect 24308 29028 24360 29034
rect 24308 28970 24360 28976
rect 24320 28529 24348 28970
rect 24412 28558 24440 34682
rect 24504 33590 24532 34870
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 24504 31754 24532 33526
rect 24492 31748 24544 31754
rect 24492 31690 24544 31696
rect 24504 31414 24532 31690
rect 24492 31408 24544 31414
rect 24492 31350 24544 31356
rect 24504 30258 24532 31350
rect 24596 30734 24624 35974
rect 24676 35624 24728 35630
rect 24676 35566 24728 35572
rect 24688 35290 24716 35566
rect 24676 35284 24728 35290
rect 24676 35226 24728 35232
rect 24780 35057 24808 37810
rect 24872 36582 24900 40038
rect 25044 39976 25096 39982
rect 25044 39918 25096 39924
rect 25056 39642 25084 39918
rect 25044 39636 25096 39642
rect 25044 39578 25096 39584
rect 25240 39370 25268 40326
rect 25332 40050 25360 42026
rect 25412 42016 25464 42022
rect 25412 41958 25464 41964
rect 25320 40044 25372 40050
rect 25320 39986 25372 39992
rect 25424 39953 25452 41958
rect 25516 40594 25544 50662
rect 25608 41546 25636 51046
rect 25688 43920 25740 43926
rect 25688 43862 25740 43868
rect 25596 41540 25648 41546
rect 25596 41482 25648 41488
rect 25504 40588 25556 40594
rect 25504 40530 25556 40536
rect 25410 39944 25466 39953
rect 25410 39879 25466 39888
rect 25228 39364 25280 39370
rect 25228 39306 25280 39312
rect 25228 38344 25280 38350
rect 25228 38286 25280 38292
rect 25044 37120 25096 37126
rect 25044 37062 25096 37068
rect 25056 36854 25084 37062
rect 25044 36848 25096 36854
rect 25044 36790 25096 36796
rect 25044 36712 25096 36718
rect 25096 36660 25176 36666
rect 25044 36654 25176 36660
rect 25056 36638 25176 36654
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 24952 36576 25004 36582
rect 24952 36518 25004 36524
rect 24964 36242 24992 36518
rect 25044 36372 25096 36378
rect 25044 36314 25096 36320
rect 24952 36236 25004 36242
rect 24952 36178 25004 36184
rect 24964 35630 24992 36178
rect 24952 35624 25004 35630
rect 24952 35566 25004 35572
rect 24766 35048 24822 35057
rect 24766 34983 24822 34992
rect 24768 34740 24820 34746
rect 24768 34682 24820 34688
rect 24676 32768 24728 32774
rect 24676 32710 24728 32716
rect 24688 32434 24716 32710
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24688 29510 24716 29582
rect 24676 29504 24728 29510
rect 24676 29446 24728 29452
rect 24400 28552 24452 28558
rect 24306 28520 24362 28529
rect 24400 28494 24452 28500
rect 24306 28455 24362 28464
rect 24308 28416 24360 28422
rect 24308 28358 24360 28364
rect 24320 27470 24348 28358
rect 24584 27940 24636 27946
rect 24584 27882 24636 27888
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 24320 25362 24348 27406
rect 24492 27328 24544 27334
rect 24492 27270 24544 27276
rect 24504 25974 24532 27270
rect 24492 25968 24544 25974
rect 24492 25910 24544 25916
rect 24308 25356 24360 25362
rect 24308 25298 24360 25304
rect 24400 24132 24452 24138
rect 24400 24074 24452 24080
rect 24308 21956 24360 21962
rect 24308 21898 24360 21904
rect 24320 16114 24348 21898
rect 24412 19854 24440 24074
rect 24596 21876 24624 27882
rect 24688 26897 24716 29446
rect 24780 29238 24808 34682
rect 24858 34232 24914 34241
rect 24858 34167 24860 34176
rect 24912 34167 24914 34176
rect 24860 34138 24912 34144
rect 24964 33318 24992 35566
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 25056 33114 25084 36314
rect 25148 35630 25176 36638
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25044 33108 25096 33114
rect 25044 33050 25096 33056
rect 24952 32836 25004 32842
rect 24952 32778 25004 32784
rect 24964 32609 24992 32778
rect 24950 32600 25006 32609
rect 24950 32535 25006 32544
rect 25148 32366 25176 34342
rect 25240 33658 25268 38286
rect 25504 37664 25556 37670
rect 25504 37606 25556 37612
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25332 34610 25360 35430
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 25332 33425 25360 34546
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 25318 33416 25374 33425
rect 25318 33351 25374 33360
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 24952 31680 25004 31686
rect 24952 31622 25004 31628
rect 24964 31414 24992 31622
rect 24952 31408 25004 31414
rect 24952 31350 25004 31356
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24768 29232 24820 29238
rect 24768 29174 24820 29180
rect 24674 26888 24730 26897
rect 24674 26823 24730 26832
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24674 25256 24730 25265
rect 24674 25191 24730 25200
rect 24688 24750 24716 25191
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24688 23798 24716 24006
rect 24676 23792 24728 23798
rect 24676 23734 24728 23740
rect 24780 22574 24808 25774
rect 24872 25294 24900 30534
rect 25240 30394 25268 32302
rect 25332 30977 25360 32846
rect 25424 31793 25452 33934
rect 25410 31784 25466 31793
rect 25410 31719 25466 31728
rect 25516 31278 25544 37606
rect 25596 35624 25648 35630
rect 25596 35566 25648 35572
rect 25608 32366 25636 35566
rect 25596 32360 25648 32366
rect 25596 32302 25648 32308
rect 25504 31272 25556 31278
rect 25504 31214 25556 31220
rect 25318 30968 25374 30977
rect 25318 30903 25374 30912
rect 25228 30388 25280 30394
rect 25228 30330 25280 30336
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 25412 30320 25464 30326
rect 25412 30262 25464 30268
rect 24964 30161 24992 30262
rect 24950 30152 25006 30161
rect 24950 30087 25006 30096
rect 25424 29850 25452 30262
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 24952 29572 25004 29578
rect 24952 29514 25004 29520
rect 24964 29345 24992 29514
rect 24950 29336 25006 29345
rect 24950 29271 25006 29280
rect 25136 28484 25188 28490
rect 25136 28426 25188 28432
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24872 24449 24900 24618
rect 24858 24440 24914 24449
rect 24858 24375 24914 24384
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24952 22024 25004 22030
rect 24766 21992 24822 22001
rect 24952 21966 25004 21972
rect 24766 21927 24822 21936
rect 24504 21848 24624 21876
rect 24504 20942 24532 21848
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24780 20398 24808 21927
rect 24964 21350 24992 21966
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24858 21176 24914 21185
rect 24858 21111 24914 21120
rect 24872 21010 24900 21111
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 25148 20466 25176 28426
rect 25700 27033 25728 43862
rect 25792 42838 25820 52566
rect 25976 51074 26004 53926
rect 25976 51046 26096 51074
rect 25872 48748 25924 48754
rect 25872 48690 25924 48696
rect 25780 42832 25832 42838
rect 25780 42774 25832 42780
rect 25884 38826 25912 48690
rect 25964 46572 26016 46578
rect 25964 46514 26016 46520
rect 25872 38820 25924 38826
rect 25872 38762 25924 38768
rect 25976 37194 26004 46514
rect 26068 43178 26096 51046
rect 26056 43172 26108 43178
rect 26056 43114 26108 43120
rect 25964 37188 26016 37194
rect 25964 37130 26016 37136
rect 25686 27024 25742 27033
rect 25686 26959 25742 26968
rect 25228 22976 25280 22982
rect 25228 22918 25280 22924
rect 25240 20874 25268 22918
rect 25228 20868 25280 20874
rect 25228 20810 25280 20816
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24768 20392 24820 20398
rect 24872 20369 24900 20402
rect 24768 20334 24820 20340
rect 24858 20360 24914 20369
rect 24858 20295 24914 20304
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24412 19378 24440 19790
rect 24872 19553 24900 19858
rect 24858 19544 24914 19553
rect 24858 19479 24914 19488
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24412 15162 24440 19314
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 25134 18728 25190 18737
rect 24596 17882 24624 18702
rect 25134 18663 25190 18672
rect 25148 18358 25176 18663
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 25134 17912 25190 17921
rect 24584 17876 24636 17882
rect 25134 17847 25190 17856
rect 24584 17818 24636 17824
rect 25148 17270 25176 17847
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25136 17264 25188 17270
rect 25136 17206 25188 17212
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 24674 16280 24730 16289
rect 24674 16215 24730 16224
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24688 14958 24716 16215
rect 24780 16046 24808 17031
rect 25240 16794 25268 17478
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 25502 15464 25558 15473
rect 25502 15399 25504 15408
rect 25556 15399 25558 15408
rect 25504 15370 25556 15376
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 25134 14648 25190 14657
rect 25134 14583 25190 14592
rect 25148 14006 25176 14583
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23308 8622 23428 8650
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22664 3738 22692 8366
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 22848 4049 22876 6122
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23020 5636 23072 5642
rect 23020 5578 23072 5584
rect 23032 5302 23060 5578
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22834 4040 22890 4049
rect 22834 3975 22890 3984
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22664 800 22692 2858
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23032 870 23152 898
rect 23032 800 23060 870
rect 13188 734 13400 762
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23124 762 23152 870
rect 23308 762 23336 7890
rect 23400 7478 23428 8622
rect 23492 8498 23520 10406
rect 23952 9586 23980 10474
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 24596 9466 24624 12854
rect 24780 12782 24808 13767
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25516 13025 25544 13194
rect 25502 13016 25558 13025
rect 25502 12951 25558 12960
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24766 11384 24822 11393
rect 24766 11319 24822 11328
rect 24780 10606 24808 11319
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24766 10432 24822 10441
rect 24766 10367 24822 10376
rect 24780 9518 24808 10367
rect 24768 9512 24820 9518
rect 24596 9438 24716 9466
rect 24768 9454 24820 9460
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23400 4865 23428 7278
rect 23952 6322 23980 8774
rect 24044 6798 24072 8774
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 24136 5234 24164 7686
rect 24596 6798 24624 9318
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 23386 4856 23442 4865
rect 23386 4791 23442 4800
rect 23754 3496 23810 3505
rect 23754 3431 23810 3440
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23400 800 23428 3334
rect 23768 800 23796 3431
rect 24688 2650 24716 9438
rect 24872 7886 24900 12038
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24964 9761 24992 9998
rect 24950 9752 25006 9761
rect 24950 9687 25006 9696
rect 25056 8974 25084 12310
rect 25134 12200 25190 12209
rect 25134 12135 25190 12144
rect 25148 11830 25176 12135
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 25148 8566 25176 8871
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 24766 7304 24822 7313
rect 24766 7239 24822 7248
rect 24780 6254 24808 7239
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24872 6497 24900 6802
rect 24858 6488 24914 6497
rect 24858 6423 24914 6432
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24766 5672 24822 5681
rect 24766 5607 24822 5616
rect 24780 5166 24808 5607
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 24676 2644 24728 2650
rect 24676 2586 24728 2592
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24136 800 24164 2314
rect 23124 734 23336 762
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 24964 785 24992 3674
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25056 1601 25084 2382
rect 25042 1592 25098 1601
rect 25042 1527 25098 1536
rect 24950 776 25006 785
rect 24950 711 25006 720
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2962 52964 3018 53000
rect 2962 52944 2964 52964
rect 2964 52944 3016 52964
rect 3016 52944 3018 52964
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 3974 55392 4030 55448
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 3330 50360 3386 50416
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 1306 43152 1362 43208
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 1306 40704 1362 40760
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 1306 38292 1308 38312
rect 1308 38292 1360 38312
rect 1360 38292 1362 38312
rect 1306 38256 1362 38292
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 1582 35808 1638 35864
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 1214 33360 1270 33416
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2778 30912 2834 30968
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2870 28464 2926 28520
rect 2778 26016 2834 26072
rect 1306 21120 1362 21176
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 4066 48048 4122 48104
rect 3974 45620 4030 45656
rect 3974 45600 3976 45620
rect 3976 45600 4028 45620
rect 4028 45600 4030 45620
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2870 23568 2926 23624
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 6366 42200 6422 42256
rect 4894 26288 4950 26344
rect 1306 18672 1362 18728
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 1306 16224 1362 16280
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 938 13812 940 13832
rect 940 13812 992 13832
rect 992 13812 994 13832
rect 938 13776 994 13812
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2778 11328 2834 11384
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2870 8880 2926 8936
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3146 6432 3202 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 1398 1536 1454 1592
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3330 3440 3386 3496
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 4066 3984 4122 4040
rect 4066 2644 4122 2680
rect 4066 2624 4068 2644
rect 4068 2624 4120 2644
rect 4120 2624 4122 2644
rect 5262 3612 5264 3632
rect 5264 3612 5316 3632
rect 5316 3612 5318 3632
rect 5262 3576 5318 3612
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 9218 44240 9274 44296
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 9402 36624 9458 36680
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 9034 26732 9036 26752
rect 9036 26732 9088 26752
rect 9088 26732 9090 26752
rect 9034 26696 9090 26732
rect 10506 44648 10562 44704
rect 10138 39480 10194 39536
rect 11242 44648 11298 44704
rect 11610 44260 11666 44296
rect 11610 44240 11612 44260
rect 11612 44240 11664 44260
rect 11664 44240 11666 44260
rect 10966 39344 11022 39400
rect 11058 34856 11114 34912
rect 11150 34740 11206 34776
rect 11150 34720 11152 34740
rect 11152 34720 11204 34740
rect 11204 34720 11206 34740
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12254 45228 12256 45248
rect 12256 45228 12308 45248
rect 12308 45228 12310 45248
rect 12254 45192 12310 45228
rect 14002 52536 14058 52592
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 10230 25100 10232 25120
rect 10232 25100 10284 25120
rect 10284 25100 10286 25120
rect 10230 25064 10286 25100
rect 10138 21292 10140 21312
rect 10140 21292 10192 21312
rect 10192 21292 10194 21312
rect 10138 21256 10194 21292
rect 10506 19796 10508 19816
rect 10508 19796 10560 19816
rect 10560 19796 10562 19816
rect 10506 19760 10562 19796
rect 10046 10920 10102 10976
rect 9218 7928 9274 7984
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 8390 3188 8446 3224
rect 8390 3168 8392 3188
rect 8392 3168 8444 3188
rect 8444 3168 8446 3188
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 10782 17312 10838 17368
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12438 38936 12494 38992
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12898 39480 12954 39536
rect 12346 38820 12402 38856
rect 12346 38800 12348 38820
rect 12348 38800 12400 38820
rect 12400 38800 12402 38820
rect 12254 38392 12310 38448
rect 12990 39344 13046 39400
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 13450 41132 13506 41168
rect 13450 41112 13452 41132
rect 13452 41112 13504 41132
rect 13504 41112 13506 41132
rect 13450 38936 13506 38992
rect 12714 35672 12770 35728
rect 11518 22616 11574 22672
rect 12346 30368 12402 30424
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 13358 33380 13414 33416
rect 13358 33360 13360 33380
rect 13360 33360 13412 33380
rect 13412 33360 13414 33380
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 14002 40724 14058 40760
rect 14002 40704 14004 40724
rect 14004 40704 14056 40724
rect 14056 40704 14058 40724
rect 13358 32272 13414 32328
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 14186 34040 14242 34096
rect 14094 33260 14096 33280
rect 14096 33260 14148 33280
rect 14148 33260 14150 33280
rect 14094 33224 14150 33260
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12346 29280 12402 29336
rect 12530 23160 12586 23216
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12438 17312 12494 17368
rect 12162 12980 12218 13016
rect 12162 12960 12164 12980
rect 12164 12960 12216 12980
rect 12216 12960 12218 12980
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 14002 21292 14004 21312
rect 14004 21292 14056 21312
rect 14056 21292 14058 21312
rect 14002 21256 14058 21292
rect 15382 38820 15438 38856
rect 15382 38800 15384 38820
rect 15384 38800 15436 38820
rect 15436 38800 15438 38820
rect 15382 38412 15438 38448
rect 15382 38392 15384 38412
rect 15384 38392 15436 38412
rect 15436 38392 15438 38412
rect 15658 38800 15714 38856
rect 14922 26424 14978 26480
rect 13634 17604 13690 17640
rect 13634 17584 13636 17604
rect 13636 17584 13688 17604
rect 13688 17584 13690 17604
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12898 13388 12954 13424
rect 12898 13368 12900 13388
rect 12900 13368 12952 13388
rect 12952 13368 12954 13388
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13542 11600 13598 11656
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 13726 11328 13782 11384
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14738 21256 14794 21312
rect 14738 18420 14794 18456
rect 14738 18400 14740 18420
rect 14740 18400 14792 18420
rect 14792 18400 14794 18420
rect 15198 26560 15254 26616
rect 15842 39480 15898 39536
rect 17038 53932 17040 53952
rect 17040 53932 17092 53952
rect 17092 53932 17094 53952
rect 17038 53896 17094 53932
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 24490 56208 24546 56264
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 16670 39072 16726 39128
rect 16394 37032 16450 37088
rect 16026 31356 16028 31376
rect 16028 31356 16080 31376
rect 16080 31356 16082 31376
rect 16026 31320 16082 31356
rect 15014 20340 15016 20360
rect 15016 20340 15068 20360
rect 15068 20340 15070 20360
rect 15014 20304 15070 20340
rect 15014 15272 15070 15328
rect 15658 28056 15714 28112
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 18234 47096 18290 47152
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17406 40704 17462 40760
rect 16394 28056 16450 28112
rect 16394 26580 16450 26616
rect 16394 26560 16396 26580
rect 16396 26560 16448 26580
rect 16448 26560 16450 26580
rect 15750 20324 15806 20360
rect 15750 20304 15752 20324
rect 15752 20304 15804 20324
rect 15804 20304 15806 20324
rect 16762 29028 16818 29064
rect 16762 29008 16764 29028
rect 16764 29008 16816 29028
rect 16816 29008 16818 29028
rect 16854 27668 16910 27704
rect 16854 27648 16856 27668
rect 16856 27648 16908 27668
rect 16908 27648 16910 27668
rect 16762 26152 16818 26208
rect 16486 19932 16488 19952
rect 16488 19932 16540 19952
rect 16540 19932 16542 19952
rect 16486 19896 16542 19932
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17498 34448 17554 34504
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 19246 47096 19302 47152
rect 19614 46996 19616 47016
rect 19616 46996 19668 47016
rect 19668 46996 19670 47016
rect 19614 46960 19670 46996
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17682 38528 17738 38584
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17682 33224 17738 33280
rect 17130 26424 17186 26480
rect 17406 30096 17462 30152
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17866 28076 17922 28112
rect 17866 28056 17868 28076
rect 17868 28056 17920 28076
rect 17920 28056 17922 28076
rect 17314 26968 17370 27024
rect 17682 26696 17738 26752
rect 17774 26288 17830 26344
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 16394 16788 16450 16824
rect 16394 16768 16396 16788
rect 16396 16768 16448 16788
rect 16448 16768 16450 16788
rect 16026 13232 16082 13288
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17498 15156 17554 15192
rect 17498 15136 17500 15156
rect 17500 15136 17552 15156
rect 17552 15136 17554 15156
rect 17498 13268 17500 13288
rect 17500 13268 17552 13288
rect 17552 13268 17554 13288
rect 17498 13232 17554 13268
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18970 30368 19026 30424
rect 19430 34604 19486 34640
rect 19430 34584 19432 34604
rect 19432 34584 19484 34604
rect 19484 34584 19486 34604
rect 18878 27820 18880 27840
rect 18880 27820 18932 27840
rect 18932 27820 18934 27840
rect 18878 27784 18934 27820
rect 19982 41112 20038 41168
rect 19982 40024 20038 40080
rect 20258 39788 20260 39808
rect 20260 39788 20312 39808
rect 20312 39788 20314 39808
rect 20258 39752 20314 39788
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18602 19352 18658 19408
rect 18786 21120 18842 21176
rect 18694 18808 18750 18864
rect 18418 17992 18474 18048
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19798 30660 19854 30696
rect 19798 30640 19800 30660
rect 19800 30640 19852 30660
rect 19852 30640 19854 30660
rect 22282 53932 22284 53952
rect 22284 53932 22336 53952
rect 22336 53932 22338 53952
rect 21362 43052 21364 43072
rect 21364 43052 21416 43072
rect 21416 43052 21418 43072
rect 21362 43016 21418 43052
rect 21178 41148 21180 41168
rect 21180 41148 21232 41168
rect 21232 41148 21234 41168
rect 21178 41112 21234 41148
rect 20626 37304 20682 37360
rect 19706 28212 19762 28248
rect 19706 28192 19708 28212
rect 19708 28192 19760 28212
rect 19760 28192 19762 28212
rect 19706 27276 19708 27296
rect 19708 27276 19760 27296
rect 19760 27276 19762 27296
rect 19706 27240 19762 27276
rect 21454 39752 21510 39808
rect 22282 53896 22338 53932
rect 21822 44684 21824 44704
rect 21824 44684 21876 44704
rect 21876 44684 21878 44704
rect 21822 44648 21878 44684
rect 21914 39752 21970 39808
rect 21822 39072 21878 39128
rect 21178 31476 21234 31512
rect 21178 31456 21180 31476
rect 21180 31456 21232 31476
rect 21232 31456 21234 31476
rect 18786 3984 18842 4040
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 20350 12824 20406 12880
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 24674 55392 24730 55448
rect 24766 54576 24822 54632
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 23846 52536 23902 52592
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22190 41520 22246 41576
rect 22190 38256 22246 38312
rect 22466 41132 22522 41168
rect 22466 41112 22468 41132
rect 22468 41112 22520 41132
rect 22520 41112 22522 41132
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22834 41112 22890 41168
rect 22466 40024 22522 40080
rect 22558 39788 22560 39808
rect 22560 39788 22612 39808
rect 22612 39788 22614 39808
rect 22558 39752 22614 39788
rect 22466 38700 22468 38720
rect 22468 38700 22520 38720
rect 22520 38700 22522 38720
rect 22466 38664 22522 38700
rect 22190 38004 22246 38040
rect 22190 37984 22192 38004
rect 22192 37984 22244 38004
rect 22244 37984 22246 38004
rect 22190 36916 22246 36952
rect 22190 36896 22192 36916
rect 22192 36896 22244 36916
rect 22244 36896 22246 36916
rect 22190 36644 22246 36680
rect 22190 36624 22192 36644
rect 22192 36624 22244 36644
rect 22244 36624 22246 36644
rect 22282 36080 22338 36136
rect 21914 32000 21970 32056
rect 22374 35808 22430 35864
rect 22742 37984 22798 38040
rect 22742 36080 22798 36136
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 23294 38392 23350 38448
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22834 34584 22890 34640
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 24490 45600 24546 45656
rect 24490 43968 24546 44024
rect 24766 44376 24822 44432
rect 24766 44276 24768 44296
rect 24768 44276 24820 44296
rect 24820 44276 24822 44296
rect 24766 44240 24822 44276
rect 24674 43152 24730 43208
rect 24490 42336 24546 42392
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 25042 46960 25098 47016
rect 24858 40704 24914 40760
rect 25318 53760 25374 53816
rect 25318 52944 25374 53000
rect 25318 52128 25374 52184
rect 25318 51348 25320 51368
rect 25320 51348 25372 51368
rect 25372 51348 25374 51368
rect 25318 51312 25374 51348
rect 25318 50496 25374 50552
rect 25318 49680 25374 49736
rect 25318 48864 25374 48920
rect 25410 48048 25466 48104
rect 25318 47232 25374 47288
rect 25226 46416 25282 46472
rect 25318 44784 25374 44840
rect 24490 37440 24546 37496
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 23294 27512 23350 27568
rect 23386 26968 23442 27024
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 23202 26036 23258 26072
rect 23202 26016 23204 26036
rect 23204 26016 23256 26036
rect 23256 26016 23258 26036
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 23386 23568 23442 23624
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22834 22752 22890 22808
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22098 11872 22154 11928
rect 21822 2352 21878 2408
rect 22190 3984 22246 4040
rect 22098 3168 22154 3224
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 25410 39888 25466 39944
rect 24766 34992 24822 35048
rect 24306 28464 24362 28520
rect 24858 34196 24914 34232
rect 24858 34176 24860 34196
rect 24860 34176 24912 34196
rect 24912 34176 24914 34196
rect 24950 32544 25006 32600
rect 25318 33360 25374 33416
rect 24674 26832 24730 26888
rect 24674 25200 24730 25256
rect 25410 31728 25466 31784
rect 25318 30912 25374 30968
rect 24950 30096 25006 30152
rect 24950 29280 25006 29336
rect 24858 24384 24914 24440
rect 24766 21936 24822 21992
rect 24858 21120 24914 21176
rect 25686 26968 25742 27024
rect 24858 20304 24914 20360
rect 24858 19488 24914 19544
rect 25134 18672 25190 18728
rect 25134 17856 25190 17912
rect 24766 17040 24822 17096
rect 24674 16224 24730 16280
rect 25502 15428 25558 15464
rect 25502 15408 25504 15428
rect 25504 15408 25556 15428
rect 25556 15408 25558 15428
rect 25134 14592 25190 14648
rect 24766 13776 24822 13832
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22834 3984 22890 4040
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 25502 12960 25558 13016
rect 24766 11328 24822 11384
rect 24766 10376 24822 10432
rect 23386 4800 23442 4856
rect 23754 3440 23810 3496
rect 24950 9696 25006 9752
rect 25134 12144 25190 12200
rect 25134 8880 25190 8936
rect 25134 8064 25190 8120
rect 24766 7248 24822 7304
rect 24858 6432 24914 6488
rect 24766 5616 24822 5672
rect 25042 1536 25098 1592
rect 24950 720 25006 776
<< metal3 >>
rect 24485 56266 24551 56269
rect 26200 56266 27000 56296
rect 24485 56264 27000 56266
rect 24485 56208 24490 56264
rect 24546 56208 27000 56264
rect 24485 56206 27000 56208
rect 24485 56203 24551 56206
rect 26200 56176 27000 56206
rect 0 55450 800 55480
rect 3969 55450 4035 55453
rect 0 55448 4035 55450
rect 0 55392 3974 55448
rect 4030 55392 4035 55448
rect 0 55390 4035 55392
rect 0 55360 800 55390
rect 3969 55387 4035 55390
rect 24669 55450 24735 55453
rect 26200 55450 27000 55480
rect 24669 55448 27000 55450
rect 24669 55392 24674 55448
rect 24730 55392 27000 55448
rect 24669 55390 27000 55392
rect 24669 55387 24735 55390
rect 26200 55360 27000 55390
rect 24761 54634 24827 54637
rect 26200 54634 27000 54664
rect 24761 54632 27000 54634
rect 24761 54576 24766 54632
rect 24822 54576 27000 54632
rect 24761 54574 27000 54576
rect 24761 54571 24827 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 17033 53954 17099 53957
rect 17166 53954 17172 53956
rect 17033 53952 17172 53954
rect 17033 53896 17038 53952
rect 17094 53896 17172 53952
rect 17033 53894 17172 53896
rect 17033 53891 17099 53894
rect 17166 53892 17172 53894
rect 17236 53892 17242 53956
rect 21950 53892 21956 53956
rect 22020 53954 22026 53956
rect 22277 53954 22343 53957
rect 22020 53952 22343 53954
rect 22020 53896 22282 53952
rect 22338 53896 22343 53952
rect 22020 53894 22343 53896
rect 22020 53892 22026 53894
rect 22277 53891 22343 53894
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 25313 53818 25379 53821
rect 26200 53818 27000 53848
rect 25313 53816 27000 53818
rect 25313 53760 25318 53816
rect 25374 53760 27000 53816
rect 25313 53758 27000 53760
rect 25313 53755 25379 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 0 53002 800 53032
rect 2957 53002 3023 53005
rect 0 53000 3023 53002
rect 0 52944 2962 53000
rect 3018 52944 3023 53000
rect 0 52942 3023 52944
rect 0 52912 800 52942
rect 2957 52939 3023 52942
rect 25313 53002 25379 53005
rect 26200 53002 27000 53032
rect 25313 53000 27000 53002
rect 25313 52944 25318 53000
rect 25374 52944 27000 53000
rect 25313 52942 27000 52944
rect 25313 52939 25379 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 13997 52596 14063 52597
rect 13997 52592 14044 52596
rect 14108 52594 14114 52596
rect 23841 52594 23907 52597
rect 23974 52594 23980 52596
rect 13997 52536 14002 52592
rect 13997 52532 14044 52536
rect 14108 52534 14154 52594
rect 23841 52592 23980 52594
rect 23841 52536 23846 52592
rect 23902 52536 23980 52592
rect 23841 52534 23980 52536
rect 14108 52532 14114 52534
rect 13997 52531 14063 52532
rect 23841 52531 23907 52534
rect 23974 52532 23980 52534
rect 24044 52532 24050 52596
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 25313 52186 25379 52189
rect 26200 52186 27000 52216
rect 25313 52184 27000 52186
rect 25313 52128 25318 52184
rect 25374 52128 27000 52184
rect 25313 52126 27000 52128
rect 25313 52123 25379 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25313 51370 25379 51373
rect 26200 51370 27000 51400
rect 25313 51368 27000 51370
rect 25313 51312 25318 51368
rect 25374 51312 27000 51368
rect 25313 51310 27000 51312
rect 25313 51307 25379 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 0 50554 800 50584
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 25313 50554 25379 50557
rect 26200 50554 27000 50584
rect 0 50494 1778 50554
rect 0 50464 800 50494
rect 1718 50418 1778 50494
rect 25313 50552 27000 50554
rect 25313 50496 25318 50552
rect 25374 50496 27000 50552
rect 25313 50494 27000 50496
rect 25313 50491 25379 50494
rect 26200 50464 27000 50494
rect 3325 50418 3391 50421
rect 1718 50416 3391 50418
rect 1718 50360 3330 50416
rect 3386 50360 3391 50416
rect 1718 50358 3391 50360
rect 3325 50355 3391 50358
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25313 49738 25379 49741
rect 26200 49738 27000 49768
rect 25313 49736 27000 49738
rect 25313 49680 25318 49736
rect 25374 49680 27000 49736
rect 25313 49678 27000 49680
rect 25313 49675 25379 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25313 48922 25379 48925
rect 26200 48922 27000 48952
rect 25313 48920 27000 48922
rect 25313 48864 25318 48920
rect 25374 48864 27000 48920
rect 25313 48862 27000 48864
rect 25313 48859 25379 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 0 48106 800 48136
rect 4061 48106 4127 48109
rect 0 48104 4127 48106
rect 0 48048 4066 48104
rect 4122 48048 4127 48104
rect 0 48046 4127 48048
rect 0 48016 800 48046
rect 4061 48043 4127 48046
rect 25405 48106 25471 48109
rect 26200 48106 27000 48136
rect 25405 48104 27000 48106
rect 25405 48048 25410 48104
rect 25466 48048 27000 48104
rect 25405 48046 27000 48048
rect 25405 48043 25471 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 18229 47154 18295 47157
rect 19241 47156 19307 47157
rect 18822 47154 18828 47156
rect 18229 47152 18828 47154
rect 18229 47096 18234 47152
rect 18290 47096 18828 47152
rect 18229 47094 18828 47096
rect 18229 47091 18295 47094
rect 18822 47092 18828 47094
rect 18892 47092 18898 47156
rect 19190 47154 19196 47156
rect 19150 47094 19196 47154
rect 19260 47152 19307 47156
rect 19302 47096 19307 47152
rect 19190 47092 19196 47094
rect 19260 47092 19307 47096
rect 19241 47091 19307 47092
rect 19609 47018 19675 47021
rect 19926 47018 19932 47020
rect 19609 47016 19932 47018
rect 19609 46960 19614 47016
rect 19670 46960 19932 47016
rect 19609 46958 19932 46960
rect 19609 46955 19675 46958
rect 19926 46956 19932 46958
rect 19996 46956 20002 47020
rect 22686 46956 22692 47020
rect 22756 47018 22762 47020
rect 25037 47018 25103 47021
rect 22756 47016 25103 47018
rect 22756 46960 25042 47016
rect 25098 46960 25103 47016
rect 22756 46958 25103 46960
rect 22756 46956 22762 46958
rect 25037 46955 25103 46958
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25221 46474 25287 46477
rect 26200 46474 27000 46504
rect 25221 46472 27000 46474
rect 25221 46416 25226 46472
rect 25282 46416 27000 46472
rect 25221 46414 27000 46416
rect 25221 46411 25287 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 0 45658 800 45688
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 3969 45658 4035 45661
rect 0 45656 4035 45658
rect 0 45600 3974 45656
rect 4030 45600 4035 45656
rect 0 45598 4035 45600
rect 0 45568 800 45598
rect 3969 45595 4035 45598
rect 24485 45658 24551 45661
rect 26200 45658 27000 45688
rect 24485 45656 27000 45658
rect 24485 45600 24490 45656
rect 24546 45600 27000 45656
rect 24485 45598 27000 45600
rect 24485 45595 24551 45598
rect 26200 45568 27000 45598
rect 12249 45252 12315 45253
rect 12198 45188 12204 45252
rect 12268 45250 12315 45252
rect 12268 45248 12360 45250
rect 12310 45192 12360 45248
rect 12268 45190 12360 45192
rect 12268 45188 12315 45190
rect 12249 45187 12315 45188
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25313 44842 25379 44845
rect 26200 44842 27000 44872
rect 25313 44840 27000 44842
rect 25313 44784 25318 44840
rect 25374 44784 27000 44840
rect 25313 44782 27000 44784
rect 25313 44779 25379 44782
rect 26200 44752 27000 44782
rect 10501 44708 10567 44709
rect 10501 44706 10548 44708
rect 10456 44704 10548 44706
rect 10456 44648 10506 44704
rect 10456 44646 10548 44648
rect 10501 44644 10548 44646
rect 10612 44644 10618 44708
rect 11094 44644 11100 44708
rect 11164 44706 11170 44708
rect 11237 44706 11303 44709
rect 21817 44708 21883 44709
rect 11164 44704 11303 44706
rect 11164 44648 11242 44704
rect 11298 44648 11303 44704
rect 11164 44646 11303 44648
rect 11164 44644 11170 44646
rect 10501 44643 10567 44644
rect 11237 44643 11303 44646
rect 21766 44644 21772 44708
rect 21836 44706 21883 44708
rect 21836 44704 21928 44706
rect 21878 44648 21928 44704
rect 21836 44646 21928 44648
rect 21836 44644 21883 44646
rect 21817 44643 21883 44644
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 23606 44372 23612 44436
rect 23676 44434 23682 44436
rect 24761 44434 24827 44437
rect 23676 44432 24827 44434
rect 23676 44376 24766 44432
rect 24822 44376 24827 44432
rect 23676 44374 24827 44376
rect 23676 44372 23682 44374
rect 24761 44371 24827 44374
rect 9213 44298 9279 44301
rect 11605 44300 11671 44301
rect 9438 44298 9444 44300
rect 9213 44296 9444 44298
rect 9213 44240 9218 44296
rect 9274 44240 9444 44296
rect 9213 44238 9444 44240
rect 9213 44235 9279 44238
rect 9438 44236 9444 44238
rect 9508 44236 9514 44300
rect 11605 44298 11652 44300
rect 11560 44296 11652 44298
rect 11560 44240 11610 44296
rect 11560 44238 11652 44240
rect 11605 44236 11652 44238
rect 11716 44236 11722 44300
rect 23422 44236 23428 44300
rect 23492 44298 23498 44300
rect 24761 44298 24827 44301
rect 23492 44296 24827 44298
rect 23492 44240 24766 44296
rect 24822 44240 24827 44296
rect 23492 44238 24827 44240
rect 23492 44236 23498 44238
rect 11605 44235 11671 44236
rect 24761 44235 24827 44238
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24485 44026 24551 44029
rect 26200 44026 27000 44056
rect 24485 44024 27000 44026
rect 24485 43968 24490 44024
rect 24546 43968 27000 44024
rect 24485 43966 27000 43968
rect 24485 43963 24551 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 0 43210 800 43240
rect 1301 43210 1367 43213
rect 0 43208 1367 43210
rect 0 43152 1306 43208
rect 1362 43152 1367 43208
rect 0 43150 1367 43152
rect 0 43120 800 43150
rect 1301 43147 1367 43150
rect 24669 43210 24735 43213
rect 26200 43210 27000 43240
rect 24669 43208 27000 43210
rect 24669 43152 24674 43208
rect 24730 43152 27000 43208
rect 24669 43150 27000 43152
rect 24669 43147 24735 43150
rect 26200 43120 27000 43150
rect 20294 43012 20300 43076
rect 20364 43074 20370 43076
rect 21357 43074 21423 43077
rect 20364 43072 21423 43074
rect 20364 43016 21362 43072
rect 21418 43016 21423 43072
rect 20364 43014 21423 43016
rect 20364 43012 20370 43014
rect 21357 43011 21423 43014
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 24485 42394 24551 42397
rect 26200 42394 27000 42424
rect 24485 42392 27000 42394
rect 24485 42336 24490 42392
rect 24546 42336 27000 42392
rect 24485 42334 27000 42336
rect 24485 42331 24551 42334
rect 26200 42304 27000 42334
rect 6361 42258 6427 42261
rect 10174 42258 10180 42260
rect 6361 42256 10180 42258
rect 6361 42200 6366 42256
rect 6422 42200 10180 42256
rect 6361 42198 10180 42200
rect 6361 42195 6427 42198
rect 10174 42196 10180 42198
rect 10244 42196 10250 42260
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 22185 41578 22251 41581
rect 26200 41578 27000 41608
rect 22185 41576 27000 41578
rect 22185 41520 22190 41576
rect 22246 41520 27000 41576
rect 22185 41518 27000 41520
rect 22185 41515 22251 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 13445 41170 13511 41173
rect 19977 41170 20043 41173
rect 21173 41170 21239 41173
rect 13445 41168 21239 41170
rect 13445 41112 13450 41168
rect 13506 41112 19982 41168
rect 20038 41112 21178 41168
rect 21234 41112 21239 41168
rect 13445 41110 21239 41112
rect 13445 41107 13511 41110
rect 19977 41107 20043 41110
rect 21173 41107 21239 41110
rect 22461 41170 22527 41173
rect 22686 41170 22692 41172
rect 22461 41168 22692 41170
rect 22461 41112 22466 41168
rect 22522 41112 22692 41168
rect 22461 41110 22692 41112
rect 22461 41107 22527 41110
rect 22686 41108 22692 41110
rect 22756 41170 22762 41172
rect 22829 41170 22895 41173
rect 22756 41168 22895 41170
rect 22756 41112 22834 41168
rect 22890 41112 22895 41168
rect 22756 41110 22895 41112
rect 22756 41108 22762 41110
rect 22829 41107 22895 41110
rect 2946 40832 3262 40833
rect 0 40762 800 40792
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 1301 40762 1367 40765
rect 0 40760 1367 40762
rect 0 40704 1306 40760
rect 1362 40704 1367 40760
rect 0 40702 1367 40704
rect 0 40672 800 40702
rect 1301 40699 1367 40702
rect 13997 40762 14063 40765
rect 17401 40762 17467 40765
rect 17718 40762 17724 40764
rect 13997 40760 17724 40762
rect 13997 40704 14002 40760
rect 14058 40704 17406 40760
rect 17462 40704 17724 40760
rect 13997 40702 17724 40704
rect 13997 40699 14063 40702
rect 17401 40699 17467 40702
rect 17718 40700 17724 40702
rect 17788 40700 17794 40764
rect 24853 40762 24919 40765
rect 26200 40762 27000 40792
rect 24853 40760 27000 40762
rect 24853 40704 24858 40760
rect 24914 40704 27000 40760
rect 24853 40702 27000 40704
rect 24853 40699 24919 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 19977 40082 20043 40085
rect 20662 40082 20668 40084
rect 19977 40080 20668 40082
rect 19977 40024 19982 40080
rect 20038 40024 20668 40080
rect 19977 40022 20668 40024
rect 19977 40019 20043 40022
rect 20662 40020 20668 40022
rect 20732 40020 20738 40084
rect 22318 40020 22324 40084
rect 22388 40082 22394 40084
rect 22461 40082 22527 40085
rect 22388 40080 22527 40082
rect 22388 40024 22466 40080
rect 22522 40024 22527 40080
rect 22388 40022 22527 40024
rect 22388 40020 22394 40022
rect 22461 40019 22527 40022
rect 25405 39946 25471 39949
rect 26200 39946 27000 39976
rect 25405 39944 27000 39946
rect 25405 39888 25410 39944
rect 25466 39888 27000 39944
rect 25405 39886 27000 39888
rect 25405 39883 25471 39886
rect 26200 39856 27000 39886
rect 18822 39748 18828 39812
rect 18892 39810 18898 39812
rect 20253 39810 20319 39813
rect 18892 39808 20319 39810
rect 18892 39752 20258 39808
rect 20314 39752 20319 39808
rect 18892 39750 20319 39752
rect 18892 39748 18898 39750
rect 20253 39747 20319 39750
rect 21449 39810 21515 39813
rect 21909 39810 21975 39813
rect 22553 39810 22619 39813
rect 21449 39808 22619 39810
rect 21449 39752 21454 39808
rect 21510 39752 21914 39808
rect 21970 39752 22558 39808
rect 22614 39752 22619 39808
rect 21449 39750 22619 39752
rect 21449 39747 21515 39750
rect 21909 39747 21975 39750
rect 22553 39747 22619 39750
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 10133 39538 10199 39541
rect 12893 39538 12959 39541
rect 15837 39538 15903 39541
rect 10133 39536 15903 39538
rect 10133 39480 10138 39536
rect 10194 39480 12898 39536
rect 12954 39480 15842 39536
rect 15898 39480 15903 39536
rect 10133 39478 15903 39480
rect 10133 39475 10199 39478
rect 12893 39475 12959 39478
rect 15837 39475 15903 39478
rect 21582 39476 21588 39540
rect 21652 39538 21658 39540
rect 23422 39538 23428 39540
rect 21652 39478 23428 39538
rect 21652 39476 21658 39478
rect 23422 39476 23428 39478
rect 23492 39476 23498 39540
rect 10961 39402 11027 39405
rect 12985 39402 13051 39405
rect 10961 39400 13051 39402
rect 10961 39344 10966 39400
rect 11022 39344 12990 39400
rect 13046 39344 13051 39400
rect 10961 39342 13051 39344
rect 10961 39339 11027 39342
rect 12985 39339 13051 39342
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 10542 39068 10548 39132
rect 10612 39130 10618 39132
rect 16665 39130 16731 39133
rect 10612 39128 16731 39130
rect 10612 39072 16670 39128
rect 16726 39072 16731 39128
rect 10612 39070 16731 39072
rect 10612 39068 10618 39070
rect 16665 39067 16731 39070
rect 21817 39130 21883 39133
rect 26200 39130 27000 39160
rect 21817 39128 27000 39130
rect 21817 39072 21822 39128
rect 21878 39072 27000 39128
rect 21817 39070 27000 39072
rect 21817 39067 21883 39070
rect 26200 39040 27000 39070
rect 12433 38994 12499 38997
rect 13445 38994 13511 38997
rect 13670 38994 13676 38996
rect 12433 38992 13676 38994
rect 12433 38936 12438 38992
rect 12494 38936 13450 38992
rect 13506 38936 13676 38992
rect 12433 38934 13676 38936
rect 12433 38931 12499 38934
rect 13445 38931 13511 38934
rect 13670 38932 13676 38934
rect 13740 38932 13746 38996
rect 12341 38858 12407 38861
rect 15377 38858 15443 38861
rect 12341 38856 15443 38858
rect 12341 38800 12346 38856
rect 12402 38800 15382 38856
rect 15438 38800 15443 38856
rect 12341 38798 15443 38800
rect 12341 38795 12407 38798
rect 15377 38795 15443 38798
rect 15510 38796 15516 38860
rect 15580 38858 15586 38860
rect 15653 38858 15719 38861
rect 15580 38856 15719 38858
rect 15580 38800 15658 38856
rect 15714 38800 15719 38856
rect 15580 38798 15719 38800
rect 15580 38796 15586 38798
rect 15653 38795 15719 38798
rect 22461 38722 22527 38725
rect 22050 38720 22527 38722
rect 22050 38664 22466 38720
rect 22522 38664 22527 38720
rect 22050 38662 22527 38664
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 17677 38586 17743 38589
rect 22050 38586 22110 38662
rect 22461 38659 22527 38662
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 17677 38584 22110 38586
rect 17677 38528 17682 38584
rect 17738 38528 22110 38584
rect 17677 38526 22110 38528
rect 17677 38523 17743 38526
rect 12249 38452 12315 38453
rect 12198 38450 12204 38452
rect 12158 38390 12204 38450
rect 12268 38448 12315 38452
rect 12310 38392 12315 38448
rect 12198 38388 12204 38390
rect 12268 38388 12315 38392
rect 12249 38387 12315 38388
rect 15377 38450 15443 38453
rect 21582 38450 21588 38452
rect 15377 38448 21588 38450
rect 15377 38392 15382 38448
rect 15438 38392 21588 38448
rect 15377 38390 21588 38392
rect 15377 38387 15443 38390
rect 21582 38388 21588 38390
rect 21652 38388 21658 38452
rect 23289 38450 23355 38453
rect 23606 38450 23612 38452
rect 23289 38448 23612 38450
rect 23289 38392 23294 38448
rect 23350 38392 23612 38448
rect 23289 38390 23612 38392
rect 23289 38387 23355 38390
rect 23606 38388 23612 38390
rect 23676 38388 23682 38452
rect 0 38314 800 38344
rect 1301 38314 1367 38317
rect 0 38312 1367 38314
rect 0 38256 1306 38312
rect 1362 38256 1367 38312
rect 0 38254 1367 38256
rect 0 38224 800 38254
rect 1301 38251 1367 38254
rect 22185 38314 22251 38317
rect 26200 38314 27000 38344
rect 22185 38312 27000 38314
rect 22185 38256 22190 38312
rect 22246 38256 27000 38312
rect 22185 38254 27000 38256
rect 22185 38251 22251 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 22185 38042 22251 38045
rect 22737 38042 22803 38045
rect 23974 38042 23980 38044
rect 22185 38040 23980 38042
rect 22185 37984 22190 38040
rect 22246 37984 22742 38040
rect 22798 37984 23980 38040
rect 22185 37982 23980 37984
rect 22185 37979 22251 37982
rect 22737 37979 22803 37982
rect 23974 37980 23980 37982
rect 24044 37980 24050 38044
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 24485 37498 24551 37501
rect 26200 37498 27000 37528
rect 24485 37496 27000 37498
rect 24485 37440 24490 37496
rect 24546 37440 27000 37496
rect 24485 37438 27000 37440
rect 24485 37435 24551 37438
rect 26200 37408 27000 37438
rect 14774 37300 14780 37364
rect 14844 37362 14850 37364
rect 20621 37362 20687 37365
rect 14844 37360 20687 37362
rect 14844 37304 20626 37360
rect 20682 37304 20687 37360
rect 14844 37302 20687 37304
rect 14844 37300 14850 37302
rect 20621 37299 20687 37302
rect 16389 37090 16455 37093
rect 10366 37088 16455 37090
rect 10366 37032 16394 37088
rect 16450 37032 16455 37088
rect 10366 37030 16455 37032
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 9397 36684 9463 36685
rect 9397 36682 9444 36684
rect 9356 36680 9444 36682
rect 9508 36682 9514 36684
rect 10366 36682 10426 37030
rect 16389 37027 16455 37030
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 22185 36954 22251 36957
rect 22318 36954 22324 36956
rect 22185 36952 22324 36954
rect 22185 36896 22190 36952
rect 22246 36896 22324 36952
rect 22185 36894 22324 36896
rect 22185 36891 22251 36894
rect 22318 36892 22324 36894
rect 22388 36892 22394 36956
rect 9356 36624 9402 36680
rect 9356 36622 9444 36624
rect 9397 36620 9444 36622
rect 9508 36622 10426 36682
rect 22185 36682 22251 36685
rect 26200 36682 27000 36712
rect 22185 36680 27000 36682
rect 22185 36624 22190 36680
rect 22246 36624 27000 36680
rect 22185 36622 27000 36624
rect 9508 36620 9514 36622
rect 9397 36619 9463 36620
rect 22185 36619 22251 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 22277 36138 22343 36141
rect 22737 36138 22803 36141
rect 22277 36136 22803 36138
rect 22277 36080 22282 36136
rect 22338 36080 22742 36136
rect 22798 36080 22803 36136
rect 22277 36078 22803 36080
rect 22277 36075 22343 36078
rect 22737 36075 22803 36078
rect 7946 35936 8262 35937
rect 0 35866 800 35896
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 1577 35866 1643 35869
rect 0 35864 1643 35866
rect 0 35808 1582 35864
rect 1638 35808 1643 35864
rect 0 35806 1643 35808
rect 0 35776 800 35806
rect 1577 35803 1643 35806
rect 22369 35866 22435 35869
rect 26200 35866 27000 35896
rect 22369 35864 27000 35866
rect 22369 35808 22374 35864
rect 22430 35808 27000 35864
rect 22369 35806 27000 35808
rect 22369 35803 22435 35806
rect 26200 35776 27000 35806
rect 12709 35730 12775 35733
rect 14774 35730 14780 35732
rect 12709 35728 14780 35730
rect 12709 35672 12714 35728
rect 12770 35672 14780 35728
rect 12709 35670 14780 35672
rect 12709 35667 12775 35670
rect 14774 35668 14780 35670
rect 14844 35668 14850 35732
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 24761 35050 24827 35053
rect 26200 35050 27000 35080
rect 24761 35048 27000 35050
rect 24761 34992 24766 35048
rect 24822 34992 27000 35048
rect 24761 34990 27000 34992
rect 24761 34987 24827 34990
rect 26200 34960 27000 34990
rect 11053 34916 11119 34917
rect 11053 34914 11100 34916
rect 11008 34912 11100 34914
rect 11008 34856 11058 34912
rect 11008 34854 11100 34856
rect 11053 34852 11100 34854
rect 11164 34852 11170 34916
rect 11053 34851 11119 34852
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 10174 34716 10180 34780
rect 10244 34778 10250 34780
rect 11145 34778 11211 34781
rect 10244 34776 11211 34778
rect 10244 34720 11150 34776
rect 11206 34720 11211 34776
rect 10244 34718 11211 34720
rect 10244 34716 10250 34718
rect 11145 34715 11211 34718
rect 14958 34580 14964 34644
rect 15028 34642 15034 34644
rect 19425 34642 19491 34645
rect 15028 34640 19491 34642
rect 15028 34584 19430 34640
rect 19486 34584 19491 34640
rect 15028 34582 19491 34584
rect 15028 34580 15034 34582
rect 19425 34579 19491 34582
rect 20662 34580 20668 34644
rect 20732 34642 20738 34644
rect 22829 34642 22895 34645
rect 20732 34640 22895 34642
rect 20732 34584 22834 34640
rect 22890 34584 22895 34640
rect 20732 34582 22895 34584
rect 20732 34580 20738 34582
rect 22829 34579 22895 34582
rect 14038 34444 14044 34508
rect 14108 34506 14114 34508
rect 17493 34506 17559 34509
rect 14108 34504 17559 34506
rect 14108 34448 17498 34504
rect 17554 34448 17559 34504
rect 14108 34446 17559 34448
rect 14108 34444 14114 34446
rect 17493 34443 17559 34446
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 24853 34234 24919 34237
rect 26200 34234 27000 34264
rect 24853 34232 27000 34234
rect 24853 34176 24858 34232
rect 24914 34176 27000 34232
rect 24853 34174 27000 34176
rect 24853 34171 24919 34174
rect 26200 34144 27000 34174
rect 14181 34098 14247 34101
rect 14958 34098 14964 34100
rect 14181 34096 14964 34098
rect 14181 34040 14186 34096
rect 14242 34040 14964 34096
rect 14181 34038 14964 34040
rect 14181 34035 14247 34038
rect 14958 34036 14964 34038
rect 15028 34036 15034 34100
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 0 33418 800 33448
rect 1209 33418 1275 33421
rect 0 33416 1275 33418
rect 0 33360 1214 33416
rect 1270 33360 1275 33416
rect 0 33358 1275 33360
rect 0 33328 800 33358
rect 1209 33355 1275 33358
rect 12566 33356 12572 33420
rect 12636 33418 12642 33420
rect 13353 33418 13419 33421
rect 12636 33416 13419 33418
rect 12636 33360 13358 33416
rect 13414 33360 13419 33416
rect 12636 33358 13419 33360
rect 12636 33356 12642 33358
rect 13353 33355 13419 33358
rect 25313 33418 25379 33421
rect 26200 33418 27000 33448
rect 25313 33416 27000 33418
rect 25313 33360 25318 33416
rect 25374 33360 27000 33416
rect 25313 33358 27000 33360
rect 25313 33355 25379 33358
rect 26200 33328 27000 33358
rect 13486 33220 13492 33284
rect 13556 33282 13562 33284
rect 14089 33282 14155 33285
rect 13556 33280 14155 33282
rect 13556 33224 14094 33280
rect 14150 33224 14155 33280
rect 13556 33222 14155 33224
rect 13556 33220 13562 33222
rect 14089 33219 14155 33222
rect 17677 33282 17743 33285
rect 19190 33282 19196 33284
rect 17677 33280 19196 33282
rect 17677 33224 17682 33280
rect 17738 33224 19196 33280
rect 17677 33222 19196 33224
rect 17677 33219 17743 33222
rect 19190 33220 19196 33222
rect 19260 33220 19266 33284
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 24945 32602 25011 32605
rect 26200 32602 27000 32632
rect 24945 32600 27000 32602
rect 24945 32544 24950 32600
rect 25006 32544 27000 32600
rect 24945 32542 27000 32544
rect 24945 32539 25011 32542
rect 26200 32512 27000 32542
rect 11646 32268 11652 32332
rect 11716 32330 11722 32332
rect 13353 32330 13419 32333
rect 11716 32328 13419 32330
rect 11716 32272 13358 32328
rect 13414 32272 13419 32328
rect 11716 32270 13419 32272
rect 11716 32268 11722 32270
rect 13353 32267 13419 32270
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 21909 32060 21975 32061
rect 21909 32058 21956 32060
rect 21864 32056 21956 32058
rect 21864 32000 21914 32056
rect 21864 31998 21956 32000
rect 21909 31996 21956 31998
rect 22020 31996 22026 32060
rect 21909 31995 21975 31996
rect 25405 31786 25471 31789
rect 26200 31786 27000 31816
rect 25405 31784 27000 31786
rect 25405 31728 25410 31784
rect 25466 31728 27000 31784
rect 25405 31726 27000 31728
rect 25405 31723 25471 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 21173 31514 21239 31517
rect 21582 31514 21588 31516
rect 21173 31512 21588 31514
rect 21173 31456 21178 31512
rect 21234 31456 21588 31512
rect 21173 31454 21588 31456
rect 21173 31451 21239 31454
rect 21582 31452 21588 31454
rect 21652 31452 21658 31516
rect 16021 31378 16087 31381
rect 17534 31378 17540 31380
rect 16021 31376 17540 31378
rect 16021 31320 16026 31376
rect 16082 31320 17540 31376
rect 16021 31318 17540 31320
rect 16021 31315 16087 31318
rect 17534 31316 17540 31318
rect 17604 31316 17610 31380
rect 2946 31040 3262 31041
rect 0 30970 800 31000
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 2773 30970 2839 30973
rect 0 30968 2839 30970
rect 0 30912 2778 30968
rect 2834 30912 2839 30968
rect 0 30910 2839 30912
rect 0 30880 800 30910
rect 2773 30907 2839 30910
rect 25313 30970 25379 30973
rect 26200 30970 27000 31000
rect 25313 30968 27000 30970
rect 25313 30912 25318 30968
rect 25374 30912 27000 30968
rect 25313 30910 27000 30912
rect 25313 30907 25379 30910
rect 26200 30880 27000 30910
rect 19793 30698 19859 30701
rect 19926 30698 19932 30700
rect 19793 30696 19932 30698
rect 19793 30640 19798 30696
rect 19854 30640 19932 30696
rect 19793 30638 19932 30640
rect 19793 30635 19859 30638
rect 19926 30636 19932 30638
rect 19996 30636 20002 30700
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 10542 30364 10548 30428
rect 10612 30426 10618 30428
rect 12341 30426 12407 30429
rect 10612 30424 12407 30426
rect 10612 30368 12346 30424
rect 12402 30368 12407 30424
rect 10612 30366 12407 30368
rect 10612 30364 10618 30366
rect 12341 30363 12407 30366
rect 18965 30426 19031 30429
rect 20294 30426 20300 30428
rect 18965 30424 20300 30426
rect 18965 30368 18970 30424
rect 19026 30368 20300 30424
rect 18965 30366 20300 30368
rect 18965 30363 19031 30366
rect 20294 30364 20300 30366
rect 20364 30364 20370 30428
rect 17401 30154 17467 30157
rect 18638 30154 18644 30156
rect 17401 30152 18644 30154
rect 17401 30096 17406 30152
rect 17462 30096 18644 30152
rect 17401 30094 18644 30096
rect 17401 30091 17467 30094
rect 18638 30092 18644 30094
rect 18708 30092 18714 30156
rect 24945 30154 25011 30157
rect 26200 30154 27000 30184
rect 24945 30152 27000 30154
rect 24945 30096 24950 30152
rect 25006 30096 27000 30152
rect 24945 30094 27000 30096
rect 24945 30091 25011 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 12198 29276 12204 29340
rect 12268 29338 12274 29340
rect 12341 29338 12407 29341
rect 12268 29336 12407 29338
rect 12268 29280 12346 29336
rect 12402 29280 12407 29336
rect 12268 29278 12407 29280
rect 12268 29276 12274 29278
rect 12341 29275 12407 29278
rect 24945 29338 25011 29341
rect 26200 29338 27000 29368
rect 24945 29336 27000 29338
rect 24945 29280 24950 29336
rect 25006 29280 27000 29336
rect 24945 29278 27000 29280
rect 24945 29275 25011 29278
rect 26200 29248 27000 29278
rect 16757 29068 16823 29069
rect 16757 29066 16804 29068
rect 16712 29064 16804 29066
rect 16712 29008 16762 29064
rect 16712 29006 16804 29008
rect 16757 29004 16804 29006
rect 16868 29004 16874 29068
rect 16757 29003 16823 29004
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 0 28522 800 28552
rect 2865 28522 2931 28525
rect 0 28520 2931 28522
rect 0 28464 2870 28520
rect 2926 28464 2931 28520
rect 0 28462 2931 28464
rect 0 28432 800 28462
rect 2865 28459 2931 28462
rect 24301 28522 24367 28525
rect 26200 28522 27000 28552
rect 24301 28520 27000 28522
rect 24301 28464 24306 28520
rect 24362 28464 27000 28520
rect 24301 28462 27000 28464
rect 24301 28459 24367 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 19701 28250 19767 28253
rect 21766 28250 21772 28252
rect 19701 28248 21772 28250
rect 19701 28192 19706 28248
rect 19762 28192 21772 28248
rect 19701 28190 21772 28192
rect 19701 28187 19767 28190
rect 21766 28188 21772 28190
rect 21836 28188 21842 28252
rect 15653 28114 15719 28117
rect 16389 28116 16455 28117
rect 16389 28114 16436 28116
rect 15653 28112 16436 28114
rect 15653 28056 15658 28112
rect 15714 28056 16394 28112
rect 15653 28054 16436 28056
rect 15653 28051 15719 28054
rect 16389 28052 16436 28054
rect 16500 28052 16506 28116
rect 17718 28052 17724 28116
rect 17788 28114 17794 28116
rect 17861 28114 17927 28117
rect 17788 28112 17927 28114
rect 17788 28056 17866 28112
rect 17922 28056 17927 28112
rect 17788 28054 17927 28056
rect 17788 28052 17794 28054
rect 16389 28051 16455 28052
rect 17861 28051 17927 28054
rect 17534 27780 17540 27844
rect 17604 27842 17610 27844
rect 18873 27842 18939 27845
rect 17604 27840 18939 27842
rect 17604 27784 18878 27840
rect 18934 27784 18939 27840
rect 17604 27782 18939 27784
rect 17604 27780 17610 27782
rect 18873 27779 18939 27782
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 16849 27706 16915 27709
rect 17166 27706 17172 27708
rect 16849 27704 17172 27706
rect 16849 27648 16854 27704
rect 16910 27648 17172 27704
rect 16849 27646 17172 27648
rect 16849 27643 16915 27646
rect 17166 27644 17172 27646
rect 17236 27644 17242 27708
rect 26200 27706 27000 27736
rect 23430 27646 27000 27706
rect 23289 27570 23355 27573
rect 23430 27570 23490 27646
rect 26200 27616 27000 27646
rect 23289 27568 23490 27570
rect 23289 27512 23294 27568
rect 23350 27512 23490 27568
rect 23289 27510 23490 27512
rect 23289 27507 23355 27510
rect 19701 27300 19767 27301
rect 19701 27298 19748 27300
rect 19656 27296 19748 27298
rect 19656 27240 19706 27296
rect 19656 27238 19748 27240
rect 19701 27236 19748 27238
rect 19812 27236 19818 27300
rect 19701 27235 19767 27236
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 17309 27026 17375 27029
rect 23381 27026 23447 27029
rect 25681 27026 25747 27029
rect 17309 27024 17602 27026
rect 17309 26968 17314 27024
rect 17370 26968 17602 27024
rect 17309 26966 17602 26968
rect 17309 26963 17375 26966
rect 9029 26756 9095 26757
rect 9029 26754 9076 26756
rect 8984 26752 9076 26754
rect 8984 26696 9034 26752
rect 8984 26694 9076 26696
rect 9029 26692 9076 26694
rect 9140 26692 9146 26756
rect 17542 26754 17602 26966
rect 23381 27024 25747 27026
rect 23381 26968 23386 27024
rect 23442 26968 25686 27024
rect 25742 26968 25747 27024
rect 23381 26966 25747 26968
rect 23381 26963 23447 26966
rect 25681 26963 25747 26966
rect 24669 26890 24735 26893
rect 26200 26890 27000 26920
rect 24669 26888 27000 26890
rect 24669 26832 24674 26888
rect 24730 26832 27000 26888
rect 24669 26830 27000 26832
rect 24669 26827 24735 26830
rect 26200 26800 27000 26830
rect 17677 26754 17743 26757
rect 17542 26752 17743 26754
rect 17542 26696 17682 26752
rect 17738 26696 17743 26752
rect 17542 26694 17743 26696
rect 9029 26691 9095 26692
rect 17677 26691 17743 26694
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 15193 26618 15259 26621
rect 16389 26618 16455 26621
rect 15193 26616 16455 26618
rect 15193 26560 15198 26616
rect 15254 26560 16394 26616
rect 16450 26560 16455 26616
rect 15193 26558 16455 26560
rect 15193 26555 15259 26558
rect 16389 26555 16455 26558
rect 14917 26482 14983 26485
rect 17125 26482 17191 26485
rect 14917 26480 17191 26482
rect 14917 26424 14922 26480
rect 14978 26424 17130 26480
rect 17186 26424 17191 26480
rect 14917 26422 17191 26424
rect 14917 26419 14983 26422
rect 17125 26419 17191 26422
rect 4889 26346 4955 26349
rect 17769 26346 17835 26349
rect 4889 26344 17835 26346
rect 4889 26288 4894 26344
rect 4950 26288 17774 26344
rect 17830 26288 17835 26344
rect 4889 26286 17835 26288
rect 4889 26283 4955 26286
rect 17769 26283 17835 26286
rect 15694 26148 15700 26212
rect 15764 26210 15770 26212
rect 16757 26210 16823 26213
rect 15764 26208 16823 26210
rect 15764 26152 16762 26208
rect 16818 26152 16823 26208
rect 15764 26150 16823 26152
rect 15764 26148 15770 26150
rect 16757 26147 16823 26150
rect 7946 26144 8262 26145
rect 0 26074 800 26104
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 2773 26074 2839 26077
rect 0 26072 2839 26074
rect 0 26016 2778 26072
rect 2834 26016 2839 26072
rect 0 26014 2839 26016
rect 0 25984 800 26014
rect 2773 26011 2839 26014
rect 23197 26074 23263 26077
rect 26200 26074 27000 26104
rect 23197 26072 27000 26074
rect 23197 26016 23202 26072
rect 23258 26016 27000 26072
rect 23197 26014 27000 26016
rect 23197 26011 23263 26014
rect 26200 25984 27000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 24669 25258 24735 25261
rect 26200 25258 27000 25288
rect 24669 25256 27000 25258
rect 24669 25200 24674 25256
rect 24730 25200 27000 25256
rect 24669 25198 27000 25200
rect 24669 25195 24735 25198
rect 26200 25168 27000 25198
rect 10225 25122 10291 25125
rect 10542 25122 10548 25124
rect 10225 25120 10548 25122
rect 10225 25064 10230 25120
rect 10286 25064 10548 25120
rect 10225 25062 10548 25064
rect 10225 25059 10291 25062
rect 10542 25060 10548 25062
rect 10612 25060 10618 25124
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24853 24442 24919 24445
rect 26200 24442 27000 24472
rect 24853 24440 27000 24442
rect 24853 24384 24858 24440
rect 24914 24384 27000 24440
rect 24853 24382 27000 24384
rect 24853 24379 24919 24382
rect 26200 24352 27000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 0 23626 800 23656
rect 2865 23626 2931 23629
rect 0 23624 2931 23626
rect 0 23568 2870 23624
rect 2926 23568 2931 23624
rect 0 23566 2931 23568
rect 0 23536 800 23566
rect 2865 23563 2931 23566
rect 23381 23626 23447 23629
rect 26200 23626 27000 23656
rect 23381 23624 27000 23626
rect 23381 23568 23386 23624
rect 23442 23568 27000 23624
rect 23381 23566 27000 23568
rect 23381 23563 23447 23566
rect 26200 23536 27000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 12525 23218 12591 23221
rect 13670 23218 13676 23220
rect 12525 23216 13676 23218
rect 12525 23160 12530 23216
rect 12586 23160 13676 23216
rect 12525 23158 13676 23160
rect 12525 23155 12591 23158
rect 13670 23156 13676 23158
rect 13740 23156 13746 23220
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 22829 22810 22895 22813
rect 26200 22810 27000 22840
rect 22829 22808 27000 22810
rect 22829 22752 22834 22808
rect 22890 22752 27000 22808
rect 22829 22750 27000 22752
rect 22829 22747 22895 22750
rect 26200 22720 27000 22750
rect 11513 22674 11579 22677
rect 12014 22674 12020 22676
rect 11513 22672 12020 22674
rect 11513 22616 11518 22672
rect 11574 22616 12020 22672
rect 11513 22614 12020 22616
rect 11513 22611 11579 22614
rect 12014 22612 12020 22614
rect 12084 22612 12090 22676
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 16798 22068 16804 22132
rect 16868 22130 16874 22132
rect 23422 22130 23428 22132
rect 16868 22070 23428 22130
rect 16868 22068 16874 22070
rect 23422 22068 23428 22070
rect 23492 22068 23498 22132
rect 24761 21994 24827 21997
rect 26200 21994 27000 22024
rect 24761 21992 27000 21994
rect 24761 21936 24766 21992
rect 24822 21936 27000 21992
rect 24761 21934 27000 21936
rect 24761 21931 24827 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 10133 21316 10199 21317
rect 13997 21316 14063 21317
rect 10133 21314 10180 21316
rect 10088 21312 10180 21314
rect 10088 21256 10138 21312
rect 10088 21254 10180 21256
rect 10133 21252 10180 21254
rect 10244 21252 10250 21316
rect 13997 21314 14044 21316
rect 13952 21312 14044 21314
rect 14108 21314 14114 21316
rect 14733 21314 14799 21317
rect 14108 21312 14799 21314
rect 13952 21256 14002 21312
rect 14108 21256 14738 21312
rect 14794 21256 14799 21312
rect 13952 21254 14044 21256
rect 13997 21252 14044 21254
rect 14108 21254 14799 21256
rect 14108 21252 14114 21254
rect 10133 21251 10199 21252
rect 13997 21251 14063 21252
rect 14733 21251 14799 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 1301 21178 1367 21181
rect 18781 21180 18847 21181
rect 18781 21178 18828 21180
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 18736 21176 18828 21178
rect 18736 21120 18786 21176
rect 18736 21118 18828 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 18781 21116 18828 21118
rect 18892 21116 18898 21180
rect 24853 21178 24919 21181
rect 26200 21178 27000 21208
rect 24853 21176 27000 21178
rect 24853 21120 24858 21176
rect 24914 21120 27000 21176
rect 24853 21118 27000 21120
rect 18781 21115 18847 21116
rect 24853 21115 24919 21118
rect 26200 21088 27000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 15009 20364 15075 20365
rect 14958 20300 14964 20364
rect 15028 20362 15075 20364
rect 15028 20360 15120 20362
rect 15070 20304 15120 20360
rect 15028 20302 15120 20304
rect 15028 20300 15075 20302
rect 15510 20300 15516 20364
rect 15580 20362 15586 20364
rect 15745 20362 15811 20365
rect 15580 20360 15811 20362
rect 15580 20304 15750 20360
rect 15806 20304 15811 20360
rect 15580 20302 15811 20304
rect 15580 20300 15586 20302
rect 15009 20299 15075 20300
rect 15745 20299 15811 20302
rect 24853 20362 24919 20365
rect 26200 20362 27000 20392
rect 24853 20360 27000 20362
rect 24853 20304 24858 20360
rect 24914 20304 27000 20360
rect 24853 20302 27000 20304
rect 24853 20299 24919 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 16481 19954 16547 19957
rect 19742 19954 19748 19956
rect 16481 19952 19748 19954
rect 16481 19896 16486 19952
rect 16542 19896 19748 19952
rect 16481 19894 19748 19896
rect 16481 19891 16547 19894
rect 19742 19892 19748 19894
rect 19812 19954 19818 19956
rect 22134 19954 22140 19956
rect 19812 19894 22140 19954
rect 19812 19892 19818 19894
rect 22134 19892 22140 19894
rect 22204 19892 22210 19956
rect 10501 19820 10567 19821
rect 10501 19818 10548 19820
rect 10456 19816 10548 19818
rect 10456 19760 10506 19816
rect 10456 19758 10548 19760
rect 10501 19756 10548 19758
rect 10612 19756 10618 19820
rect 10501 19755 10567 19756
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 24853 19546 24919 19549
rect 26200 19546 27000 19576
rect 24853 19544 27000 19546
rect 24853 19488 24858 19544
rect 24914 19488 27000 19544
rect 24853 19486 27000 19488
rect 24853 19483 24919 19486
rect 26200 19456 27000 19486
rect 18597 19410 18663 19413
rect 18822 19410 18828 19412
rect 18597 19408 18828 19410
rect 18597 19352 18602 19408
rect 18658 19352 18828 19408
rect 18597 19350 18828 19352
rect 18597 19347 18663 19350
rect 18822 19348 18828 19350
rect 18892 19348 18898 19412
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 18689 18868 18755 18869
rect 18638 18804 18644 18868
rect 18708 18866 18755 18868
rect 18708 18864 18800 18866
rect 18750 18808 18800 18864
rect 18708 18806 18800 18808
rect 18708 18804 18755 18806
rect 18689 18803 18755 18804
rect 0 18730 800 18760
rect 1301 18730 1367 18733
rect 0 18728 1367 18730
rect 0 18672 1306 18728
rect 1362 18672 1367 18728
rect 0 18670 1367 18672
rect 0 18640 800 18670
rect 1301 18667 1367 18670
rect 25129 18730 25195 18733
rect 26200 18730 27000 18760
rect 25129 18728 27000 18730
rect 25129 18672 25134 18728
rect 25190 18672 27000 18728
rect 25129 18670 27000 18672
rect 25129 18667 25195 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 14733 18460 14799 18461
rect 14733 18458 14780 18460
rect 14688 18456 14780 18458
rect 14688 18400 14738 18456
rect 14688 18398 14780 18400
rect 14733 18396 14780 18398
rect 14844 18396 14850 18460
rect 14733 18395 14799 18396
rect 18413 18050 18479 18053
rect 19926 18050 19932 18052
rect 18413 18048 19932 18050
rect 18413 17992 18418 18048
rect 18474 17992 19932 18048
rect 18413 17990 19932 17992
rect 18413 17987 18479 17990
rect 19926 17988 19932 17990
rect 19996 17988 20002 18052
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 25129 17914 25195 17917
rect 26200 17914 27000 17944
rect 25129 17912 27000 17914
rect 25129 17856 25134 17912
rect 25190 17856 27000 17912
rect 25129 17854 27000 17856
rect 25129 17851 25195 17854
rect 26200 17824 27000 17854
rect 13486 17580 13492 17644
rect 13556 17642 13562 17644
rect 13629 17642 13695 17645
rect 13556 17640 13695 17642
rect 13556 17584 13634 17640
rect 13690 17584 13695 17640
rect 13556 17582 13695 17584
rect 13556 17580 13562 17582
rect 13629 17579 13695 17582
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 10777 17370 10843 17373
rect 12433 17370 12499 17373
rect 10777 17368 12499 17370
rect 10777 17312 10782 17368
rect 10838 17312 12438 17368
rect 12494 17312 12499 17368
rect 10777 17310 12499 17312
rect 10777 17307 10843 17310
rect 12433 17307 12499 17310
rect 24761 17098 24827 17101
rect 26200 17098 27000 17128
rect 24761 17096 27000 17098
rect 24761 17040 24766 17096
rect 24822 17040 27000 17096
rect 24761 17038 27000 17040
rect 24761 17035 24827 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 16389 16828 16455 16829
rect 16389 16826 16436 16828
rect 16344 16824 16436 16826
rect 16344 16768 16394 16824
rect 16344 16766 16436 16768
rect 16389 16764 16436 16766
rect 16500 16764 16506 16828
rect 16389 16763 16455 16764
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 24669 16282 24735 16285
rect 26200 16282 27000 16312
rect 24669 16280 27000 16282
rect 24669 16224 24674 16280
rect 24730 16224 27000 16280
rect 24669 16222 27000 16224
rect 24669 16219 24735 16222
rect 26200 16192 27000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 25497 15466 25563 15469
rect 26200 15466 27000 15496
rect 25497 15464 27000 15466
rect 25497 15408 25502 15464
rect 25558 15408 27000 15464
rect 25497 15406 27000 15408
rect 25497 15403 25563 15406
rect 26200 15376 27000 15406
rect 15009 15330 15075 15333
rect 15694 15330 15700 15332
rect 15009 15328 15700 15330
rect 15009 15272 15014 15328
rect 15070 15272 15700 15328
rect 15009 15270 15700 15272
rect 15009 15267 15075 15270
rect 15694 15268 15700 15270
rect 15764 15268 15770 15332
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 17493 15196 17559 15197
rect 17493 15194 17540 15196
rect 17448 15192 17540 15194
rect 17448 15136 17498 15192
rect 17448 15134 17540 15136
rect 17493 15132 17540 15134
rect 17604 15132 17610 15196
rect 17493 15131 17559 15132
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 25129 14650 25195 14653
rect 26200 14650 27000 14680
rect 25129 14648 27000 14650
rect 25129 14592 25134 14648
rect 25190 14592 27000 14648
rect 25129 14590 27000 14592
rect 25129 14587 25195 14590
rect 26200 14560 27000 14590
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 0 13834 800 13864
rect 933 13834 999 13837
rect 0 13832 999 13834
rect 0 13776 938 13832
rect 994 13776 999 13832
rect 0 13774 999 13776
rect 0 13744 800 13774
rect 933 13771 999 13774
rect 24761 13834 24827 13837
rect 26200 13834 27000 13864
rect 24761 13832 27000 13834
rect 24761 13776 24766 13832
rect 24822 13776 27000 13832
rect 24761 13774 27000 13776
rect 24761 13771 24827 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 12566 13364 12572 13428
rect 12636 13426 12642 13428
rect 12893 13426 12959 13429
rect 12636 13424 12959 13426
rect 12636 13368 12898 13424
rect 12954 13368 12959 13424
rect 12636 13366 12959 13368
rect 12636 13364 12642 13366
rect 12893 13363 12959 13366
rect 16021 13290 16087 13293
rect 17493 13290 17559 13293
rect 16021 13288 17559 13290
rect 16021 13232 16026 13288
rect 16082 13232 17498 13288
rect 17554 13232 17559 13288
rect 16021 13230 17559 13232
rect 16021 13227 16087 13230
rect 17493 13227 17559 13230
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 12014 12956 12020 13020
rect 12084 13018 12090 13020
rect 12157 13018 12223 13021
rect 12084 13016 12223 13018
rect 12084 12960 12162 13016
rect 12218 12960 12223 13016
rect 12084 12958 12223 12960
rect 12084 12956 12090 12958
rect 12157 12955 12223 12958
rect 25497 13018 25563 13021
rect 26200 13018 27000 13048
rect 25497 13016 27000 13018
rect 25497 12960 25502 13016
rect 25558 12960 27000 13016
rect 25497 12958 27000 12960
rect 25497 12955 25563 12958
rect 26200 12928 27000 12958
rect 20345 12882 20411 12885
rect 22318 12882 22324 12884
rect 20345 12880 22324 12882
rect 20345 12824 20350 12880
rect 20406 12824 22324 12880
rect 20345 12822 22324 12824
rect 20345 12819 20411 12822
rect 22318 12820 22324 12822
rect 22388 12820 22394 12884
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 25129 12202 25195 12205
rect 26200 12202 27000 12232
rect 25129 12200 27000 12202
rect 25129 12144 25134 12200
rect 25190 12144 27000 12200
rect 25129 12142 27000 12144
rect 25129 12139 25195 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 22093 11932 22159 11933
rect 22093 11930 22140 11932
rect 22048 11928 22140 11930
rect 22048 11872 22098 11928
rect 22048 11870 22140 11872
rect 22093 11868 22140 11870
rect 22204 11868 22210 11932
rect 22093 11867 22159 11868
rect 13537 11658 13603 11661
rect 13537 11656 13738 11658
rect 13537 11600 13542 11656
rect 13598 11600 13738 11656
rect 13537 11598 13738 11600
rect 13537 11595 13603 11598
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 13678 11389 13738 11598
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 2773 11386 2839 11389
rect 0 11384 2839 11386
rect 0 11328 2778 11384
rect 2834 11328 2839 11384
rect 0 11326 2839 11328
rect 13678 11384 13787 11389
rect 13678 11328 13726 11384
rect 13782 11328 13787 11384
rect 13678 11326 13787 11328
rect 0 11296 800 11326
rect 2773 11323 2839 11326
rect 13721 11323 13787 11326
rect 24761 11386 24827 11389
rect 26200 11386 27000 11416
rect 24761 11384 27000 11386
rect 24761 11328 24766 11384
rect 24822 11328 27000 11384
rect 24761 11326 27000 11328
rect 24761 11323 24827 11326
rect 26200 11296 27000 11326
rect 10041 10978 10107 10981
rect 14958 10978 14964 10980
rect 10041 10976 14964 10978
rect 10041 10920 10046 10976
rect 10102 10920 14964 10976
rect 10041 10918 14964 10920
rect 10041 10915 10107 10918
rect 14958 10916 14964 10918
rect 15028 10916 15034 10980
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 26200 10570 27000 10600
rect 24902 10510 27000 10570
rect 24761 10434 24827 10437
rect 24902 10434 24962 10510
rect 26200 10480 27000 10510
rect 24761 10432 24962 10434
rect 24761 10376 24766 10432
rect 24822 10376 24962 10432
rect 24761 10374 24962 10376
rect 24761 10371 24827 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24945 9754 25011 9757
rect 26200 9754 27000 9784
rect 24945 9752 27000 9754
rect 24945 9696 24950 9752
rect 25006 9696 27000 9752
rect 24945 9694 27000 9696
rect 24945 9691 25011 9694
rect 26200 9664 27000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 0 8938 800 8968
rect 2865 8938 2931 8941
rect 0 8936 2931 8938
rect 0 8880 2870 8936
rect 2926 8880 2931 8936
rect 0 8878 2931 8880
rect 0 8848 800 8878
rect 2865 8875 2931 8878
rect 25129 8938 25195 8941
rect 26200 8938 27000 8968
rect 25129 8936 27000 8938
rect 25129 8880 25134 8936
rect 25190 8880 27000 8936
rect 25129 8878 27000 8880
rect 25129 8875 25195 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 9213 7986 9279 7989
rect 14038 7986 14044 7988
rect 9213 7984 14044 7986
rect 9213 7928 9218 7984
rect 9274 7928 14044 7984
rect 9213 7926 14044 7928
rect 9213 7923 9279 7926
rect 14038 7924 14044 7926
rect 14108 7924 14114 7988
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 24761 7306 24827 7309
rect 26200 7306 27000 7336
rect 24761 7304 27000 7306
rect 24761 7248 24766 7304
rect 24822 7248 27000 7304
rect 24761 7246 27000 7248
rect 24761 7243 24827 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3141 6490 3207 6493
rect 0 6488 3207 6490
rect 0 6432 3146 6488
rect 3202 6432 3207 6488
rect 0 6430 3207 6432
rect 0 6400 800 6430
rect 3141 6427 3207 6430
rect 24853 6490 24919 6493
rect 26200 6490 27000 6520
rect 24853 6488 27000 6490
rect 24853 6432 24858 6488
rect 24914 6432 27000 6488
rect 24853 6430 27000 6432
rect 24853 6427 24919 6430
rect 26200 6400 27000 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 24761 5674 24827 5677
rect 26200 5674 27000 5704
rect 24761 5672 27000 5674
rect 24761 5616 24766 5672
rect 24822 5616 27000 5672
rect 24761 5614 27000 5616
rect 24761 5611 24827 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23381 4858 23447 4861
rect 26200 4858 27000 4888
rect 23381 4856 27000 4858
rect 23381 4800 23386 4856
rect 23442 4800 27000 4856
rect 23381 4798 27000 4800
rect 23381 4795 23447 4798
rect 26200 4768 27000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 0 4042 800 4072
rect 4061 4042 4127 4045
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 0 3952 800 3982
rect 4061 3979 4127 3982
rect 18781 4044 18847 4045
rect 18781 4040 18828 4044
rect 18892 4042 18898 4044
rect 22185 4042 22251 4045
rect 22318 4042 22324 4044
rect 18781 3984 18786 4040
rect 18781 3980 18828 3984
rect 18892 3982 18938 4042
rect 22185 4040 22324 4042
rect 22185 3984 22190 4040
rect 22246 3984 22324 4040
rect 22185 3982 22324 3984
rect 18892 3980 18898 3982
rect 18781 3979 18847 3980
rect 22185 3979 22251 3982
rect 22318 3980 22324 3982
rect 22388 3980 22394 4044
rect 22829 4042 22895 4045
rect 26200 4042 27000 4072
rect 22829 4040 27000 4042
rect 22829 3984 22834 4040
rect 22890 3984 27000 4040
rect 22829 3982 27000 3984
rect 22829 3979 22895 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 5257 3634 5323 3637
rect 10174 3634 10180 3636
rect 5257 3632 10180 3634
rect 5257 3576 5262 3632
rect 5318 3576 10180 3632
rect 5257 3574 10180 3576
rect 5257 3571 5323 3574
rect 10174 3572 10180 3574
rect 10244 3572 10250 3636
rect 3325 3498 3391 3501
rect 10542 3498 10548 3500
rect 3325 3496 10548 3498
rect 3325 3440 3330 3496
rect 3386 3440 10548 3496
rect 3325 3438 10548 3440
rect 3325 3435 3391 3438
rect 10542 3436 10548 3438
rect 10612 3436 10618 3500
rect 23422 3436 23428 3500
rect 23492 3498 23498 3500
rect 23749 3498 23815 3501
rect 23492 3496 23815 3498
rect 23492 3440 23754 3496
rect 23810 3440 23815 3496
rect 23492 3438 23815 3440
rect 23492 3436 23498 3438
rect 23749 3435 23815 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 8385 3226 8451 3229
rect 12198 3226 12204 3228
rect 8385 3224 12204 3226
rect 8385 3168 8390 3224
rect 8446 3168 12204 3224
rect 8385 3166 12204 3168
rect 8385 3163 8451 3166
rect 12198 3164 12204 3166
rect 12268 3164 12274 3228
rect 22093 3226 22159 3229
rect 26200 3226 27000 3256
rect 22093 3224 27000 3226
rect 22093 3168 22098 3224
rect 22154 3168 27000 3224
rect 22093 3166 27000 3168
rect 22093 3163 22159 3166
rect 26200 3136 27000 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 4061 2682 4127 2685
rect 9070 2682 9076 2684
rect 4061 2680 9076 2682
rect 4061 2624 4066 2680
rect 4122 2624 9076 2680
rect 4061 2622 9076 2624
rect 4061 2619 4127 2622
rect 9070 2620 9076 2622
rect 9140 2620 9146 2684
rect 21817 2410 21883 2413
rect 26200 2410 27000 2440
rect 21817 2408 27000 2410
rect 21817 2352 21822 2408
rect 21878 2352 27000 2408
rect 21817 2350 27000 2352
rect 21817 2347 21883 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1594 800 1624
rect 1393 1594 1459 1597
rect 0 1592 1459 1594
rect 0 1536 1398 1592
rect 1454 1536 1459 1592
rect 0 1534 1459 1536
rect 0 1504 800 1534
rect 1393 1531 1459 1534
rect 25037 1594 25103 1597
rect 26200 1594 27000 1624
rect 25037 1592 27000 1594
rect 25037 1536 25042 1592
rect 25098 1536 27000 1592
rect 25037 1534 27000 1536
rect 25037 1531 25103 1534
rect 26200 1504 27000 1534
rect 24945 778 25011 781
rect 26200 778 27000 808
rect 24945 776 27000 778
rect 24945 720 24950 776
rect 25006 720 27000 776
rect 24945 718 27000 720
rect 24945 715 25011 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 17172 53892 17236 53956
rect 21956 53892 22020 53956
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 14044 52592 14108 52596
rect 14044 52536 14058 52592
rect 14058 52536 14108 52592
rect 14044 52532 14108 52536
rect 23980 52532 24044 52596
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 18828 47092 18892 47156
rect 19196 47152 19260 47156
rect 19196 47096 19246 47152
rect 19246 47096 19260 47152
rect 19196 47092 19260 47096
rect 19932 46956 19996 47020
rect 22692 46956 22756 47020
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 12204 45248 12268 45252
rect 12204 45192 12254 45248
rect 12254 45192 12268 45248
rect 12204 45188 12268 45192
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 10548 44704 10612 44708
rect 10548 44648 10562 44704
rect 10562 44648 10612 44704
rect 10548 44644 10612 44648
rect 11100 44644 11164 44708
rect 21772 44704 21836 44708
rect 21772 44648 21822 44704
rect 21822 44648 21836 44704
rect 21772 44644 21836 44648
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 23612 44372 23676 44436
rect 9444 44236 9508 44300
rect 11652 44296 11716 44300
rect 11652 44240 11666 44296
rect 11666 44240 11716 44296
rect 11652 44236 11716 44240
rect 23428 44236 23492 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 20300 43012 20364 43076
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 10180 42196 10244 42260
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 22692 41108 22756 41172
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 17724 40700 17788 40764
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 20668 40020 20732 40084
rect 22324 40020 22388 40084
rect 18828 39748 18892 39812
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 21588 39476 21652 39540
rect 23428 39476 23492 39540
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 10548 39068 10612 39132
rect 13676 38932 13740 38996
rect 15516 38796 15580 38860
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 12204 38448 12268 38452
rect 12204 38392 12254 38448
rect 12254 38392 12268 38448
rect 12204 38388 12268 38392
rect 21588 38388 21652 38452
rect 23612 38388 23676 38452
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 23980 37980 24044 38044
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 14780 37300 14844 37364
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 9444 36680 9508 36684
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 22324 36892 22388 36956
rect 9444 36624 9458 36680
rect 9458 36624 9508 36680
rect 9444 36620 9508 36624
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 14780 35668 14844 35732
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 11100 34912 11164 34916
rect 11100 34856 11114 34912
rect 11114 34856 11164 34912
rect 11100 34852 11164 34856
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 10180 34716 10244 34780
rect 14964 34580 15028 34644
rect 20668 34580 20732 34644
rect 14044 34444 14108 34508
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 14964 34036 15028 34100
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 12572 33356 12636 33420
rect 13492 33220 13556 33284
rect 19196 33220 19260 33284
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 11652 32268 11716 32332
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 21956 32056 22020 32060
rect 21956 32000 21970 32056
rect 21970 32000 22020 32056
rect 21956 31996 22020 32000
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 21588 31452 21652 31516
rect 17540 31316 17604 31380
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 19932 30636 19996 30700
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 10548 30364 10612 30428
rect 20300 30364 20364 30428
rect 18644 30092 18708 30156
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 12204 29276 12268 29340
rect 16804 29064 16868 29068
rect 16804 29008 16818 29064
rect 16818 29008 16868 29064
rect 16804 29004 16868 29008
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 21772 28188 21836 28252
rect 16436 28112 16500 28116
rect 16436 28056 16450 28112
rect 16450 28056 16500 28112
rect 16436 28052 16500 28056
rect 17724 28052 17788 28116
rect 17540 27780 17604 27844
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 17172 27644 17236 27708
rect 19748 27296 19812 27300
rect 19748 27240 19762 27296
rect 19762 27240 19812 27296
rect 19748 27236 19812 27240
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 9076 26752 9140 26756
rect 9076 26696 9090 26752
rect 9090 26696 9140 26752
rect 9076 26692 9140 26696
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 15700 26148 15764 26212
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 10548 25060 10612 25124
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 13676 23156 13740 23220
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 12020 22612 12084 22676
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 16804 22068 16868 22132
rect 23428 22068 23492 22132
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 10180 21312 10244 21316
rect 10180 21256 10194 21312
rect 10194 21256 10244 21312
rect 10180 21252 10244 21256
rect 14044 21312 14108 21316
rect 14044 21256 14058 21312
rect 14058 21256 14108 21312
rect 14044 21252 14108 21256
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 18828 21176 18892 21180
rect 18828 21120 18842 21176
rect 18842 21120 18892 21176
rect 18828 21116 18892 21120
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 14964 20360 15028 20364
rect 14964 20304 15014 20360
rect 15014 20304 15028 20360
rect 14964 20300 15028 20304
rect 15516 20300 15580 20364
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 19748 19892 19812 19956
rect 22140 19892 22204 19956
rect 10548 19816 10612 19820
rect 10548 19760 10562 19816
rect 10562 19760 10612 19816
rect 10548 19756 10612 19760
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18828 19348 18892 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 18644 18864 18708 18868
rect 18644 18808 18694 18864
rect 18694 18808 18708 18864
rect 18644 18804 18708 18808
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 14780 18456 14844 18460
rect 14780 18400 14794 18456
rect 14794 18400 14844 18456
rect 14780 18396 14844 18400
rect 19932 17988 19996 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 13492 17580 13556 17644
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 16436 16824 16500 16828
rect 16436 16768 16450 16824
rect 16450 16768 16500 16824
rect 16436 16764 16500 16768
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 15700 15268 15764 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 17540 15192 17604 15196
rect 17540 15136 17554 15192
rect 17554 15136 17604 15192
rect 17540 15132 17604 15136
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 12572 13364 12636 13428
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 12020 12956 12084 13020
rect 22324 12820 22388 12884
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 22140 11928 22204 11932
rect 22140 11872 22154 11928
rect 22154 11872 22204 11928
rect 22140 11868 22204 11872
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 14964 10916 15028 10980
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 14044 7924 14108 7988
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18828 4040 18892 4044
rect 18828 3984 18842 4040
rect 18842 3984 18892 4040
rect 18828 3980 18892 3984
rect 22324 3980 22388 4044
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 10180 3572 10244 3636
rect 10548 3436 10612 3500
rect 23428 3436 23492 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 12204 3164 12268 3228
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 9076 2620 9140 2684
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 12944 53888 13264 54448
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17171 53956 17237 53957
rect 17171 53892 17172 53956
rect 17236 53892 17237 53956
rect 17171 53891 17237 53892
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 14043 52596 14109 52597
rect 14043 52532 14044 52596
rect 14108 52532 14109 52596
rect 14043 52531 14109 52532
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12203 45252 12269 45253
rect 12203 45188 12204 45252
rect 12268 45188 12269 45252
rect 12203 45187 12269 45188
rect 10547 44708 10613 44709
rect 10547 44644 10548 44708
rect 10612 44644 10613 44708
rect 10547 44643 10613 44644
rect 11099 44708 11165 44709
rect 11099 44644 11100 44708
rect 11164 44644 11165 44708
rect 11099 44643 11165 44644
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 9443 44300 9509 44301
rect 9443 44236 9444 44300
rect 9508 44236 9509 44300
rect 9443 44235 9509 44236
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 9446 36685 9506 44235
rect 10179 42260 10245 42261
rect 10179 42196 10180 42260
rect 10244 42196 10245 42260
rect 10179 42195 10245 42196
rect 9443 36684 9509 36685
rect 9443 36620 9444 36684
rect 9508 36620 9509 36684
rect 9443 36619 9509 36620
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 10182 34781 10242 42195
rect 10550 39133 10610 44643
rect 10547 39132 10613 39133
rect 10547 39068 10548 39132
rect 10612 39068 10613 39132
rect 10547 39067 10613 39068
rect 10179 34780 10245 34781
rect 10179 34716 10180 34780
rect 10244 34716 10245 34780
rect 10179 34715 10245 34716
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 10550 30429 10610 39067
rect 11102 34917 11162 44643
rect 11651 44300 11717 44301
rect 11651 44236 11652 44300
rect 11716 44236 11717 44300
rect 11651 44235 11717 44236
rect 11099 34916 11165 34917
rect 11099 34852 11100 34916
rect 11164 34852 11165 34916
rect 11099 34851 11165 34852
rect 11654 32333 11714 44235
rect 12206 38453 12266 45187
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 13675 38996 13741 38997
rect 13675 38932 13676 38996
rect 13740 38932 13741 38996
rect 13675 38931 13741 38932
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12203 38452 12269 38453
rect 12203 38388 12204 38452
rect 12268 38388 12269 38452
rect 12203 38387 12269 38388
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12571 33420 12637 33421
rect 12571 33356 12572 33420
rect 12636 33356 12637 33420
rect 12571 33355 12637 33356
rect 11651 32332 11717 32333
rect 11651 32268 11652 32332
rect 11716 32268 11717 32332
rect 11651 32267 11717 32268
rect 10547 30428 10613 30429
rect 10547 30364 10548 30428
rect 10612 30364 10613 30428
rect 10547 30363 10613 30364
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 12203 29340 12269 29341
rect 12203 29276 12204 29340
rect 12268 29276 12269 29340
rect 12203 29275 12269 29276
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 9075 26756 9141 26757
rect 9075 26692 9076 26756
rect 9140 26692 9141 26756
rect 9075 26691 9141 26692
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 9078 2685 9138 26691
rect 10547 25124 10613 25125
rect 10547 25060 10548 25124
rect 10612 25060 10613 25124
rect 10547 25059 10613 25060
rect 10179 21316 10245 21317
rect 10179 21252 10180 21316
rect 10244 21252 10245 21316
rect 10179 21251 10245 21252
rect 10182 3637 10242 21251
rect 10550 19821 10610 25059
rect 12019 22676 12085 22677
rect 12019 22612 12020 22676
rect 12084 22612 12085 22676
rect 12019 22611 12085 22612
rect 10547 19820 10613 19821
rect 10547 19756 10548 19820
rect 10612 19756 10613 19820
rect 10547 19755 10613 19756
rect 10179 3636 10245 3637
rect 10179 3572 10180 3636
rect 10244 3572 10245 3636
rect 10179 3571 10245 3572
rect 10550 3501 10610 19755
rect 12022 13021 12082 22611
rect 12019 13020 12085 13021
rect 12019 12956 12020 13020
rect 12084 12956 12085 13020
rect 12019 12955 12085 12956
rect 10547 3500 10613 3501
rect 10547 3436 10548 3500
rect 10612 3436 10613 3500
rect 10547 3435 10613 3436
rect 12206 3229 12266 29275
rect 12574 13429 12634 33355
rect 12944 33216 13264 34240
rect 13491 33284 13557 33285
rect 13491 33220 13492 33284
rect 13556 33220 13557 33284
rect 13491 33219 13557 33220
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 13494 17645 13554 33219
rect 13678 23221 13738 38931
rect 14046 34509 14106 52531
rect 15515 38860 15581 38861
rect 15515 38796 15516 38860
rect 15580 38796 15581 38860
rect 15515 38795 15581 38796
rect 14779 37364 14845 37365
rect 14779 37300 14780 37364
rect 14844 37300 14845 37364
rect 14779 37299 14845 37300
rect 14782 35733 14842 37299
rect 14779 35732 14845 35733
rect 14779 35668 14780 35732
rect 14844 35668 14845 35732
rect 14779 35667 14845 35668
rect 14043 34508 14109 34509
rect 14043 34444 14044 34508
rect 14108 34444 14109 34508
rect 14043 34443 14109 34444
rect 13675 23220 13741 23221
rect 13675 23156 13676 23220
rect 13740 23156 13741 23220
rect 13675 23155 13741 23156
rect 14043 21316 14109 21317
rect 14043 21252 14044 21316
rect 14108 21252 14109 21316
rect 14043 21251 14109 21252
rect 13491 17644 13557 17645
rect 13491 17580 13492 17644
rect 13556 17580 13557 17644
rect 13491 17579 13557 17580
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12571 13428 12637 13429
rect 12571 13364 12572 13428
rect 12636 13364 12637 13428
rect 12571 13363 12637 13364
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 14046 7989 14106 21251
rect 14782 18461 14842 35667
rect 14963 34644 15029 34645
rect 14963 34580 14964 34644
rect 15028 34580 15029 34644
rect 14963 34579 15029 34580
rect 14966 34101 15026 34579
rect 14963 34100 15029 34101
rect 14963 34036 14964 34100
rect 15028 34036 15029 34100
rect 14963 34035 15029 34036
rect 14966 20365 15026 34035
rect 15518 20365 15578 38795
rect 16803 29068 16869 29069
rect 16803 29004 16804 29068
rect 16868 29004 16869 29068
rect 16803 29003 16869 29004
rect 16435 28116 16501 28117
rect 16435 28052 16436 28116
rect 16500 28052 16501 28116
rect 16435 28051 16501 28052
rect 15699 26212 15765 26213
rect 15699 26148 15700 26212
rect 15764 26148 15765 26212
rect 15699 26147 15765 26148
rect 14963 20364 15029 20365
rect 14963 20300 14964 20364
rect 15028 20300 15029 20364
rect 14963 20299 15029 20300
rect 15515 20364 15581 20365
rect 15515 20300 15516 20364
rect 15580 20300 15581 20364
rect 15515 20299 15581 20300
rect 14779 18460 14845 18461
rect 14779 18396 14780 18460
rect 14844 18396 14845 18460
rect 14779 18395 14845 18396
rect 14966 10981 15026 20299
rect 15702 15333 15762 26147
rect 16438 16829 16498 28051
rect 16806 22133 16866 29003
rect 17174 27709 17234 53891
rect 17944 53344 18264 54368
rect 21955 53956 22021 53957
rect 21955 53892 21956 53956
rect 22020 53892 22021 53956
rect 21955 53891 22021 53892
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 18827 47156 18893 47157
rect 18827 47092 18828 47156
rect 18892 47092 18893 47156
rect 18827 47091 18893 47092
rect 19195 47156 19261 47157
rect 19195 47092 19196 47156
rect 19260 47092 19261 47156
rect 19195 47091 19261 47092
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17723 40764 17789 40765
rect 17723 40700 17724 40764
rect 17788 40700 17789 40764
rect 17723 40699 17789 40700
rect 17539 31380 17605 31381
rect 17539 31316 17540 31380
rect 17604 31316 17605 31380
rect 17539 31315 17605 31316
rect 17542 27845 17602 31315
rect 17726 28117 17786 40699
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 18830 39813 18890 47091
rect 18827 39812 18893 39813
rect 18827 39748 18828 39812
rect 18892 39748 18893 39812
rect 18827 39747 18893 39748
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 18643 30156 18709 30157
rect 18643 30092 18644 30156
rect 18708 30092 18709 30156
rect 18643 30091 18709 30092
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17723 28116 17789 28117
rect 17723 28052 17724 28116
rect 17788 28052 17789 28116
rect 17723 28051 17789 28052
rect 17539 27844 17605 27845
rect 17539 27780 17540 27844
rect 17604 27780 17605 27844
rect 17539 27779 17605 27780
rect 17171 27708 17237 27709
rect 17171 27644 17172 27708
rect 17236 27644 17237 27708
rect 17171 27643 17237 27644
rect 16803 22132 16869 22133
rect 16803 22068 16804 22132
rect 16868 22068 16869 22132
rect 16803 22067 16869 22068
rect 16435 16828 16501 16829
rect 16435 16764 16436 16828
rect 16500 16764 16501 16828
rect 16435 16763 16501 16764
rect 15699 15332 15765 15333
rect 15699 15268 15700 15332
rect 15764 15268 15765 15332
rect 15699 15267 15765 15268
rect 17542 15197 17602 27779
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 18646 18869 18706 30091
rect 18830 21181 18890 39747
rect 19198 33285 19258 47091
rect 19931 47020 19997 47021
rect 19931 46956 19932 47020
rect 19996 46956 19997 47020
rect 19931 46955 19997 46956
rect 19195 33284 19261 33285
rect 19195 33220 19196 33284
rect 19260 33220 19261 33284
rect 19195 33219 19261 33220
rect 19934 30701 19994 46955
rect 21771 44708 21837 44709
rect 21771 44644 21772 44708
rect 21836 44644 21837 44708
rect 21771 44643 21837 44644
rect 20299 43076 20365 43077
rect 20299 43012 20300 43076
rect 20364 43012 20365 43076
rect 20299 43011 20365 43012
rect 19931 30700 19997 30701
rect 19931 30636 19932 30700
rect 19996 30636 19997 30700
rect 19931 30635 19997 30636
rect 19747 27300 19813 27301
rect 19747 27236 19748 27300
rect 19812 27236 19813 27300
rect 19747 27235 19813 27236
rect 18827 21180 18893 21181
rect 18827 21116 18828 21180
rect 18892 21116 18893 21180
rect 18827 21115 18893 21116
rect 19750 19957 19810 27235
rect 19747 19956 19813 19957
rect 19747 19892 19748 19956
rect 19812 19892 19813 19956
rect 19747 19891 19813 19892
rect 18827 19412 18893 19413
rect 18827 19348 18828 19412
rect 18892 19348 18893 19412
rect 18827 19347 18893 19348
rect 18643 18868 18709 18869
rect 18643 18804 18644 18868
rect 18708 18804 18709 18868
rect 18643 18803 18709 18804
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17539 15196 17605 15197
rect 17539 15132 17540 15196
rect 17604 15132 17605 15196
rect 17539 15131 17605 15132
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 14963 10980 15029 10981
rect 14963 10916 14964 10980
rect 15028 10916 15029 10980
rect 14963 10915 15029 10916
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 14043 7988 14109 7989
rect 14043 7924 14044 7988
rect 14108 7924 14109 7988
rect 14043 7923 14109 7924
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12203 3228 12269 3229
rect 12203 3164 12204 3228
rect 12268 3164 12269 3228
rect 12203 3163 12269 3164
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 9075 2684 9141 2685
rect 9075 2620 9076 2684
rect 9140 2620 9141 2684
rect 9075 2619 9141 2620
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 2128 13264 2688
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 18830 4045 18890 19347
rect 19934 18053 19994 30635
rect 20302 30429 20362 43011
rect 20667 40084 20733 40085
rect 20667 40020 20668 40084
rect 20732 40020 20733 40084
rect 20667 40019 20733 40020
rect 20670 34645 20730 40019
rect 21587 39540 21653 39541
rect 21587 39476 21588 39540
rect 21652 39476 21653 39540
rect 21587 39475 21653 39476
rect 21590 38453 21650 39475
rect 21587 38452 21653 38453
rect 21587 38388 21588 38452
rect 21652 38388 21653 38452
rect 21587 38387 21653 38388
rect 20667 34644 20733 34645
rect 20667 34580 20668 34644
rect 20732 34580 20733 34644
rect 20667 34579 20733 34580
rect 21590 31517 21650 38387
rect 21587 31516 21653 31517
rect 21587 31452 21588 31516
rect 21652 31452 21653 31516
rect 21587 31451 21653 31452
rect 20299 30428 20365 30429
rect 20299 30364 20300 30428
rect 20364 30364 20365 30428
rect 20299 30363 20365 30364
rect 21774 28253 21834 44643
rect 21958 32061 22018 53891
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 23979 52596 24045 52597
rect 23979 52532 23980 52596
rect 24044 52532 24045 52596
rect 23979 52531 24045 52532
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22691 47020 22757 47021
rect 22691 46956 22692 47020
rect 22756 46956 22757 47020
rect 22691 46955 22757 46956
rect 22694 41173 22754 46955
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 23611 44436 23677 44437
rect 23611 44372 23612 44436
rect 23676 44372 23677 44436
rect 23611 44371 23677 44372
rect 23427 44300 23493 44301
rect 23427 44236 23428 44300
rect 23492 44236 23493 44300
rect 23427 44235 23493 44236
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22691 41172 22757 41173
rect 22691 41108 22692 41172
rect 22756 41108 22757 41172
rect 22691 41107 22757 41108
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22323 40084 22389 40085
rect 22323 40020 22324 40084
rect 22388 40020 22389 40084
rect 22323 40019 22389 40020
rect 22326 36957 22386 40019
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 23430 39541 23490 44235
rect 23427 39540 23493 39541
rect 23427 39476 23428 39540
rect 23492 39476 23493 39540
rect 23427 39475 23493 39476
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 23614 38453 23674 44371
rect 23611 38452 23677 38453
rect 23611 38388 23612 38452
rect 23676 38388 23677 38452
rect 23611 38387 23677 38388
rect 23982 38045 24042 52531
rect 23979 38044 24045 38045
rect 23979 37980 23980 38044
rect 24044 37980 24045 38044
rect 23979 37979 24045 37980
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22323 36956 22389 36957
rect 22323 36892 22324 36956
rect 22388 36892 22389 36956
rect 22323 36891 22389 36892
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 21955 32060 22021 32061
rect 21955 31996 21956 32060
rect 22020 31996 22021 32060
rect 21955 31995 22021 31996
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 21771 28252 21837 28253
rect 21771 28188 21772 28252
rect 21836 28188 21837 28252
rect 21771 28187 21837 28188
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 23427 22132 23493 22133
rect 23427 22068 23428 22132
rect 23492 22068 23493 22132
rect 23427 22067 23493 22068
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22139 19956 22205 19957
rect 22139 19892 22140 19956
rect 22204 19892 22205 19956
rect 22139 19891 22205 19892
rect 19931 18052 19997 18053
rect 19931 17988 19932 18052
rect 19996 17988 19997 18052
rect 19931 17987 19997 17988
rect 22142 11933 22202 19891
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22323 12884 22389 12885
rect 22323 12820 22324 12884
rect 22388 12820 22389 12884
rect 22323 12819 22389 12820
rect 22139 11932 22205 11933
rect 22139 11868 22140 11932
rect 22204 11868 22205 11932
rect 22139 11867 22205 11868
rect 22326 4045 22386 12819
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 18827 4044 18893 4045
rect 18827 3980 18828 4044
rect 18892 3980 18893 4044
rect 18827 3979 18893 3980
rect 22323 4044 22389 4045
rect 22323 3980 22324 4044
rect 22388 3980 22389 4044
rect 22323 3979 22389 3980
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 23430 3501 23490 22067
rect 23427 3500 23493 3501
rect 23427 3436 23428 3500
rect 23492 3436 23493 3500
rect 23427 3435 23493 3436
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 24932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _110_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23184 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform -1 0 24932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1679235063
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1679235063
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1679235063
transform -1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 16008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1679235063
transform -1 0 23552 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1679235063
transform -1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1679235063
transform -1 0 22264 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 23276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 22632 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 23184 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1679235063
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 23552 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1679235063
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 23736 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1679235063
transform -1 0 24104 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform -1 0 22632 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1679235063
transform -1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 24564 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1679235063
transform 1 0 24656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform -1 0 24932 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform -1 0 24932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _137_
timestamp 1679235063
transform -1 0 21528 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform -1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform -1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 13248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 11868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform -1 0 14628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform -1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 15640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform -1 0 21068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1679235063
transform 1 0 21988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1679235063
transform 1 0 18308 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 20424 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1679235063
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1679235063
transform -1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1679235063
transform -1 0 3772 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1679235063
transform -1 0 4508 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1679235063
transform -1 0 4876 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1679235063
transform -1 0 7912 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1679235063
transform -1 0 5060 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1679235063
transform -1 0 5244 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1679235063
transform -1 0 6072 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1679235063
transform -1 0 9476 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1679235063
transform -1 0 6900 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1679235063
transform -1 0 6900 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1679235063
transform -1 0 7636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_
timestamp 1679235063
transform -1 0 7544 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1679235063
transform -1 0 8096 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1679235063
transform -1 0 8372 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1679235063
transform -1 0 9476 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp 1679235063
transform -1 0 7176 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1679235063
transform -1 0 9476 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1679235063
transform -1 0 9384 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1679235063
transform -1 0 10672 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1679235063
transform 1 0 9200 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1679235063
transform -1 0 11224 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1679235063
transform -1 0 11408 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1679235063
transform -1 0 12052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1679235063
transform 1 0 9200 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1679235063
transform 1 0 9292 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1679235063
transform -1 0 12328 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1679235063
transform 1 0 10212 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1679235063
transform -1 0 11960 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1679235063
transform 1 0 12604 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1679235063
transform -1 0 12604 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1679235063
transform -1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _199_
timestamp 1679235063
transform -1 0 2392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1679235063
transform 1 0 1748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 14168 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1679235063
transform -1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform -1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform -1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform -1 0 16468 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform -1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform -1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform -1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 18860 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 18216 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1679235063
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1679235063
transform -1 0 23368 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1679235063
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1679235063
transform 1 0 3036 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1679235063
transform 1 0 3956 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1679235063
transform -1 0 5244 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1679235063
transform -1 0 5428 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1679235063
transform 1 0 5428 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1679235063
transform -1 0 6440 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1679235063
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1679235063
transform -1 0 6532 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1679235063
transform 1 0 7084 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1679235063
transform -1 0 8464 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1679235063
transform 1 0 7636 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1679235063
transform -1 0 9844 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1679235063
transform -1 0 9844 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1679235063
transform 1 0 8648 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1679235063
transform -1 0 10120 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1679235063
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1679235063
transform -1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1679235063
transform 1 0 12236 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1679235063
transform -1 0 11776 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8464 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform -1 0 11408 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8740 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11500 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14628 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 14444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 13708 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12328 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1679235063
transform -1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 10396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14352 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 14996 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform -1 0 9384 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 12512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform -1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13248 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 15180 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform -1 0 13524 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 13064 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 10764 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 2484 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5796 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 4324 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1679235063
transform 1 0 7176 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform -1 0 6256 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 12052 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 9660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 11776 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform -1 0 21896 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 20332 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 19320 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 10488 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 13248 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 20976 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 21252 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform -1 0 21068 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout203_A
timestamp 1679235063
transform 1 0 22264 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout204_A
timestamp 1679235063
transform 1 0 16284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout205_A
timestamp 1679235063
transform 1 0 13524 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout206_A
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout207_A
timestamp 1679235063
transform -1 0 25484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout208_A
timestamp 1679235063
transform -1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout209_A
timestamp 1679235063
transform 1 0 15272 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout210_A
timestamp 1679235063
transform 1 0 11040 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout211_A
timestamp 1679235063
transform -1 0 25576 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout212_A
timestamp 1679235063
transform 1 0 16192 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout213_A
timestamp 1679235063
transform 1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout214_A
timestamp 1679235063
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout215_A
timestamp 1679235063
transform -1 0 24748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold126_A
timestamp 1679235063
transform -1 0 7636 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold129_A
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform -1 0 21988 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform -1 0 24288 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform -1 0 20976 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 21436 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform -1 0 24288 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform -1 0 21712 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform -1 0 20884 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform -1 0 23184 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 23368 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform -1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform -1 0 25208 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform -1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform -1 0 23184 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform -1 0 24288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform -1 0 25576 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform -1 0 24564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 25208 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform -1 0 25576 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform -1 0 24932 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform -1 0 24932 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform -1 0 24748 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform -1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 24196 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform -1 0 23644 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform -1 0 22816 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform -1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform -1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform -1 0 24564 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform -1 0 25576 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform -1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform -1 0 6256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform -1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform -1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform -1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform -1 0 8832 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform -1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform -1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform -1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform -1 0 9844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform -1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform -1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform -1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform -1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform -1 0 11408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform -1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform -1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform -1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform -1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform -1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform -1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform -1 0 4232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform -1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform -1 0 5980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform -1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform -1 0 14260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform -1 0 16468 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform -1 0 19044 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform -1 0 17388 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform -1 0 19044 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform -1 0 18860 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform -1 0 19872 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform -1 0 19504 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform -1 0 19688 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform -1 0 21620 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform -1 0 20884 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform -1 0 13340 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform -1 0 20976 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform -1 0 21344 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1679235063
transform -1 0 21160 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1679235063
transform -1 0 23460 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform -1 0 21988 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform -1 0 22448 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1679235063
transform -1 0 22724 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1679235063
transform -1 0 24564 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1679235063
transform -1 0 23092 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1679235063
transform -1 0 24564 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1679235063
transform -1 0 14260 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1679235063
transform -1 0 14996 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1679235063
transform -1 0 15088 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1679235063
transform -1 0 14628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1679235063
transform -1 0 16284 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1679235063
transform -1 0 16284 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1679235063
transform -1 0 16560 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1679235063
transform -1 0 16560 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1679235063
transform -1 0 2208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1679235063
transform -1 0 2208 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1679235063
transform -1 0 2208 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1679235063
transform -1 0 2208 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1679235063
transform -1 0 2300 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1679235063
transform -1 0 25300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1679235063
transform -1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1679235063
transform -1 0 25576 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1679235063
transform -1 0 24840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1679235063
transform -1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1679235063
transform -1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1679235063
transform -1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1679235063
transform -1 0 24748 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1679235063
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output107_A
timestamp 1679235063
transform -1 0 21712 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output108_A
timestamp 1679235063
transform -1 0 3404 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output141_A
timestamp 1679235063
transform -1 0 18676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output147_A
timestamp 1679235063
transform -1 0 21712 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21160 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19504 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 22080 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform -1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14628 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform -1 0 16468 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16928 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform -1 0 21620 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform -1 0 16008 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10488 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24656 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15088 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14444 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12604 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11776 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11132 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15272 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform -1 0 16284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform -1 0 24288 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8648 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11868 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16284 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform -1 0 14352 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform -1 0 16192 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11408 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11776 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 9476 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 6992 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7820 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10120 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11868 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 7452 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9016 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8280 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10120 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17112 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18492 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1679235063
transform -1 0 19964 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 19780 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 16008 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 20608 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21160 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 21712 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 17848 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19044 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 23184 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 20424 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 18768 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 20700 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 19504 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11776 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17020 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 17848 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19320 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 21344 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 23368 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17756 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 21436 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20608 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 20976 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11592 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20240 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21896 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21896 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 23000 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23460 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 20884 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21988 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 21160 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 20424 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21436 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21804 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24012 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 19504 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21344 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 23184 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 20884 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20884 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 22448 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18676 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 21436 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 21988 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20608 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 20240 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1
timestamp 1679235063
transform -1 0 18584 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 18216 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16192 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18216 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 18400 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 14168 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17664 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 18584 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1
timestamp 1679235063
transform -1 0 14260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16192 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 15640 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11960 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13800 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 13800 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11684 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15272 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10948 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16192 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8924 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13248 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 7636 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14260 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10120 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 17848 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12144 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15456 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15640 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 15364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 20240 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8004 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9568 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 10212 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18308 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 16744 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14536 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 14628 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 9200 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 9384 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18124 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 18492 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 12052 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 12236 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17848 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 18308 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 10856 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8832 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8648 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18400 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 17020 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 13616 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__S
timestamp 1679235063
transform -1 0 13984 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 7636 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 9016 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 10304 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 10856 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__S
timestamp 1679235063
transform -1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16928 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 15916 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 12236 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__S
timestamp 1679235063
transform -1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 6900 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13616 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 12052 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 8004 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 8004 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15732 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14352 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 8648 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 8832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13708 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12328 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 14076 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 4876 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12696 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform -1 0 13432 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 8004 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10396 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3956 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 10948 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 8372 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 5336 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7544 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 13524 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 8648 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6716 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7912 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 11224 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 8004 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 5060 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9384 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 8464 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform -1 0 7176 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12880 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10212 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10304 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10028 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__262 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9568 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7452 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 6532 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14720 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14720 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 13984 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12604 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9568 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__263
timestamp 1679235063
transform 1 0 12880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10304 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7912 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7360 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4324 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13984 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10028 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__264
timestamp 1679235063
transform -1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9108 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 8832 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7268 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 5980 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3680 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13616 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13432 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13524 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12052 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 8832 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__265
timestamp 1679235063
transform -1 0 10028 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 8648 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 5428 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 4140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3772 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 4600 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform -1 0 3496 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 6256 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 4048 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform -1 0 3496 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform -1 0 3772 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 5612 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 4232 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform -1 0 5152 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform -1 0 3496 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 4324 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 3956 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 4048 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform -1 0 7176 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform -1 0 4324 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9844 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 16560 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 10120 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform -1 0 11868 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform -1 0 9476 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 10764 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform -1 0 18952 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 20424 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform -1 0 20884 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 19872 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform -1 0 10120 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform -1 0 11224 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 9660 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 12052 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform -1 0 20424 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 21436 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform -1 0 20424 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 21436 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout202
timestamp 1679235063
transform -1 0 15364 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout203
timestamp 1679235063
transform 1 0 21068 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout204
timestamp 1679235063
transform 1 0 14812 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout205 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 13340 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout206
timestamp 1679235063
transform 1 0 24196 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout207
timestamp 1679235063
transform -1 0 25116 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout208
timestamp 1679235063
transform -1 0 21528 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout209 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14260 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout210 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 10672 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout211
timestamp 1679235063
transform -1 0 25392 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout212
timestamp 1679235063
transform 1 0 14444 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout213
timestamp 1679235063
transform -1 0 25392 0 -1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout214
timestamp 1679235063
transform -1 0 23920 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout215
timestamp 1679235063
transform 1 0 24564 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1679235063
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1679235063
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61
timestamp 1679235063
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1679235063
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1679235063
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90
timestamp 1679235063
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1679235063
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1679235063
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1679235063
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1679235063
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1679235063
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1679235063
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1679235063
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1679235063
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1679235063
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1679235063
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1679235063
transform 1 0 24932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263
timestamp 1679235063
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1679235063
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35
timestamp 1679235063
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1679235063
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1679235063
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_59
timestamp 1679235063
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1679235063
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1679235063
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1679235063
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1679235063
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1679235063
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1679235063
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1679235063
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1679235063
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_219
timestamp 1679235063
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1679235063
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_263
timestamp 1679235063
transform 1 0 25300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_5
timestamp 1679235063
transform 1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_20
timestamp 1679235063
transform 1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1679235063
transform 1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1679235063
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_51
timestamp 1679235063
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1679235063
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_63
timestamp 1679235063
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_68
timestamp 1679235063
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_73
timestamp 1679235063
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_79
timestamp 1679235063
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 1679235063
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1679235063
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1679235063
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1679235063
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1679235063
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1679235063
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1679235063
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_235
timestamp 1679235063
transform 1 0 22724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1679235063
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1679235063
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_265
timestamp 1679235063
transform 1 0 25484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1679235063
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_17
timestamp 1679235063
transform 1 0 2668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_28
timestamp 1679235063
transform 1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_34
timestamp 1679235063
transform 1 0 4232 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_37
timestamp 1679235063
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59
timestamp 1679235063
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_71
timestamp 1679235063
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_83
timestamp 1679235063
transform 1 0 8740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_95
timestamp 1679235063
transform 1 0 9844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_98
timestamp 1679235063
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1679235063
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1679235063
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_151
timestamp 1679235063
transform 1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_159
timestamp 1679235063
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1679235063
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1679235063
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1679235063
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1679235063
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1679235063
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1679235063
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 1679235063
transform 1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_14
timestamp 1679235063
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1679235063
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1679235063
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_34
timestamp 1679235063
transform 1 0 4232 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_46
timestamp 1679235063
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 1679235063
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1679235063
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1679235063
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1679235063
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_239
timestamp 1679235063
transform 1 0 23092 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1679235063
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_5
timestamp 1679235063
transform 1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_10
timestamp 1679235063
transform 1 0 2024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_14
timestamp 1679235063
transform 1 0 2392 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1679235063
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1679235063
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1679235063
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_199
timestamp 1679235063
transform 1 0 19412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1679235063
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1679235063
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1679235063
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1679235063
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1679235063
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1679235063
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1679235063
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_205
timestamp 1679235063
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1679235063
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_243
timestamp 1679235063
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1679235063
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1679235063
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_29
timestamp 1679235063
transform 1 0 3772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_41
timestamp 1679235063
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1679235063
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1679235063
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_197
timestamp 1679235063
transform 1 0 19228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1679235063
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1679235063
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1679235063
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_204
timestamp 1679235063
transform 1 0 19872 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1679235063
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1679235063
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_258
timestamp 1679235063
transform 1 0 24840 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1679235063
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_181
timestamp 1679235063
transform 1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_191
timestamp 1679235063
transform 1 0 18676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_203
timestamp 1679235063
transform 1 0 19780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_209
timestamp 1679235063
transform 1 0 20332 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_213
timestamp 1679235063
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1679235063
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_54
timestamp 1679235063
transform 1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1679235063
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_70
timestamp 1679235063
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1679235063
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1679235063
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1679235063
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1679235063
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1679235063
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_203
timestamp 1679235063
transform 1 0 19780 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_215
timestamp 1679235063
transform 1 0 20884 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1679235063
transform 1 0 21436 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_225
timestamp 1679235063
transform 1 0 21804 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_233
timestamp 1679235063
transform 1 0 22540 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1679235063
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1679235063
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_65
timestamp 1679235063
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_77
timestamp 1679235063
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_89
timestamp 1679235063
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_101
timestamp 1679235063
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1679235063
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1679235063
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1679235063
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1679235063
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1679235063
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1679235063
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1679235063
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_217
timestamp 1679235063
transform 1 0 21068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_221
timestamp 1679235063
transform 1 0 21436 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_65
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1679235063
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1679235063
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1679235063
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1679235063
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1679235063
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1679235063
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1679235063
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_171
timestamp 1679235063
transform 1 0 16836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_183
timestamp 1679235063
transform 1 0 17940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1679235063
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_203
timestamp 1679235063
transform 1 0 19780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_215
timestamp 1679235063
transform 1 0 20884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_227
timestamp 1679235063
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_239
timestamp 1679235063
transform 1 0 23092 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_245
timestamp 1679235063
transform 1 0 23644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1679235063
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_259
timestamp 1679235063
transform 1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1679235063
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1679235063
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1679235063
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1679235063
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1679235063
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_137
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1679235063
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1679235063
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1679235063
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1679235063
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1679235063
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1679235063
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1679235063
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1679235063
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_233
timestamp 1679235063
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1679235063
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1679235063
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1679235063
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1679235063
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1679235063
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1679235063
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1679235063
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1679235063
transform 1 0 16652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_174
timestamp 1679235063
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp 1679235063
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1679235063
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_221
timestamp 1679235063
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1679235063
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_259
timestamp 1679235063
transform 1 0 24932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_265
timestamp 1679235063
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1679235063
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1679235063
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_115
timestamp 1679235063
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_121
timestamp 1679235063
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_126
timestamp 1679235063
transform 1 0 12696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_138
timestamp 1679235063
transform 1 0 13800 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1679235063
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1679235063
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1679235063
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1679235063
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1679235063
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_206
timestamp 1679235063
transform 1 0 20056 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_213
timestamp 1679235063
transform 1 0 20700 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1679235063
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_230
timestamp 1679235063
transform 1 0 22264 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_238
timestamp 1679235063
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1679235063
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1679235063
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_103
timestamp 1679235063
transform 1 0 10580 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_124
timestamp 1679235063
transform 1 0 12512 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_136
timestamp 1679235063
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1679235063
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1679235063
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1679235063
transform 1 0 16008 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_169
timestamp 1679235063
transform 1 0 16652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_181
timestamp 1679235063
transform 1 0 17756 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1679235063
transform 1 0 18676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1679235063
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1679235063
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1679235063
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_223
timestamp 1679235063
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_227
timestamp 1679235063
transform 1 0 21988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_239
timestamp 1679235063
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1679235063
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1679235063
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1679235063
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1679235063
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1679235063
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1679235063
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1679235063
transform 1 0 15364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1679235063
transform 1 0 16100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1679235063
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1679235063
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1679235063
transform 1 0 18032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1679235063
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1679235063
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1679235063
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_231
timestamp 1679235063
transform 1 0 22356 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_238
timestamp 1679235063
transform 1 0 23000 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_242
timestamp 1679235063
transform 1 0 23368 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1679235063
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_110
timestamp 1679235063
transform 1 0 11224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_122
timestamp 1679235063
transform 1 0 12328 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_163
timestamp 1679235063
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_175
timestamp 1679235063
transform 1 0 17204 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1679235063
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1679235063
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1679235063
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_231
timestamp 1679235063
transform 1 0 22356 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_239
timestamp 1679235063
transform 1 0 23092 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_243
timestamp 1679235063
transform 1 0 23460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1679235063
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1679235063
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1679235063
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1679235063
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1679235063
transform 1 0 10764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1679235063
transform 1 0 11132 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1679235063
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_122
timestamp 1679235063
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_128
timestamp 1679235063
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_136
timestamp 1679235063
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_149
timestamp 1679235063
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1679235063
transform 1 0 15364 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1679235063
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1679235063
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1679235063
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1679235063
transform 1 0 18032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_205
timestamp 1679235063
transform 1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_209
timestamp 1679235063
transform 1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_214
timestamp 1679235063
transform 1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1679235063
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1679235063
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_247
timestamp 1679235063
transform 1 0 23828 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1679235063
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1679235063
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1679235063
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1679235063
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1679235063
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_95
timestamp 1679235063
transform 1 0 9844 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_107
timestamp 1679235063
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 1679235063
transform 1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1679235063
transform 1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1679235063
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1679235063
transform 1 0 14444 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1679235063
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1679235063
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1679235063
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_199
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_205
timestamp 1679235063
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1679235063
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_214
timestamp 1679235063
transform 1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_228
timestamp 1679235063
transform 1 0 22080 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1679235063
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1679235063
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1679235063
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1679235063
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1679235063
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1679235063
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_73
timestamp 1679235063
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1679235063
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_101
timestamp 1679235063
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1679235063
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1679235063
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1679235063
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1679235063
transform 1 0 14536 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_150
timestamp 1679235063
transform 1 0 14904 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_155
timestamp 1679235063
transform 1 0 15364 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1679235063
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1679235063
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1679235063
transform 1 0 17388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_185
timestamp 1679235063
transform 1 0 18124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_189
timestamp 1679235063
transform 1 0 18492 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_200
timestamp 1679235063
transform 1 0 19504 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1679235063
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1679235063
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1679235063
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_244
timestamp 1679235063
transform 1 0 23552 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1679235063
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_87
timestamp 1679235063
transform 1 0 9108 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1679235063
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_120
timestamp 1679235063
transform 1 0 12144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1679235063
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1679235063
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1679235063
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_189
timestamp 1679235063
transform 1 0 18492 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_193
timestamp 1679235063
transform 1 0 18860 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1679235063
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_216
timestamp 1679235063
transform 1 0 20976 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_237
timestamp 1679235063
transform 1 0 22908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1679235063
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1679235063
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1679235063
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1679235063
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1679235063
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1679235063
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1679235063
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1679235063
transform 1 0 8556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_85
timestamp 1679235063
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1679235063
transform 1 0 12420 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_131
timestamp 1679235063
transform 1 0 13156 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_134
timestamp 1679235063
transform 1 0 13432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1679235063
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1679235063
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_157
timestamp 1679235063
transform 1 0 15548 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1679235063
transform 1 0 17204 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1679235063
transform 1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1679235063
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_194
timestamp 1679235063
transform 1 0 18952 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1679235063
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_227
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_233
timestamp 1679235063
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_238
timestamp 1679235063
transform 1 0 23000 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_246
timestamp 1679235063
transform 1 0 23736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1679235063
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1679235063
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1679235063
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_61
timestamp 1679235063
transform 1 0 6716 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1679235063
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1679235063
transform 1 0 9384 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_101
timestamp 1679235063
transform 1 0 10396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_109
timestamp 1679235063
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1679235063
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_135
timestamp 1679235063
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1679235063
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1679235063
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1679235063
transform 1 0 15548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1679235063
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1679235063
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1679235063
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1679235063
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_232
timestamp 1679235063
transform 1 0 22448 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1679235063
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1679235063
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1679235063
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1679235063
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1679235063
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1679235063
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_65
timestamp 1679235063
transform 1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_77
timestamp 1679235063
transform 1 0 8188 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_83
timestamp 1679235063
transform 1 0 8740 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_93
timestamp 1679235063
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_98
timestamp 1679235063
transform 1 0 10120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1679235063
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_123
timestamp 1679235063
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_135
timestamp 1679235063
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_147
timestamp 1679235063
transform 1 0 14628 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1679235063
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1679235063
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1679235063
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_181
timestamp 1679235063
transform 1 0 17756 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1679235063
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1679235063
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_197
timestamp 1679235063
transform 1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_210
timestamp 1679235063
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1679235063
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_247
timestamp 1679235063
transform 1 0 23828 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1679235063
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_53
timestamp 1679235063
transform 1 0 5980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_75
timestamp 1679235063
transform 1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_79
timestamp 1679235063
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_96
timestamp 1679235063
transform 1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_109
timestamp 1679235063
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_133
timestamp 1679235063
transform 1 0 13340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_137
timestamp 1679235063
transform 1 0 13708 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1679235063
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_165
timestamp 1679235063
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_168
timestamp 1679235063
transform 1 0 16560 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1679235063
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1679235063
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_199
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1679235063
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_209
timestamp 1679235063
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_215
timestamp 1679235063
transform 1 0 20884 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1679235063
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1679235063
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp 1679235063
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_11
timestamp 1679235063
transform 1 0 2116 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_16
timestamp 1679235063
transform 1 0 2576 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_28
timestamp 1679235063
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_40
timestamp 1679235063
transform 1 0 4784 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1679235063
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1679235063
transform 1 0 7544 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_83
timestamp 1679235063
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1679235063
transform 1 0 9936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_100
timestamp 1679235063
transform 1 0 10304 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_117
timestamp 1679235063
transform 1 0 11868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1679235063
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_136
timestamp 1679235063
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 1679235063
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_155
timestamp 1679235063
transform 1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_191
timestamp 1679235063
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_203
timestamp 1679235063
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1679235063
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1679235063
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1679235063
transform 1 0 23460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1679235063
transform 1 0 23828 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1679235063
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1679235063
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1679235063
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_63
timestamp 1679235063
transform 1 0 6900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1679235063
transform 1 0 8096 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1679235063
transform 1 0 10120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_104
timestamp 1679235063
transform 1 0 10672 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_117
timestamp 1679235063
transform 1 0 11868 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_121
timestamp 1679235063
transform 1 0 12236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1679235063
transform 1 0 12788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1679235063
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1679235063
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1679235063
transform 1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1679235063
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_199
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1679235063
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_245
timestamp 1679235063
transform 1 0 23644 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_249
timestamp 1679235063
transform 1 0 24012 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_263
timestamp 1679235063
transform 1 0 25300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1679235063
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1679235063
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1679235063
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1679235063
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1679235063
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1679235063
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_107
timestamp 1679235063
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1679235063
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_124
timestamp 1679235063
transform 1 0 12512 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1679235063
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1679235063
transform 1 0 14260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1679235063
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1679235063
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1679235063
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_204
timestamp 1679235063
transform 1 0 19872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_208
timestamp 1679235063
transform 1 0 20240 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1679235063
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1679235063
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1679235063
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1679235063
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1679235063
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1679235063
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1679235063
transform 1 0 6808 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_68
timestamp 1679235063
transform 1 0 7360 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_95
timestamp 1679235063
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_108
timestamp 1679235063
transform 1 0 11040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1679235063
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1679235063
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1679235063
transform 1 0 14996 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_155
timestamp 1679235063
transform 1 0 15364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_159
timestamp 1679235063
transform 1 0 15732 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_164
timestamp 1679235063
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_168
timestamp 1679235063
transform 1 0 16560 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_171
timestamp 1679235063
transform 1 0 16836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1679235063
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1679235063
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1679235063
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_220
timestamp 1679235063
transform 1 0 21344 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1679235063
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1679235063
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1679235063
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_14
timestamp 1679235063
transform 1 0 2392 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_26
timestamp 1679235063
transform 1 0 3496 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_38
timestamp 1679235063
transform 1 0 4600 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_50
timestamp 1679235063
transform 1 0 5704 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_66
timestamp 1679235063
transform 1 0 7176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1679235063
transform 1 0 9660 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1679235063
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_124
timestamp 1679235063
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_131
timestamp 1679235063
transform 1 0 13156 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1679235063
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_148
timestamp 1679235063
transform 1 0 14720 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_160
timestamp 1679235063
transform 1 0 15824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1679235063
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1679235063
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_185
timestamp 1679235063
transform 1 0 18124 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_189
timestamp 1679235063
transform 1 0 18492 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1679235063
transform 1 0 20976 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1679235063
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1679235063
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1679235063
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1679235063
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_53
timestamp 1679235063
transform 1 0 5980 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_62
timestamp 1679235063
transform 1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_70
timestamp 1679235063
transform 1 0 7544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1679235063
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1679235063
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1679235063
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_110
timestamp 1679235063
transform 1 0 11224 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_120
timestamp 1679235063
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_126
timestamp 1679235063
transform 1 0 12696 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_132
timestamp 1679235063
transform 1 0 13248 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1679235063
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1679235063
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1679235063
transform 1 0 16100 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_167
timestamp 1679235063
transform 1 0 16468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_173
timestamp 1679235063
transform 1 0 17020 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_181
timestamp 1679235063
transform 1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1679235063
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1679235063
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1679235063
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_218
timestamp 1679235063
transform 1 0 21160 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1679235063
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_257
timestamp 1679235063
transform 1 0 24748 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1679235063
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_31
timestamp 1679235063
transform 1 0 3956 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_38
timestamp 1679235063
transform 1 0 4600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_50
timestamp 1679235063
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1679235063
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_83
timestamp 1679235063
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1679235063
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_97
timestamp 1679235063
transform 1 0 10028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_124
timestamp 1679235063
transform 1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_128
timestamp 1679235063
transform 1 0 12880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_140
timestamp 1679235063
transform 1 0 13984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_146
timestamp 1679235063
transform 1 0 14536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_161
timestamp 1679235063
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1679235063
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1679235063
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_178
timestamp 1679235063
transform 1 0 17480 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1679235063
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1679235063
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1679235063
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_205
timestamp 1679235063
transform 1 0 19964 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_213
timestamp 1679235063
transform 1 0 20700 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_244
timestamp 1679235063
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1679235063
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1679235063
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1679235063
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_45
timestamp 1679235063
transform 1 0 5244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_66
timestamp 1679235063
transform 1 0 7176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_78
timestamp 1679235063
transform 1 0 8280 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_87
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_111
timestamp 1679235063
transform 1 0 11316 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_117
timestamp 1679235063
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_125
timestamp 1679235063
transform 1 0 12604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp 1679235063
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1679235063
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_175
timestamp 1679235063
transform 1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_179
timestamp 1679235063
transform 1 0 17572 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1679235063
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1679235063
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_202
timestamp 1679235063
transform 1 0 19688 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_226
timestamp 1679235063
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1679235063
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_10
timestamp 1679235063
transform 1 0 2024 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_35
timestamp 1679235063
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 1679235063
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1679235063
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_59
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_67
timestamp 1679235063
transform 1 0 7268 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_78
timestamp 1679235063
transform 1 0 8280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_91
timestamp 1679235063
transform 1 0 9476 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_99
timestamp 1679235063
transform 1 0 10212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_115
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1679235063
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_124
timestamp 1679235063
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_135
timestamp 1679235063
transform 1 0 13524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_141
timestamp 1679235063
transform 1 0 14076 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_152
timestamp 1679235063
transform 1 0 15088 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_156
timestamp 1679235063
transform 1 0 15456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1679235063
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_180
timestamp 1679235063
transform 1 0 17664 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_184
timestamp 1679235063
transform 1 0 18032 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_207
timestamp 1679235063
transform 1 0 20148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1679235063
transform 1 0 21252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1679235063
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_260
timestamp 1679235063
transform 1 0 25024 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_264
timestamp 1679235063
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1679235063
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_55
timestamp 1679235063
transform 1 0 6164 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_68
timestamp 1679235063
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1679235063
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1679235063
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_116
timestamp 1679235063
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_120
timestamp 1679235063
transform 1 0 12144 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1679235063
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1679235063
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_152
timestamp 1679235063
transform 1 0 15088 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_162
timestamp 1679235063
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_175
timestamp 1679235063
transform 1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1679235063
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_202
timestamp 1679235063
transform 1 0 19688 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1679235063
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1679235063
transform 1 0 23184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_248
timestamp 1679235063
transform 1 0 23920 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_263
timestamp 1679235063
transform 1 0 25300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1679235063
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_27
timestamp 1679235063
transform 1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_33
timestamp 1679235063
transform 1 0 4140 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1679235063
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_65
timestamp 1679235063
transform 1 0 7084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_76
timestamp 1679235063
transform 1 0 8096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_91
timestamp 1679235063
transform 1 0 9476 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_95
timestamp 1679235063
transform 1 0 9844 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_103
timestamp 1679235063
transform 1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1679235063
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1679235063
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_125
timestamp 1679235063
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_147
timestamp 1679235063
transform 1 0 14628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 1679235063
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_174
timestamp 1679235063
transform 1 0 17112 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_200
timestamp 1679235063
transform 1 0 19504 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1679235063
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1679235063
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_251
timestamp 1679235063
transform 1 0 24196 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_255
timestamp 1679235063
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_263
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_37
timestamp 1679235063
transform 1 0 4508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_45
timestamp 1679235063
transform 1 0 5244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_56
timestamp 1679235063
transform 1 0 6256 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_80
timestamp 1679235063
transform 1 0 8464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1679235063
transform 1 0 9476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_101
timestamp 1679235063
transform 1 0 10396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_108
timestamp 1679235063
transform 1 0 11040 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_115
timestamp 1679235063
transform 1 0 11684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_128
timestamp 1679235063
transform 1 0 12880 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1679235063
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_152
timestamp 1679235063
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_156
timestamp 1679235063
transform 1 0 15456 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_168
timestamp 1679235063
transform 1 0 16560 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_173
timestamp 1679235063
transform 1 0 17020 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1679235063
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1679235063
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_207
timestamp 1679235063
transform 1 0 20148 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1679235063
transform 1 0 20516 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_217
timestamp 1679235063
transform 1 0 21068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1679235063
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_263
timestamp 1679235063
transform 1 0 25300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1679235063
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_27
timestamp 1679235063
transform 1 0 3588 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_31
timestamp 1679235063
transform 1 0 3956 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_35
timestamp 1679235063
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1679235063
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1679235063
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_65
timestamp 1679235063
transform 1 0 7084 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_68
timestamp 1679235063
transform 1 0 7360 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_80
timestamp 1679235063
transform 1 0 8464 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_88
timestamp 1679235063
transform 1 0 9200 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_92
timestamp 1679235063
transform 1 0 9568 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1679235063
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1679235063
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_139
timestamp 1679235063
transform 1 0 13892 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_151
timestamp 1679235063
transform 1 0 14996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_155
timestamp 1679235063
transform 1 0 15364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1679235063
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_187
timestamp 1679235063
transform 1 0 18308 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_195
timestamp 1679235063
transform 1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_218
timestamp 1679235063
transform 1 0 21160 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1679235063
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_257
timestamp 1679235063
transform 1 0 24748 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_265
timestamp 1679235063
transform 1 0 25484 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1679235063
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_13
timestamp 1679235063
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1679235063
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_33
timestamp 1679235063
transform 1 0 4140 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_42
timestamp 1679235063
transform 1 0 4968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_66
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1679235063
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_93
timestamp 1679235063
transform 1 0 9660 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_103
timestamp 1679235063
transform 1 0 10580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_107
timestamp 1679235063
transform 1 0 10948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_111
timestamp 1679235063
transform 1 0 11316 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1679235063
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_153
timestamp 1679235063
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1679235063
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_187
timestamp 1679235063
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1679235063
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_203
timestamp 1679235063
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_224
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_232
timestamp 1679235063
transform 1 0 22448 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_261
timestamp 1679235063
transform 1 0 25116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_265
timestamp 1679235063
transform 1 0 25484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1679235063
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_7
timestamp 1679235063
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_29
timestamp 1679235063
transform 1 0 3772 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_36
timestamp 1679235063
transform 1 0 4416 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_48
timestamp 1679235063
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_59
timestamp 1679235063
transform 1 0 6532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_73
timestamp 1679235063
transform 1 0 7820 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_81
timestamp 1679235063
transform 1 0 8556 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_86
timestamp 1679235063
transform 1 0 9016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1679235063
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1679235063
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1679235063
transform 1 0 12420 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_133
timestamp 1679235063
transform 1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1679235063
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_149
timestamp 1679235063
transform 1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1679235063
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_171
timestamp 1679235063
transform 1 0 16836 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1679235063
transform 1 0 19044 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_199
timestamp 1679235063
transform 1 0 19412 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_209
timestamp 1679235063
transform 1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1679235063
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1679235063
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_244
timestamp 1679235063
transform 1 0 23552 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1679235063
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1679235063
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_17
timestamp 1679235063
transform 1 0 2668 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1679235063
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_29
timestamp 1679235063
transform 1 0 3772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_35
timestamp 1679235063
transform 1 0 4324 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_56
timestamp 1679235063
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_68
timestamp 1679235063
transform 1 0 7360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_72
timestamp 1679235063
transform 1 0 7728 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1679235063
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1679235063
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_96
timestamp 1679235063
transform 1 0 9936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_100
timestamp 1679235063
transform 1 0 10304 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_112
timestamp 1679235063
transform 1 0 11408 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_118
timestamp 1679235063
transform 1 0 11960 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1679235063
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1679235063
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1679235063
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_154
timestamp 1679235063
transform 1 0 15272 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_158
timestamp 1679235063
transform 1 0 15640 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_167
timestamp 1679235063
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_180
timestamp 1679235063
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_187
timestamp 1679235063
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1679235063
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1679235063
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1679235063
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_221
timestamp 1679235063
transform 1 0 21436 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_238
timestamp 1679235063
transform 1 0 23000 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1679235063
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1679235063
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_259
timestamp 1679235063
transform 1 0 24932 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_265
timestamp 1679235063
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1679235063
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_15
timestamp 1679235063
transform 1 0 2484 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_21
timestamp 1679235063
transform 1 0 3036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_25
timestamp 1679235063
transform 1 0 3404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_49
timestamp 1679235063
transform 1 0 5612 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1679235063
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1679235063
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_69
timestamp 1679235063
transform 1 0 7452 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_73
timestamp 1679235063
transform 1 0 7820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1679235063
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1679235063
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1679235063
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1679235063
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_121
timestamp 1679235063
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_134
timestamp 1679235063
transform 1 0 13432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_142
timestamp 1679235063
transform 1 0 14168 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1679235063
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_171
timestamp 1679235063
transform 1 0 16836 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_179
timestamp 1679235063
transform 1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_191
timestamp 1679235063
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_206
timestamp 1679235063
transform 1 0 20056 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_212
timestamp 1679235063
transform 1 0 20608 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_218
timestamp 1679235063
transform 1 0 21160 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1679235063
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_227
timestamp 1679235063
transform 1 0 21988 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_234
timestamp 1679235063
transform 1 0 22632 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_258
timestamp 1679235063
transform 1 0 24840 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1679235063
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1679235063
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1679235063
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_31
timestamp 1679235063
transform 1 0 3956 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_39
timestamp 1679235063
transform 1 0 4692 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_49
timestamp 1679235063
transform 1 0 5612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_61
timestamp 1679235063
transform 1 0 6716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1679235063
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1679235063
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_97
timestamp 1679235063
transform 1 0 10028 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1679235063
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_115
timestamp 1679235063
transform 1 0 11684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_127
timestamp 1679235063
transform 1 0 12788 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1679235063
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1679235063
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1679235063
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_165
timestamp 1679235063
transform 1 0 16284 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1679235063
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_179
timestamp 1679235063
transform 1 0 17572 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_184
timestamp 1679235063
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_197
timestamp 1679235063
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_207
timestamp 1679235063
transform 1 0 20148 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_229
timestamp 1679235063
transform 1 0 22172 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_242
timestamp 1679235063
transform 1 0 23368 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1679235063
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1679235063
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_259
timestamp 1679235063
transform 1 0 24932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_265
timestamp 1679235063
transform 1 0 25484 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1679235063
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_15
timestamp 1679235063
transform 1 0 2484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_23
timestamp 1679235063
transform 1 0 3220 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_27
timestamp 1679235063
transform 1 0 3588 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_38
timestamp 1679235063
transform 1 0 4600 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_50
timestamp 1679235063
transform 1 0 5704 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1679235063
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_79
timestamp 1679235063
transform 1 0 8372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_87
timestamp 1679235063
transform 1 0 9108 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_98
timestamp 1679235063
transform 1 0 10120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_105
timestamp 1679235063
transform 1 0 10764 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1679235063
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1679235063
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_118
timestamp 1679235063
transform 1 0 11960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1679235063
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_163
timestamp 1679235063
transform 1 0 16100 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1679235063
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1679235063
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_180
timestamp 1679235063
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_193
timestamp 1679235063
transform 1 0 18860 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_199
timestamp 1679235063
transform 1 0 19412 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_203
timestamp 1679235063
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_216
timestamp 1679235063
transform 1 0 20976 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1679235063
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_236
timestamp 1679235063
transform 1 0 22816 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_248
timestamp 1679235063
transform 1 0 23920 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_260
timestamp 1679235063
transform 1 0 25024 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1679235063
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1679235063
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1679235063
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1679235063
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_52
timestamp 1679235063
transform 1 0 5888 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_60
timestamp 1679235063
transform 1 0 6624 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_70
timestamp 1679235063
transform 1 0 7544 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1679235063
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1679235063
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_109
timestamp 1679235063
transform 1 0 11132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_113
timestamp 1679235063
transform 1 0 11500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_123
timestamp 1679235063
transform 1 0 12420 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1679235063
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_145
timestamp 1679235063
transform 1 0 14444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_149
timestamp 1679235063
transform 1 0 14812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1679235063
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_187
timestamp 1679235063
transform 1 0 18308 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1679235063
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1679235063
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_208
timestamp 1679235063
transform 1 0 20240 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_212
timestamp 1679235063
transform 1 0 20608 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_218
timestamp 1679235063
transform 1 0 21160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_243
timestamp 1679235063
transform 1 0 23460 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1679235063
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1679235063
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_263
timestamp 1679235063
transform 1 0 25300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1679235063
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1679235063
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1679235063
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1679235063
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1679235063
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1679235063
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1679235063
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_61
timestamp 1679235063
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_82
timestamp 1679235063
transform 1 0 8648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_106
timestamp 1679235063
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1679235063
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_123
timestamp 1679235063
transform 1 0 12420 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_147
timestamp 1679235063
transform 1 0 14628 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1679235063
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1679235063
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1679235063
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_176
timestamp 1679235063
transform 1 0 17296 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_187
timestamp 1679235063
transform 1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_191
timestamp 1679235063
transform 1 0 18676 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_197
timestamp 1679235063
transform 1 0 19228 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_208
timestamp 1679235063
transform 1 0 20240 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1679235063
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1679235063
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_248
timestamp 1679235063
transform 1 0 23920 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_254
timestamp 1679235063
transform 1 0 24472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1679235063
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_265
timestamp 1679235063
transform 1 0 25484 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1679235063
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1679235063
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1679235063
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1679235063
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_33
timestamp 1679235063
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_55
timestamp 1679235063
transform 1 0 6164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_61
timestamp 1679235063
transform 1 0 6716 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1679235063
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1679235063
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_95
timestamp 1679235063
transform 1 0 9844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_107
timestamp 1679235063
transform 1 0 10948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_113
timestamp 1679235063
transform 1 0 11500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_117
timestamp 1679235063
transform 1 0 11868 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_130
timestamp 1679235063
transform 1 0 13064 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1679235063
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1679235063
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_152
timestamp 1679235063
transform 1 0 15088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_158
timestamp 1679235063
transform 1 0 15640 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_175
timestamp 1679235063
transform 1 0 17204 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_188
timestamp 1679235063
transform 1 0 18400 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1679235063
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_219
timestamp 1679235063
transform 1 0 21252 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_223
timestamp 1679235063
transform 1 0 21620 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_229
timestamp 1679235063
transform 1 0 22172 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1679235063
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1679235063
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_259
timestamp 1679235063
transform 1 0 24932 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_265
timestamp 1679235063
transform 1 0 25484 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1679235063
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_15
timestamp 1679235063
transform 1 0 2484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_23
timestamp 1679235063
transform 1 0 3220 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_28
timestamp 1679235063
transform 1 0 3680 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_40
timestamp 1679235063
transform 1 0 4784 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1679235063
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_57
timestamp 1679235063
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_63
timestamp 1679235063
transform 1 0 6900 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_72
timestamp 1679235063
transform 1 0 7728 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_77
timestamp 1679235063
transform 1 0 8188 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_88
timestamp 1679235063
transform 1 0 9200 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_92
timestamp 1679235063
transform 1 0 9568 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_101
timestamp 1679235063
transform 1 0 10396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1679235063
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1679235063
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_116
timestamp 1679235063
transform 1 0 11776 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_127
timestamp 1679235063
transform 1 0 12788 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_133
timestamp 1679235063
transform 1 0 13340 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_143
timestamp 1679235063
transform 1 0 14260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1679235063
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_171
timestamp 1679235063
transform 1 0 16836 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_177
timestamp 1679235063
transform 1 0 17388 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_187
timestamp 1679235063
transform 1 0 18308 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_200
timestamp 1679235063
transform 1 0 19504 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_212
timestamp 1679235063
transform 1 0 20608 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_218
timestamp 1679235063
transform 1 0 21160 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1679235063
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1679235063
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_235
timestamp 1679235063
transform 1 0 22724 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_242
timestamp 1679235063
transform 1 0 23368 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_249
timestamp 1679235063
transform 1 0 24012 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_253
timestamp 1679235063
transform 1 0 24380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_259
timestamp 1679235063
transform 1 0 24932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_265
timestamp 1679235063
transform 1 0 25484 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1679235063
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1679235063
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1679235063
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_29
timestamp 1679235063
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1679235063
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_65
timestamp 1679235063
transform 1 0 7084 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_73
timestamp 1679235063
transform 1 0 7820 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1679235063
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1679235063
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1679235063
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_93
timestamp 1679235063
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_114
timestamp 1679235063
transform 1 0 11592 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_118
timestamp 1679235063
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_130
timestamp 1679235063
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1679235063
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1679235063
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1679235063
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1679235063
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_192
timestamp 1679235063
transform 1 0 18768 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_197
timestamp 1679235063
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_209
timestamp 1679235063
transform 1 0 20332 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_217
timestamp 1679235063
transform 1 0 21068 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_228
timestamp 1679235063
transform 1 0 22080 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_241
timestamp 1679235063
transform 1 0 23276 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_245
timestamp 1679235063
transform 1 0 23644 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1679235063
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1679235063
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_258
timestamp 1679235063
transform 1 0 24840 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_262
timestamp 1679235063
transform 1 0 25208 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1679235063
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1679235063
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1679235063
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1679235063
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1679235063
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1679235063
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1679235063
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1679235063
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_81
timestamp 1679235063
transform 1 0 8556 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_86
timestamp 1679235063
transform 1 0 9016 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_97
timestamp 1679235063
transform 1 0 10028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1679235063
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_117
timestamp 1679235063
transform 1 0 11868 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_123
timestamp 1679235063
transform 1 0 12420 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_134
timestamp 1679235063
transform 1 0 13432 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_146
timestamp 1679235063
transform 1 0 14536 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1679235063
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1679235063
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_171
timestamp 1679235063
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_175
timestamp 1679235063
transform 1 0 17204 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_186
timestamp 1679235063
transform 1 0 18216 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_190
timestamp 1679235063
transform 1 0 18584 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1679235063
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_211
timestamp 1679235063
transform 1 0 20516 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_218
timestamp 1679235063
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_225
timestamp 1679235063
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_233
timestamp 1679235063
transform 1 0 22540 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_236
timestamp 1679235063
transform 1 0 22816 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_241
timestamp 1679235063
transform 1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_248
timestamp 1679235063
transform 1 0 23920 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_252
timestamp 1679235063
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_264
timestamp 1679235063
transform 1 0 25392 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1679235063
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1679235063
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1679235063
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1679235063
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1679235063
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1679235063
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_65
timestamp 1679235063
transform 1 0 7084 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_69
timestamp 1679235063
transform 1 0 7452 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp 1679235063
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1679235063
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1679235063
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_113
timestamp 1679235063
transform 1 0 11500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_120
timestamp 1679235063
transform 1 0 12144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_124
timestamp 1679235063
transform 1 0 12512 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_134
timestamp 1679235063
transform 1 0 13432 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1679235063
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1679235063
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_152
timestamp 1679235063
transform 1 0 15088 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_158
timestamp 1679235063
transform 1 0 15640 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_169
timestamp 1679235063
transform 1 0 16652 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_173
timestamp 1679235063
transform 1 0 17020 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1679235063
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_197
timestamp 1679235063
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1679235063
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_216
timestamp 1679235063
transform 1 0 20976 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_220
timestamp 1679235063
transform 1 0 21344 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_224
timestamp 1679235063
transform 1 0 21712 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_228
timestamp 1679235063
transform 1 0 22080 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_236
timestamp 1679235063
transform 1 0 22816 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1679235063
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1679235063
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_258
timestamp 1679235063
transform 1 0 24840 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1679235063
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1679235063
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_27
timestamp 1679235063
transform 1 0 3588 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1679235063
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_57
timestamp 1679235063
transform 1 0 6348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_67
timestamp 1679235063
transform 1 0 7268 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_78
timestamp 1679235063
transform 1 0 8280 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_90
timestamp 1679235063
transform 1 0 9384 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1679235063
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1679235063
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_145
timestamp 1679235063
transform 1 0 14444 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_158
timestamp 1679235063
transform 1 0 15640 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1679235063
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1679235063
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_180
timestamp 1679235063
transform 1 0 17664 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_186
timestamp 1679235063
transform 1 0 18216 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1679235063
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_209
timestamp 1679235063
transform 1 0 20332 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1679235063
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1679235063
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_236
timestamp 1679235063
transform 1 0 22816 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_240
timestamp 1679235063
transform 1 0 23184 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_263
timestamp 1679235063
transform 1 0 25300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1679235063
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1679235063
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1679235063
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1679235063
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1679235063
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_53
timestamp 1679235063
transform 1 0 5980 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_59
timestamp 1679235063
transform 1 0 6532 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_80
timestamp 1679235063
transform 1 0 8464 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1679235063
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_90
timestamp 1679235063
transform 1 0 9384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_94
timestamp 1679235063
transform 1 0 9752 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_115
timestamp 1679235063
transform 1 0 11684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_119
timestamp 1679235063
transform 1 0 12052 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_130
timestamp 1679235063
transform 1 0 13064 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1679235063
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_152
timestamp 1679235063
transform 1 0 15088 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_176
timestamp 1679235063
transform 1 0 17296 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1679235063
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_197
timestamp 1679235063
transform 1 0 19228 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_200
timestamp 1679235063
transform 1 0 19504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_205
timestamp 1679235063
transform 1 0 19964 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_213
timestamp 1679235063
transform 1 0 20700 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_224
timestamp 1679235063
transform 1 0 21712 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_228
timestamp 1679235063
transform 1 0 22080 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1679235063
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1679235063
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_263
timestamp 1679235063
transform 1 0 25300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1679235063
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1679235063
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1679235063
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1679235063
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1679235063
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1679235063
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1679235063
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_65
timestamp 1679235063
transform 1 0 7084 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_71
timestamp 1679235063
transform 1 0 7636 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_96
timestamp 1679235063
transform 1 0 9936 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_100
timestamp 1679235063
transform 1 0 10304 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1679235063
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_117
timestamp 1679235063
transform 1 0 11868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_120
timestamp 1679235063
transform 1 0 12144 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_131
timestamp 1679235063
transform 1 0 13156 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_139
timestamp 1679235063
transform 1 0 13892 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_150
timestamp 1679235063
transform 1 0 14904 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_162
timestamp 1679235063
transform 1 0 16008 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_169
timestamp 1679235063
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_177
timestamp 1679235063
transform 1 0 17388 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_188
timestamp 1679235063
transform 1 0 18400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_201
timestamp 1679235063
transform 1 0 19596 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1679235063
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_218
timestamp 1679235063
transform 1 0 21160 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1679235063
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1679235063
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_237
timestamp 1679235063
transform 1 0 22908 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_251
timestamp 1679235063
transform 1 0 24196 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1679235063
transform 1 0 25392 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1679235063
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1679235063
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1679235063
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1679235063
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 1679235063
transform 1 0 4876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_49
timestamp 1679235063
transform 1 0 5612 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_71
timestamp 1679235063
transform 1 0 7636 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_75
timestamp 1679235063
transform 1 0 8004 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1679235063
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1679235063
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_95
timestamp 1679235063
transform 1 0 9844 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_107
timestamp 1679235063
transform 1 0 10948 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_119
timestamp 1679235063
transform 1 0 12052 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_131
timestamp 1679235063
transform 1 0 13156 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1679235063
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1679235063
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_163
timestamp 1679235063
transform 1 0 16100 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_168
timestamp 1679235063
transform 1 0 16560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_179
timestamp 1679235063
transform 1 0 17572 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_183
timestamp 1679235063
transform 1 0 17940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1679235063
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_197
timestamp 1679235063
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_206
timestamp 1679235063
transform 1 0 20056 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_213
timestamp 1679235063
transform 1 0 20700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_217
timestamp 1679235063
transform 1 0 21068 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_227
timestamp 1679235063
transform 1 0 21988 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_234
timestamp 1679235063
transform 1 0 22632 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_241
timestamp 1679235063
transform 1 0 23276 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_245
timestamp 1679235063
transform 1 0 23644 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1679235063
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_259
timestamp 1679235063
transform 1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1679235063
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1679235063
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_8
timestamp 1679235063
transform 1 0 1840 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_12
timestamp 1679235063
transform 1 0 2208 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_24
timestamp 1679235063
transform 1 0 3312 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_36
timestamp 1679235063
transform 1 0 4416 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_48
timestamp 1679235063
transform 1 0 5520 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1679235063
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 1679235063
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_73
timestamp 1679235063
transform 1 0 7820 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_84
timestamp 1679235063
transform 1 0 8832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_88
timestamp 1679235063
transform 1 0 9200 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_103
timestamp 1679235063
transform 1 0 10580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1679235063
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1679235063
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_124
timestamp 1679235063
transform 1 0 12512 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_136
timestamp 1679235063
transform 1 0 13616 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_140
timestamp 1679235063
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_143
timestamp 1679235063
transform 1 0 14260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_153
timestamp 1679235063
transform 1 0 15180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1679235063
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1679235063
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_181
timestamp 1679235063
transform 1 0 17756 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_204
timestamp 1679235063
transform 1 0 19872 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_218
timestamp 1679235063
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1679235063
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_236
timestamp 1679235063
transform 1 0 22816 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_240
timestamp 1679235063
transform 1 0 23184 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1679235063
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1679235063
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1679235063
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1679235063
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1679235063
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_41
timestamp 1679235063
transform 1 0 4876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_49
timestamp 1679235063
transform 1 0 5612 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_54
timestamp 1679235063
transform 1 0 6072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_66
timestamp 1679235063
transform 1 0 7176 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1679235063
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1679235063
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1679235063
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_104
timestamp 1679235063
transform 1 0 10672 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_117
timestamp 1679235063
transform 1 0 11868 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1679235063
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1679235063
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_152
timestamp 1679235063
transform 1 0 15088 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_156
timestamp 1679235063
transform 1 0 15456 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1679235063
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1679235063
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1679235063
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_199
timestamp 1679235063
transform 1 0 19412 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_210
timestamp 1679235063
transform 1 0 20424 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1679235063
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_235
timestamp 1679235063
transform 1 0 22724 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_242
timestamp 1679235063
transform 1 0 23368 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_246
timestamp 1679235063
transform 1 0 23736 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1679235063
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_255
timestamp 1679235063
transform 1 0 24564 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_259
timestamp 1679235063
transform 1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_264
timestamp 1679235063
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1679235063
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1679235063
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1679235063
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_39
timestamp 1679235063
transform 1 0 4692 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_43
timestamp 1679235063
transform 1 0 5060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1679235063
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1679235063
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_80
timestamp 1679235063
transform 1 0 8464 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_104
timestamp 1679235063
transform 1 0 10672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1679235063
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_135
timestamp 1679235063
transform 1 0 13524 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_148
timestamp 1679235063
transform 1 0 14720 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_160
timestamp 1679235063
transform 1 0 15824 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_169
timestamp 1679235063
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_183
timestamp 1679235063
transform 1 0 17940 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_196
timestamp 1679235063
transform 1 0 19136 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_202
timestamp 1679235063
transform 1 0 19688 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_213
timestamp 1679235063
transform 1 0 20700 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1679235063
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1679235063
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_227
timestamp 1679235063
transform 1 0 21988 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_238
timestamp 1679235063
transform 1 0 23000 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_242
timestamp 1679235063
transform 1 0 23368 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_249
timestamp 1679235063
transform 1 0 24012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1679235063
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_260
timestamp 1679235063
transform 1 0 25024 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1679235063
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1679235063
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1679235063
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1679235063
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1679235063
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_41
timestamp 1679235063
transform 1 0 4876 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_47
timestamp 1679235063
transform 1 0 5428 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_68
timestamp 1679235063
transform 1 0 7360 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_72
timestamp 1679235063
transform 1 0 7728 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1679235063
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_87
timestamp 1679235063
transform 1 0 9108 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_98
timestamp 1679235063
transform 1 0 10120 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_102
timestamp 1679235063
transform 1 0 10488 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_123
timestamp 1679235063
transform 1 0 12420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_127
timestamp 1679235063
transform 1 0 12788 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1679235063
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_143
timestamp 1679235063
transform 1 0 14260 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_155
timestamp 1679235063
transform 1 0 15364 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_176
timestamp 1679235063
transform 1 0 17296 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_184
timestamp 1679235063
transform 1 0 18032 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1679235063
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1679235063
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_219
timestamp 1679235063
transform 1 0 21252 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_236
timestamp 1679235063
transform 1 0 22816 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_249
timestamp 1679235063
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1679235063
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_263
timestamp 1679235063
transform 1 0 25300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1679235063
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1679235063
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_27
timestamp 1679235063
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_33
timestamp 1679235063
transform 1 0 4140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1679235063
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_59
timestamp 1679235063
transform 1 0 6532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_63
timestamp 1679235063
transform 1 0 6900 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_66
timestamp 1679235063
transform 1 0 7176 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_76
timestamp 1679235063
transform 1 0 8096 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1679235063
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1679235063
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_135
timestamp 1679235063
transform 1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_139
timestamp 1679235063
transform 1 0 13892 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_151
timestamp 1679235063
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_163
timestamp 1679235063
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1679235063
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1679235063
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_181
timestamp 1679235063
transform 1 0 17756 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_202
timestamp 1679235063
transform 1 0 19688 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_214
timestamp 1679235063
transform 1 0 20792 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1679235063
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1679235063
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1679235063
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1679235063
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_260
timestamp 1679235063
transform 1 0 25024 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1679235063
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_8
timestamp 1679235063
transform 1 0 1840 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_12
timestamp 1679235063
transform 1 0 2208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1679235063
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1679235063
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1679235063
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_53
timestamp 1679235063
transform 1 0 5980 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_59
timestamp 1679235063
transform 1 0 6532 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1679235063
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_85
timestamp 1679235063
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_100
timestamp 1679235063
transform 1 0 10304 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_108
timestamp 1679235063
transform 1 0 11040 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_119
timestamp 1679235063
transform 1 0 12052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_132
timestamp 1679235063
transform 1 0 13248 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1679235063
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_152
timestamp 1679235063
transform 1 0 15088 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_159
timestamp 1679235063
transform 1 0 15732 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_171
timestamp 1679235063
transform 1 0 16836 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_174
timestamp 1679235063
transform 1 0 17112 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_186
timestamp 1679235063
transform 1 0 18216 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1679235063
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1679235063
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_208
timestamp 1679235063
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_223
timestamp 1679235063
transform 1 0 21620 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_229
timestamp 1679235063
transform 1 0 22172 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1679235063
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1679235063
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1679235063
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1679235063
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1679235063
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1679235063
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1679235063
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1679235063
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1679235063
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1679235063
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_89
timestamp 1679235063
transform 1 0 9292 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_93
timestamp 1679235063
transform 1 0 9660 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1679235063
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_115
timestamp 1679235063
transform 1 0 11684 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_123
timestamp 1679235063
transform 1 0 12420 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_134
timestamp 1679235063
transform 1 0 13432 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_138
timestamp 1679235063
transform 1 0 13800 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_146
timestamp 1679235063
transform 1 0 14536 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_156
timestamp 1679235063
transform 1 0 15456 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_160
timestamp 1679235063
transform 1 0 15824 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_163
timestamp 1679235063
transform 1 0 16100 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1679235063
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_180
timestamp 1679235063
transform 1 0 17664 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_192
timestamp 1679235063
transform 1 0 18768 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1679235063
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_207
timestamp 1679235063
transform 1 0 20148 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_217
timestamp 1679235063
transform 1 0 21068 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1679235063
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1679235063
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_236
timestamp 1679235063
transform 1 0 22816 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_242
timestamp 1679235063
transform 1 0 23368 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1679235063
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1679235063
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1679235063
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1679235063
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1679235063
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1679235063
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1679235063
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_65
timestamp 1679235063
transform 1 0 7084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_78
timestamp 1679235063
transform 1 0 8280 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1679235063
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_98
timestamp 1679235063
transform 1 0 10120 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_111
timestamp 1679235063
transform 1 0 11316 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1679235063
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1679235063
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_143
timestamp 1679235063
transform 1 0 14260 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_146
timestamp 1679235063
transform 1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_157
timestamp 1679235063
transform 1 0 15548 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_161
timestamp 1679235063
transform 1 0 15916 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1679235063
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_179
timestamp 1679235063
transform 1 0 17572 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_183
timestamp 1679235063
transform 1 0 17940 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1679235063
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1679235063
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_210
timestamp 1679235063
transform 1 0 20424 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_218
timestamp 1679235063
transform 1 0 21160 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_232
timestamp 1679235063
transform 1 0 22448 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_244
timestamp 1679235063
transform 1 0 23552 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1679235063
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_263
timestamp 1679235063
transform 1 0 25300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1679235063
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1679235063
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_27
timestamp 1679235063
transform 1 0 3588 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_33
timestamp 1679235063
transform 1 0 4140 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1679235063
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1679235063
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_82
timestamp 1679235063
transform 1 0 8648 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_86
timestamp 1679235063
transform 1 0 9016 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_90
timestamp 1679235063
transform 1 0 9384 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_100
timestamp 1679235063
transform 1 0 10304 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_104
timestamp 1679235063
transform 1 0 10672 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1679235063
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_124
timestamp 1679235063
transform 1 0 12512 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_136
timestamp 1679235063
transform 1 0 13616 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_143
timestamp 1679235063
transform 1 0 14260 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_148
timestamp 1679235063
transform 1 0 14720 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_159
timestamp 1679235063
transform 1 0 15732 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1679235063
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1679235063
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_191
timestamp 1679235063
transform 1 0 18676 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_204
timestamp 1679235063
transform 1 0 19872 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_217
timestamp 1679235063
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1679235063
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1679235063
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_230
timestamp 1679235063
transform 1 0 22264 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_254
timestamp 1679235063
transform 1 0 24472 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_258
timestamp 1679235063
transform 1 0 24840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1679235063
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1679235063
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_8
timestamp 1679235063
transform 1 0 1840 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_12
timestamp 1679235063
transform 1 0 2208 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1679235063
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1679235063
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_41
timestamp 1679235063
transform 1 0 4876 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_69
timestamp 1679235063
transform 1 0 7452 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_81
timestamp 1679235063
transform 1 0 8556 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_85
timestamp 1679235063
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_92
timestamp 1679235063
transform 1 0 9568 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_103
timestamp 1679235063
transform 1 0 10580 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_116
timestamp 1679235063
transform 1 0 11776 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_124
timestamp 1679235063
transform 1 0 12512 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_135
timestamp 1679235063
transform 1 0 13524 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1679235063
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_141
timestamp 1679235063
transform 1 0 14076 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_149
timestamp 1679235063
transform 1 0 14812 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_160
timestamp 1679235063
transform 1 0 15824 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_173
timestamp 1679235063
transform 1 0 17020 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_186
timestamp 1679235063
transform 1 0 18216 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_190
timestamp 1679235063
transform 1 0 18584 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_193
timestamp 1679235063
transform 1 0 18860 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1679235063
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_208
timestamp 1679235063
transform 1 0 20240 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_212
timestamp 1679235063
transform 1 0 20608 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_216
timestamp 1679235063
transform 1 0 20976 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_221
timestamp 1679235063
transform 1 0 21436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_234
timestamp 1679235063
transform 1 0 22632 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_247
timestamp 1679235063
transform 1 0 23828 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1679235063
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1679235063
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_263
timestamp 1679235063
transform 1 0 25300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1679235063
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1679235063
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1679235063
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_39
timestamp 1679235063
transform 1 0 4692 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_45
timestamp 1679235063
transform 1 0 5244 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1679235063
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 1679235063
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_68
timestamp 1679235063
transform 1 0 7360 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_74
timestamp 1679235063
transform 1 0 7912 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_77
timestamp 1679235063
transform 1 0 8188 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_88
timestamp 1679235063
transform 1 0 9200 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_97
timestamp 1679235063
transform 1 0 10028 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1679235063
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_113
timestamp 1679235063
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_118
timestamp 1679235063
transform 1 0 11960 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_122
timestamp 1679235063
transform 1 0 12328 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_143
timestamp 1679235063
transform 1 0 14260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_147
timestamp 1679235063
transform 1 0 14628 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_160
timestamp 1679235063
transform 1 0 15824 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1679235063
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_169
timestamp 1679235063
transform 1 0 16652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_175
timestamp 1679235063
transform 1 0 17204 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_186
timestamp 1679235063
transform 1 0 18216 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_190
timestamp 1679235063
transform 1 0 18584 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_202
timestamp 1679235063
transform 1 0 19688 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_215
timestamp 1679235063
transform 1 0 20884 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1679235063
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1679235063
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_236
timestamp 1679235063
transform 1 0 22816 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_249
timestamp 1679235063
transform 1 0 24012 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_264
timestamp 1679235063
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1679235063
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1679235063
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1679235063
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1679235063
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_41
timestamp 1679235063
transform 1 0 4876 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_67
timestamp 1679235063
transform 1 0 7268 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_71
timestamp 1679235063
transform 1 0 7636 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_82
timestamp 1679235063
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1679235063
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_96
timestamp 1679235063
transform 1 0 9936 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_100
timestamp 1679235063
transform 1 0 10304 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_103
timestamp 1679235063
transform 1 0 10580 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_114
timestamp 1679235063
transform 1 0 11592 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_118
timestamp 1679235063
transform 1 0 11960 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_130
timestamp 1679235063
transform 1 0 13064 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_134
timestamp 1679235063
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_141
timestamp 1679235063
transform 1 0 14076 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_149
timestamp 1679235063
transform 1 0 14812 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_161
timestamp 1679235063
transform 1 0 15916 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_165
timestamp 1679235063
transform 1 0 16284 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_175
timestamp 1679235063
transform 1 0 17204 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_189
timestamp 1679235063
transform 1 0 18492 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1679235063
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1679235063
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_202
timestamp 1679235063
transform 1 0 19688 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_206
timestamp 1679235063
transform 1 0 20056 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_216
timestamp 1679235063
transform 1 0 20976 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_224
timestamp 1679235063
transform 1 0 21712 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1679235063
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_253
timestamp 1679235063
transform 1 0 24380 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1679235063
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1679235063
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1679235063
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1679235063
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1679235063
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1679235063
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1679235063
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1679235063
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1679235063
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_81
timestamp 1679235063
transform 1 0 8556 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_107
timestamp 1679235063
transform 1 0 10948 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1679235063
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_135
timestamp 1679235063
transform 1 0 13524 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_139
timestamp 1679235063
transform 1 0 13892 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_144
timestamp 1679235063
transform 1 0 14352 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_155
timestamp 1679235063
transform 1 0 15364 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_162
timestamp 1679235063
transform 1 0 16008 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_166
timestamp 1679235063
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_169
timestamp 1679235063
transform 1 0 16652 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_180
timestamp 1679235063
transform 1 0 17664 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_187
timestamp 1679235063
transform 1 0 18308 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_195
timestamp 1679235063
transform 1 0 19044 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_206
timestamp 1679235063
transform 1 0 20056 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_210
timestamp 1679235063
transform 1 0 20424 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_225
timestamp 1679235063
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_236
timestamp 1679235063
transform 1 0 22816 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_240
timestamp 1679235063
transform 1 0 23184 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1679235063
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1679235063
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1679235063
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1679235063
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1679235063
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1679235063
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1679235063
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_65
timestamp 1679235063
transform 1 0 7084 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_71
timestamp 1679235063
transform 1 0 7636 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_80
timestamp 1679235063
transform 1 0 8464 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_85
timestamp 1679235063
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_97
timestamp 1679235063
transform 1 0 10028 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_110
timestamp 1679235063
transform 1 0 11224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_123
timestamp 1679235063
transform 1 0 12420 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_136
timestamp 1679235063
transform 1 0 13616 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_141
timestamp 1679235063
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_156
timestamp 1679235063
transform 1 0 15456 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_169
timestamp 1679235063
transform 1 0 16652 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_173
timestamp 1679235063
transform 1 0 17020 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 1679235063
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 1679235063
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_205
timestamp 1679235063
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_210
timestamp 1679235063
transform 1 0 20424 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_222
timestamp 1679235063
transform 1 0 21528 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_229
timestamp 1679235063
transform 1 0 22172 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_242
timestamp 1679235063
transform 1 0 23368 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_246
timestamp 1679235063
transform 1 0 23736 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1679235063
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1679235063
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_263
timestamp 1679235063
transform 1 0 25300 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1679235063
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_8
timestamp 1679235063
transform 1 0 1840 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_12
timestamp 1679235063
transform 1 0 2208 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_24
timestamp 1679235063
transform 1 0 3312 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_36
timestamp 1679235063
transform 1 0 4416 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_48
timestamp 1679235063
transform 1 0 5520 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_57
timestamp 1679235063
transform 1 0 6348 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_80
timestamp 1679235063
transform 1 0 8464 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_88
timestamp 1679235063
transform 1 0 9200 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_92
timestamp 1679235063
transform 1 0 9568 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_104
timestamp 1679235063
transform 1 0 10672 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1679235063
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_124
timestamp 1679235063
transform 1 0 12512 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_128
timestamp 1679235063
transform 1 0 12880 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_152
timestamp 1679235063
transform 1 0 15088 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_165
timestamp 1679235063
transform 1 0 16284 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1679235063
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_180
timestamp 1679235063
transform 1 0 17664 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_184
timestamp 1679235063
transform 1 0 18032 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_195
timestamp 1679235063
transform 1 0 19044 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_208
timestamp 1679235063
transform 1 0 20240 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_221
timestamp 1679235063
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_229
timestamp 1679235063
transform 1 0 22172 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_240
timestamp 1679235063
transform 1 0 23184 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_244
timestamp 1679235063
transform 1 0 23552 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_249
timestamp 1679235063
transform 1 0 24012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_253
timestamp 1679235063
transform 1 0 24380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1679235063
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1679235063
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1679235063
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1679235063
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_29
timestamp 1679235063
transform 1 0 3772 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_33
timestamp 1679235063
transform 1 0 4140 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_41
timestamp 1679235063
transform 1 0 4876 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_45
timestamp 1679235063
transform 1 0 5244 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_53
timestamp 1679235063
transform 1 0 5980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_76
timestamp 1679235063
transform 1 0 8096 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_80
timestamp 1679235063
transform 1 0 8464 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_85
timestamp 1679235063
transform 1 0 8924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_89
timestamp 1679235063
transform 1 0 9292 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_110
timestamp 1679235063
transform 1 0 11224 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_114
timestamp 1679235063
transform 1 0 11592 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_118
timestamp 1679235063
transform 1 0 11960 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_130
timestamp 1679235063
transform 1 0 13064 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_134
timestamp 1679235063
transform 1 0 13432 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_141
timestamp 1679235063
transform 1 0 14076 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_163
timestamp 1679235063
transform 1 0 16100 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_176
timestamp 1679235063
transform 1 0 17296 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_188
timestamp 1679235063
transform 1 0 18400 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_192
timestamp 1679235063
transform 1 0 18768 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1679235063
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_210
timestamp 1679235063
transform 1 0 20424 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_217
timestamp 1679235063
transform 1 0 21068 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_232
timestamp 1679235063
transform 1 0 22448 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_245
timestamp 1679235063
transform 1 0 23644 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1679235063
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1679235063
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1679235063
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_15
timestamp 1679235063
transform 1 0 2484 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_23
timestamp 1679235063
transform 1 0 3220 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_29
timestamp 1679235063
transform 1 0 3772 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_37
timestamp 1679235063
transform 1 0 4508 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_45
timestamp 1679235063
transform 1 0 5244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1679235063
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1679235063
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1679235063
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_69
timestamp 1679235063
transform 1 0 7452 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_93
timestamp 1679235063
transform 1 0 9660 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1679235063
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1679235063
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_113
timestamp 1679235063
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_124
timestamp 1679235063
transform 1 0 12512 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_128
timestamp 1679235063
transform 1 0 12880 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_138
timestamp 1679235063
transform 1 0 13800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_150
timestamp 1679235063
transform 1 0 14904 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_154
timestamp 1679235063
transform 1 0 15272 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1679235063
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_169
timestamp 1679235063
transform 1 0 16652 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_172
timestamp 1679235063
transform 1 0 16928 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_183
timestamp 1679235063
transform 1 0 17940 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_189
timestamp 1679235063
transform 1 0 18492 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_211
timestamp 1679235063
transform 1 0 20516 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_217
timestamp 1679235063
transform 1 0 21068 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1679235063
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1679235063
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_230
timestamp 1679235063
transform 1 0 22264 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_234
timestamp 1679235063
transform 1 0 22632 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_257
timestamp 1679235063
transform 1 0 24748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_264
timestamp 1679235063
transform 1 0 25392 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1679235063
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1679235063
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1679235063
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 1679235063
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_37
timestamp 1679235063
transform 1 0 4508 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_43
timestamp 1679235063
transform 1 0 5060 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_47
timestamp 1679235063
transform 1 0 5428 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_54
timestamp 1679235063
transform 1 0 6072 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_58
timestamp 1679235063
transform 1 0 6440 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_70
timestamp 1679235063
transform 1 0 7544 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1679235063
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_85
timestamp 1679235063
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_96
timestamp 1679235063
transform 1 0 9936 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_100
timestamp 1679235063
transform 1 0 10304 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_104
timestamp 1679235063
transform 1 0 10672 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_128
timestamp 1679235063
transform 1 0 12880 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_132
timestamp 1679235063
transform 1 0 13248 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_136
timestamp 1679235063
transform 1 0 13616 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_141
timestamp 1679235063
transform 1 0 14076 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_149
timestamp 1679235063
transform 1 0 14812 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_170
timestamp 1679235063
transform 1 0 16744 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_183
timestamp 1679235063
transform 1 0 17940 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1679235063
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1679235063
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_197
timestamp 1679235063
transform 1 0 19228 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_210
timestamp 1679235063
transform 1 0 20424 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_225
timestamp 1679235063
transform 1 0 21804 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_229
timestamp 1679235063
transform 1 0 22172 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1679235063
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_253
timestamp 1679235063
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_263
timestamp 1679235063
transform 1 0 25300 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1679235063
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_9
timestamp 1679235063
transform 1 0 1932 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_13
timestamp 1679235063
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_25
timestamp 1679235063
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_37
timestamp 1679235063
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1679235063
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1679235063
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1679235063
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_69
timestamp 1679235063
transform 1 0 7452 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_73
timestamp 1679235063
transform 1 0 7820 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_77
timestamp 1679235063
transform 1 0 8188 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_102
timestamp 1679235063
transform 1 0 10488 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_106
timestamp 1679235063
transform 1 0 10856 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1679235063
transform 1 0 11224 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1679235063
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_125
timestamp 1679235063
transform 1 0 12604 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_147
timestamp 1679235063
transform 1 0 14628 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_160
timestamp 1679235063
transform 1 0 15824 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1679235063
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_169
timestamp 1679235063
transform 1 0 16652 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_181
timestamp 1679235063
transform 1 0 17756 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_205
timestamp 1679235063
transform 1 0 19964 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_217
timestamp 1679235063
transform 1 0 21068 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1679235063
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_236
timestamp 1679235063
transform 1 0 22816 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_240
timestamp 1679235063
transform 1 0 23184 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_263
timestamp 1679235063
transform 1 0 25300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1679235063
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1679235063
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1679235063
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1679235063
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1679235063
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1679235063
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_65
timestamp 1679235063
transform 1 0 7084 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_73
timestamp 1679235063
transform 1 0 7820 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_77
timestamp 1679235063
transform 1 0 8188 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1679235063
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_85
timestamp 1679235063
transform 1 0 8924 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_97
timestamp 1679235063
transform 1 0 10028 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_101
timestamp 1679235063
transform 1 0 10396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_113
timestamp 1679235063
transform 1 0 11500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_117
timestamp 1679235063
transform 1 0 11868 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_127
timestamp 1679235063
transform 1 0 12788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1679235063
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_141
timestamp 1679235063
transform 1 0 14076 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_151
timestamp 1679235063
transform 1 0 14996 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_164
timestamp 1679235063
transform 1 0 16192 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_172
timestamp 1679235063
transform 1 0 16928 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_184
timestamp 1679235063
transform 1 0 18032 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_190
timestamp 1679235063
transform 1 0 18584 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_197
timestamp 1679235063
transform 1 0 19228 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_201
timestamp 1679235063
transform 1 0 19596 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_222
timestamp 1679235063
transform 1 0 21528 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_235
timestamp 1679235063
transform 1 0 22724 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_240
timestamp 1679235063
transform 1 0 23184 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_248
timestamp 1679235063
transform 1 0 23920 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_253
timestamp 1679235063
transform 1 0 24380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_263
timestamp 1679235063
transform 1 0 25300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1679235063
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1679235063
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1679235063
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1679235063
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_51
timestamp 1679235063
transform 1 0 5796 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1679235063
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_63
timestamp 1679235063
transform 1 0 6900 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_67
timestamp 1679235063
transform 1 0 7268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_79
timestamp 1679235063
transform 1 0 8372 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_84
timestamp 1679235063
transform 1 0 8832 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_90
timestamp 1679235063
transform 1 0 9384 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_94
timestamp 1679235063
transform 1 0 9752 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1679235063
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_115
timestamp 1679235063
transform 1 0 11684 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_126
timestamp 1679235063
transform 1 0 12696 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_130
timestamp 1679235063
transform 1 0 13064 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_151
timestamp 1679235063
transform 1 0 14996 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_163
timestamp 1679235063
transform 1 0 16100 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1679235063
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_169
timestamp 1679235063
transform 1 0 16652 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_191
timestamp 1679235063
transform 1 0 18676 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_203
timestamp 1679235063
transform 1 0 19780 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_211
timestamp 1679235063
transform 1 0 20516 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_221
timestamp 1679235063
transform 1 0 21436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_77_225
timestamp 1679235063
transform 1 0 21804 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_237
timestamp 1679235063
transform 1 0 22908 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_249
timestamp 1679235063
transform 1 0 24012 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_253
timestamp 1679235063
transform 1 0 24380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1679235063
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1679235063
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1679235063
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1679235063
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1679235063
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_41
timestamp 1679235063
transform 1 0 4876 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_49
timestamp 1679235063
transform 1 0 5612 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_55
timestamp 1679235063
transform 1 0 6164 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_63
timestamp 1679235063
transform 1 0 6900 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_71
timestamp 1679235063
transform 1 0 7636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_78
timestamp 1679235063
transform 1 0 8280 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1679235063
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_91
timestamp 1679235063
transform 1 0 9476 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_95
timestamp 1679235063
transform 1 0 9844 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_98
timestamp 1679235063
transform 1 0 10120 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_104
timestamp 1679235063
transform 1 0 10672 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_112
timestamp 1679235063
transform 1 0 11408 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_116
timestamp 1679235063
transform 1 0 11776 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_122
timestamp 1679235063
transform 1 0 12328 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_134
timestamp 1679235063
transform 1 0 13432 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1679235063
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_153
timestamp 1679235063
transform 1 0 15180 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_174
timestamp 1679235063
transform 1 0 17112 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1679235063
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_197
timestamp 1679235063
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_219
timestamp 1679235063
transform 1 0 21252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_227
timestamp 1679235063
transform 1 0 21988 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_249
timestamp 1679235063
transform 1 0 24012 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1679235063
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_263
timestamp 1679235063
transform 1 0 25300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1679235063
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1679235063
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1679235063
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1679235063
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1679235063
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1679235063
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_59
timestamp 1679235063
transform 1 0 6532 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_71
timestamp 1679235063
transform 1 0 7636 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_79
timestamp 1679235063
transform 1 0 8372 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_84
timestamp 1679235063
transform 1 0 8832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_106
timestamp 1679235063
transform 1 0 10856 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1679235063
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_119
timestamp 1679235063
transform 1 0 12052 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_123
timestamp 1679235063
transform 1 0 12420 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_131
timestamp 1679235063
transform 1 0 13156 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_142
timestamp 1679235063
transform 1 0 14168 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_154
timestamp 1679235063
transform 1 0 15272 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_166
timestamp 1679235063
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_169
timestamp 1679235063
transform 1 0 16652 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_179
timestamp 1679235063
transform 1 0 17572 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_193
timestamp 1679235063
transform 1 0 18860 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1679235063
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1679235063
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1679235063
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_247
timestamp 1679235063
transform 1 0 23828 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_252
timestamp 1679235063
transform 1 0 24288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1679235063
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1679235063
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1679235063
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1679235063
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1679235063
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1679235063
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1679235063
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_65
timestamp 1679235063
transform 1 0 7084 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_71
timestamp 1679235063
transform 1 0 7636 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_76
timestamp 1679235063
transform 1 0 8096 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1679235063
transform 1 0 8464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_85
timestamp 1679235063
transform 1 0 8924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_91
timestamp 1679235063
transform 1 0 9476 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_95
timestamp 1679235063
transform 1 0 9844 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_103
timestamp 1679235063
transform 1 0 10580 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_113
timestamp 1679235063
transform 1 0 11500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1679235063
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_143
timestamp 1679235063
transform 1 0 14260 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_165
timestamp 1679235063
transform 1 0 16284 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_177
timestamp 1679235063
transform 1 0 17388 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1679235063
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1679235063
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 1679235063
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_205
timestamp 1679235063
transform 1 0 19964 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_217
timestamp 1679235063
transform 1 0 21068 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_221
timestamp 1679235063
transform 1 0 21436 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_229
timestamp 1679235063
transform 1 0 22172 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1679235063
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1679235063
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_263
timestamp 1679235063
transform 1 0 25300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1679235063
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1679235063
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1679235063
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1679235063
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1679235063
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1679235063
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1679235063
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_69
timestamp 1679235063
transform 1 0 7452 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_73
timestamp 1679235063
transform 1 0 7820 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_79
timestamp 1679235063
transform 1 0 8372 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_83
timestamp 1679235063
transform 1 0 8740 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_87
timestamp 1679235063
transform 1 0 9108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1679235063
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_106
timestamp 1679235063
transform 1 0 10856 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_113
timestamp 1679235063
transform 1 0 11500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_119
timestamp 1679235063
transform 1 0 12052 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1679235063
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1679235063
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1679235063
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1679235063
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_215
timestamp 1679235063
transform 1 0 20884 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1679235063
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_225
timestamp 1679235063
transform 1 0 21804 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_229
timestamp 1679235063
transform 1 0 22172 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_240
timestamp 1679235063
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_252
timestamp 1679235063
transform 1 0 24288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1679235063
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1679235063
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1679235063
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1679235063
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1679235063
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1679235063
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1679235063
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_65
timestamp 1679235063
transform 1 0 7084 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_71
timestamp 1679235063
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1679235063
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1679235063
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_117
timestamp 1679235063
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_129
timestamp 1679235063
transform 1 0 12972 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1679235063
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_141
timestamp 1679235063
transform 1 0 14076 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_144
timestamp 1679235063
transform 1 0 14352 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_156
timestamp 1679235063
transform 1 0 15456 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_178
timestamp 1679235063
transform 1 0 17480 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_182
timestamp 1679235063
transform 1 0 17848 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1679235063
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_199
timestamp 1679235063
transform 1 0 19412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_210
timestamp 1679235063
transform 1 0 20424 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_214
timestamp 1679235063
transform 1 0 20792 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_217
timestamp 1679235063
transform 1 0 21068 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_228
timestamp 1679235063
transform 1 0 22080 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1679235063
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_255
timestamp 1679235063
transform 1 0 24564 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_263
timestamp 1679235063
transform 1 0 25300 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1679235063
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1679235063
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1679235063
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1679235063
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1679235063
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1679235063
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1679235063
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1679235063
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_81
timestamp 1679235063
transform 1 0 8556 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_87
timestamp 1679235063
transform 1 0 9108 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_91
timestamp 1679235063
transform 1 0 9476 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_103
timestamp 1679235063
transform 1 0 10580 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1679235063
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_113
timestamp 1679235063
transform 1 0 11500 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_118
timestamp 1679235063
transform 1 0 11960 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_130
timestamp 1679235063
transform 1 0 13064 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_142
timestamp 1679235063
transform 1 0 14168 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_154
timestamp 1679235063
transform 1 0 15272 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_166
timestamp 1679235063
transform 1 0 16376 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_169
timestamp 1679235063
transform 1 0 16652 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_180
timestamp 1679235063
transform 1 0 17664 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_204
timestamp 1679235063
transform 1 0 19872 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_216
timestamp 1679235063
transform 1 0 20976 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1679235063
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1679235063
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_249
timestamp 1679235063
transform 1 0 24012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_253
timestamp 1679235063
transform 1 0 24380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1679235063
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1679235063
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1679235063
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1679235063
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1679235063
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1679235063
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1679235063
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1679235063
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1679235063
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1679235063
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1679235063
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1679235063
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1679235063
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1679235063
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1679235063
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1679235063
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1679235063
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1679235063
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_165
timestamp 1679235063
transform 1 0 16284 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_173
timestamp 1679235063
transform 1 0 17020 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_184
timestamp 1679235063
transform 1 0 18032 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_188
timestamp 1679235063
transform 1 0 18400 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_197
timestamp 1679235063
transform 1 0 19228 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_207
timestamp 1679235063
transform 1 0 20148 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_219
timestamp 1679235063
transform 1 0 21252 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_231
timestamp 1679235063
transform 1 0 22356 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_243
timestamp 1679235063
transform 1 0 23460 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1679235063
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_253
timestamp 1679235063
transform 1 0 24380 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_261
timestamp 1679235063
transform 1 0 25116 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1679235063
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1679235063
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1679235063
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1679235063
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1679235063
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1679235063
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1679235063
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1679235063
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1679235063
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1679235063
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1679235063
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1679235063
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1679235063
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1679235063
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1679235063
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1679235063
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1679235063
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1679235063
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1679235063
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1679235063
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1679235063
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1679235063
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1679235063
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1679235063
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1679235063
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1679235063
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_249
timestamp 1679235063
transform 1 0 24012 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_253
timestamp 1679235063
transform 1 0 24380 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_264
timestamp 1679235063
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1679235063
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_21
timestamp 1679235063
transform 1 0 3036 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_86_25
timestamp 1679235063
transform 1 0 3404 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1679235063
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1679235063
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1679235063
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1679235063
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1679235063
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1679235063
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1679235063
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1679235063
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1679235063
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_121
timestamp 1679235063
transform 1 0 12236 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_86_130
timestamp 1679235063
transform 1 0 13064 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_138
timestamp 1679235063
transform 1 0 13800 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1679235063
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1679235063
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1679235063
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1679235063
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1679235063
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1679235063
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1679235063
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1679235063
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1679235063
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1679235063
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1679235063
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1679235063
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_253
timestamp 1679235063
transform 1 0 24380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_259
timestamp 1679235063
transform 1 0 24932 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1679235063
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_87_3
timestamp 1679235063
transform 1 0 1380 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_25
timestamp 1679235063
transform 1 0 3404 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1679235063
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_59
timestamp 1679235063
transform 1 0 6532 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_71
timestamp 1679235063
transform 1 0 7636 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_83
timestamp 1679235063
transform 1 0 8740 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_87
timestamp 1679235063
transform 1 0 9108 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_92
timestamp 1679235063
transform 1 0 9568 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_104
timestamp 1679235063
transform 1 0 10672 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_113
timestamp 1679235063
transform 1 0 11500 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_118
timestamp 1679235063
transform 1 0 11960 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_130
timestamp 1679235063
transform 1 0 13064 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_142
timestamp 1679235063
transform 1 0 14168 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_154
timestamp 1679235063
transform 1 0 15272 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_166
timestamp 1679235063
transform 1 0 16376 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1679235063
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1679235063
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1679235063
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1679235063
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1679235063
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1679235063
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1679235063
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1679235063
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1679235063
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1679235063
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1679235063
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_3
timestamp 1679235063
transform 1 0 1380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_9
timestamp 1679235063
transform 1 0 1932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1679235063
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_29
timestamp 1679235063
transform 1 0 3772 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_39
timestamp 1679235063
transform 1 0 4692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_51
timestamp 1679235063
transform 1 0 5796 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_59
timestamp 1679235063
transform 1 0 6532 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_70
timestamp 1679235063
transform 1 0 7544 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_82
timestamp 1679235063
transform 1 0 8648 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_88_85
timestamp 1679235063
transform 1 0 8924 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_91
timestamp 1679235063
transform 1 0 9476 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_103
timestamp 1679235063
transform 1 0 10580 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_115
timestamp 1679235063
transform 1 0 11684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_127
timestamp 1679235063
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1679235063
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1679235063
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1679235063
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1679235063
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1679235063
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1679235063
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1679235063
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1679235063
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1679235063
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1679235063
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1679235063
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1679235063
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1679235063
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_253
timestamp 1679235063
transform 1 0 24380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_259
timestamp 1679235063
transform 1 0 24932 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_264
timestamp 1679235063
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1679235063
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_8
timestamp 1679235063
transform 1 0 1840 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_12
timestamp 1679235063
transform 1 0 2208 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_29
timestamp 1679235063
transform 1 0 3772 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_49
timestamp 1679235063
transform 1 0 5612 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1679235063
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_57
timestamp 1679235063
transform 1 0 6348 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_61
timestamp 1679235063
transform 1 0 6716 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_66
timestamp 1679235063
transform 1 0 7176 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_74
timestamp 1679235063
transform 1 0 7912 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_86
timestamp 1679235063
transform 1 0 9016 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1679235063
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1679235063
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1679235063
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1679235063
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1679235063
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1679235063
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1679235063
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1679235063
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1679235063
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1679235063
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1679235063
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1679235063
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1679235063
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1679235063
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1679235063
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1679235063
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1679235063
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_249
timestamp 1679235063
transform 1 0 24012 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_255
timestamp 1679235063
transform 1 0 24564 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_258
timestamp 1679235063
transform 1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1679235063
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_3
timestamp 1679235063
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_9
timestamp 1679235063
transform 1 0 1932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1679235063
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_29
timestamp 1679235063
transform 1 0 3772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_39
timestamp 1679235063
transform 1 0 4692 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_61
timestamp 1679235063
transform 1 0 6716 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1679235063
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1679235063
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_97
timestamp 1679235063
transform 1 0 10028 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_102
timestamp 1679235063
transform 1 0 10488 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_114
timestamp 1679235063
transform 1 0 11592 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_126
timestamp 1679235063
transform 1 0 12696 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1679235063
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1679235063
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1679235063
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1679235063
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1679235063
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1679235063
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1679235063
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1679235063
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1679235063
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1679235063
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1679235063
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1679235063
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1679235063
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_253
timestamp 1679235063
transform 1 0 24380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_259
timestamp 1679235063
transform 1 0 24932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1679235063
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1679235063
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_13
timestamp 1679235063
transform 1 0 2300 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_17
timestamp 1679235063
transform 1 0 2668 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_34
timestamp 1679235063
transform 1 0 4232 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1679235063
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_57
timestamp 1679235063
transform 1 0 6348 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_67
timestamp 1679235063
transform 1 0 7268 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_71
timestamp 1679235063
transform 1 0 7636 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_89
timestamp 1679235063
transform 1 0 9292 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_91_109
timestamp 1679235063
transform 1 0 11132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_113
timestamp 1679235063
transform 1 0 11500 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_118
timestamp 1679235063
transform 1 0 11960 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_125
timestamp 1679235063
transform 1 0 12604 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_133
timestamp 1679235063
transform 1 0 13340 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_145
timestamp 1679235063
transform 1 0 14444 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_157
timestamp 1679235063
transform 1 0 15548 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_165
timestamp 1679235063
transform 1 0 16284 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1679235063
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1679235063
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1679235063
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1679235063
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1679235063
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1679235063
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1679235063
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1679235063
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1679235063
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_261
timestamp 1679235063
transform 1 0 25116 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_3
timestamp 1679235063
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_9
timestamp 1679235063
transform 1 0 1932 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1679235063
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_29
timestamp 1679235063
transform 1 0 3772 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_39
timestamp 1679235063
transform 1 0 4692 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 1679235063
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_62
timestamp 1679235063
transform 1 0 6808 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1679235063
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_85
timestamp 1679235063
transform 1 0 8924 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_91
timestamp 1679235063
transform 1 0 9476 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_103
timestamp 1679235063
transform 1 0 10580 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_121
timestamp 1679235063
transform 1 0 12236 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_128
timestamp 1679235063
transform 1 0 12880 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_132
timestamp 1679235063
transform 1 0 13248 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1679235063
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_143
timestamp 1679235063
transform 1 0 14260 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_155
timestamp 1679235063
transform 1 0 15364 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_167
timestamp 1679235063
transform 1 0 16468 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_179
timestamp 1679235063
transform 1 0 17572 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_191
timestamp 1679235063
transform 1 0 18676 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1679235063
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1679235063
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1679235063
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1679235063
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1679235063
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1679235063
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1679235063
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1679235063
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_258
timestamp 1679235063
transform 1 0 24840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1679235063
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_93_3
timestamp 1679235063
transform 1 0 1380 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_14
timestamp 1679235063
transform 1 0 2392 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_34
timestamp 1679235063
transform 1 0 4232 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1679235063
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1679235063
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_67
timestamp 1679235063
transform 1 0 7268 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_73
timestamp 1679235063
transform 1 0 7820 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_90
timestamp 1679235063
transform 1 0 9384 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1679235063
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_113
timestamp 1679235063
transform 1 0 11500 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_133
timestamp 1679235063
transform 1 0 13340 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_141
timestamp 1679235063
transform 1 0 14076 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_148
timestamp 1679235063
transform 1 0 14720 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_152
timestamp 1679235063
transform 1 0 15088 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_160
timestamp 1679235063
transform 1 0 15824 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_164
timestamp 1679235063
transform 1 0 16192 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_169
timestamp 1679235063
transform 1 0 16652 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_177
timestamp 1679235063
transform 1 0 17388 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_189
timestamp 1679235063
transform 1 0 18492 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_196
timestamp 1679235063
transform 1 0 19136 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_204
timestamp 1679235063
transform 1 0 19872 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_208
timestamp 1679235063
transform 1 0 20240 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_212
timestamp 1679235063
transform 1 0 20608 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_220
timestamp 1679235063
transform 1 0 21344 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_227
timestamp 1679235063
transform 1 0 21988 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_93_232
timestamp 1679235063
transform 1 0 22448 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_235
timestamp 1679235063
transform 1 0 22724 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_239
timestamp 1679235063
transform 1 0 23092 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_244
timestamp 1679235063
transform 1 0 23552 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_251
timestamp 1679235063
transform 1 0 24196 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_255
timestamp 1679235063
transform 1 0 24564 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1679235063
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1679235063
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1679235063
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1679235063
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1679235063
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1679235063
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_39
timestamp 1679235063
transform 1 0 4692 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_45
timestamp 1679235063
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1679235063
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1679235063
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_85
timestamp 1679235063
transform 1 0 8924 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_95
timestamp 1679235063
transform 1 0 9844 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_117
timestamp 1679235063
transform 1 0 11868 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1679235063
transform 1 0 13708 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1679235063
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_147
timestamp 1679235063
transform 1 0 14628 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_151
timestamp 1679235063
transform 1 0 14996 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_161
timestamp 1679235063
transform 1 0 15916 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_167
timestamp 1679235063
transform 1 0 16468 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_173
timestamp 1679235063
transform 1 0 17020 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_180
timestamp 1679235063
transform 1 0 17664 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_184
timestamp 1679235063
transform 1 0 18032 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_189
timestamp 1679235063
transform 1 0 18492 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1679235063
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_197
timestamp 1679235063
transform 1 0 19228 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_203
timestamp 1679235063
transform 1 0 19780 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_211
timestamp 1679235063
transform 1 0 20516 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_215
timestamp 1679235063
transform 1 0 20884 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_221
timestamp 1679235063
transform 1 0 21436 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_228
timestamp 1679235063
transform 1 0 22080 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_235
timestamp 1679235063
transform 1 0 22724 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1679235063
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1679235063
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_255
timestamp 1679235063
transform 1 0 24564 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1679235063
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1679235063
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1679235063
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1679235063
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1679235063
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1679235063
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1679235063
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1679235063
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1679235063
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1679235063
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1679235063
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1679235063
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1679235063
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_113
timestamp 1679235063
transform 1 0 11500 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_118
timestamp 1679235063
transform 1 0 11960 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1679235063
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_143
timestamp 1679235063
transform 1 0 14260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_147
timestamp 1679235063
transform 1 0 14628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_153
timestamp 1679235063
transform 1 0 15180 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_161
timestamp 1679235063
transform 1 0 15916 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_165
timestamp 1679235063
transform 1 0 16284 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1679235063
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_175
timestamp 1679235063
transform 1 0 17204 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_183
timestamp 1679235063
transform 1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_191
timestamp 1679235063
transform 1 0 18676 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1679235063
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1679235063
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_203
timestamp 1679235063
transform 1 0 19780 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_211
timestamp 1679235063
transform 1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_219
timestamp 1679235063
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1679235063
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1679235063
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_231
timestamp 1679235063
transform 1 0 22356 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_239
timestamp 1679235063
transform 1 0 23092 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_243
timestamp 1679235063
transform 1 0 23460 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1679235063
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_257
timestamp 1679235063
transform 1 0 24748 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1679235063
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1679235063
transform 1 0 3036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 9108 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform -1 0 4692 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 20608 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 20332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 18032 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 12236 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 24656 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 19412 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 14260 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 16468 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform -1 0 17572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 11592 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 17388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform -1 0 20148 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform -1 0 16192 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 14444 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform -1 0 14996 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform -1 0 14904 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 20700 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 18768 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 17664 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 7544 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform -1 0 18952 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform -1 0 17388 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 17756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 6808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 7728 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform -1 0 11132 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform -1 0 13616 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform -1 0 8648 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform -1 0 18492 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform -1 0 13800 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 23460 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform -1 0 16468 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform -1 0 13892 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform -1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 24564 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform -1 0 6072 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform -1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform -1 0 7360 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 17664 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 20240 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 9108 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform -1 0 12420 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform -1 0 13800 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform -1 0 8648 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform -1 0 13432 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 10028 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 6440 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 23184 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold68
timestamp 1679235063
transform 1 0 24564 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform -1 0 9844 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform -1 0 18860 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 7820 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1679235063
transform 1 0 24564 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold73
timestamp 1679235063
transform 1 0 17480 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform -1 0 12052 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform -1 0 7544 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1679235063
transform -1 0 17940 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold78
timestamp 1679235063
transform -1 0 7728 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1679235063
transform -1 0 8096 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold80
timestamp 1679235063
transform -1 0 25024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold81
timestamp 1679235063
transform 1 0 19872 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 21988 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform -1 0 16008 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1679235063
transform -1 0 9844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold87
timestamp 1679235063
transform 1 0 17756 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold88
timestamp 1679235063
transform 1 0 19044 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1679235063
transform 1 0 20332 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1679235063
transform -1 0 10396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1679235063
transform 1 0 24564 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold92
timestamp 1679235063
transform -1 0 25300 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold93
timestamp 1679235063
transform -1 0 16100 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform -1 0 12604 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold95
timestamp 1679235063
transform 1 0 24564 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1679235063
transform -1 0 12420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform -1 0 8648 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform -1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1679235063
transform 1 0 18676 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold100
timestamp 1679235063
transform -1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold101
timestamp 1679235063
transform -1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold102
timestamp 1679235063
transform -1 0 21160 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold103 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 13616 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold104
timestamp 1679235063
transform 1 0 21988 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold105
timestamp 1679235063
transform 1 0 24564 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold106
timestamp 1679235063
transform -1 0 8280 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold107
timestamp 1679235063
transform 1 0 24564 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold108
timestamp 1679235063
transform 1 0 24564 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold109
timestamp 1679235063
transform -1 0 25300 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold110
timestamp 1679235063
transform -1 0 7544 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold111
timestamp 1679235063
transform 1 0 23276 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold112
timestamp 1679235063
transform 1 0 22816 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold113
timestamp 1679235063
transform -1 0 6072 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold114
timestamp 1679235063
transform -1 0 12420 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold115
timestamp 1679235063
transform -1 0 20516 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold116
timestamp 1679235063
transform 1 0 20516 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold117
timestamp 1679235063
transform -1 0 15272 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold118
timestamp 1679235063
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold119
timestamp 1679235063
transform 1 0 1748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold120
timestamp 1679235063
transform -1 0 3220 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold121
timestamp 1679235063
transform 1 0 3956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold122
timestamp 1679235063
transform -1 0 7268 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold123
timestamp 1679235063
transform -1 0 2392 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold124
timestamp 1679235063
transform 1 0 3956 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold125
timestamp 1679235063
transform 1 0 3956 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold126
timestamp 1679235063
transform 1 0 6532 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold127
timestamp 1679235063
transform 1 0 1564 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold128
timestamp 1679235063
transform -1 0 4692 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold129
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold130
timestamp 1679235063
transform -1 0 2300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold131
timestamp 1679235063
transform -1 0 2484 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform -1 0 1840 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 23828 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 25116 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 21988 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 21160 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 23828 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 21252 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 21252 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 25116 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform -1 0 21068 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 21896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 24564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 24472 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1679235063
transform 1 0 24472 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1679235063
transform 1 0 24472 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1679235063
transform -1 0 25392 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1679235063
transform -1 0 24104 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1679235063
transform -1 0 25392 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1679235063
transform -1 0 25392 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1679235063
transform -1 0 25392 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 25116 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1679235063
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 23828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 23000 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 23828 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform -1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1679235063
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1679235063
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform -1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1679235063
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1679235063
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1679235063
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1679235063
transform 1 0 7636 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1679235063
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1679235063
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1679235063
transform -1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1679235063
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1679235063
transform -1 0 9936 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1679235063
transform -1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1679235063
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1679235063
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1679235063
transform -1 0 11224 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1679235063
transform 1 0 10948 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1679235063
transform 1 0 11684 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform -1 0 11224 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1679235063
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1679235063
transform 1 0 3956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1679235063
transform -1 0 3680 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1679235063
transform 1 0 3128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1679235063
transform 1 0 3956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1679235063
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1679235063
transform -1 0 5612 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1679235063
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform -1 0 11960 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1679235063
transform 1 0 16652 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1679235063
transform -1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform -1 0 17664 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1679235063
transform -1 0 18676 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1679235063
transform -1 0 18492 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1679235063
transform -1 0 19780 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1679235063
transform 1 0 18860 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1679235063
transform 1 0 19412 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1679235063
transform -1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1679235063
transform -1 0 20516 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1679235063
transform 1 0 13340 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1679235063
transform 1 0 20332 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1679235063
transform -1 0 21252 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1679235063
transform 1 0 21068 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1679235063
transform -1 0 22356 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1679235063
transform 1 0 21804 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1679235063
transform 1 0 22448 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1679235063
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1679235063
transform 1 0 23092 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1679235063
transform 1 0 23276 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1679235063
transform 1 0 23920 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1679235063
transform 1 0 13708 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1679235063
transform -1 0 14628 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1679235063
transform -1 0 14720 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1679235063
transform 1 0 14812 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1679235063
transform -1 0 15916 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1679235063
transform -1 0 15916 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1679235063
transform -1 0 16192 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1679235063
transform 1 0 16836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1679235063
transform -1 0 1840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1679235063
transform -1 0 1840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1679235063
transform -1 0 1840 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1679235063
transform -1 0 1840 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1679235063
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1679235063
transform -1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1679235063
transform -1 0 25392 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1679235063
transform -1 0 25392 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1679235063
transform -1 0 25392 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1679235063
transform -1 0 25392 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1679235063
transform -1 0 25392 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input104
timestamp 1679235063
transform -1 0 25392 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1679235063
transform -1 0 24104 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1679235063
transform -1 0 24104 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  left_tile_216
timestamp 1679235063
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output107 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform -1 0 3036 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 22632 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 23920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform -1 0 19412 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform -1 0 24104 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 22080 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform -1 0 24104 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform -1 0 25392 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform -1 0 24104 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform -1 0 24104 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform -1 0 23552 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 23920 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform -1 0 18952 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform -1 0 21528 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform -1 0 23552 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform -1 0 24104 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform -1 0 13800 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 21988 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform -1 0 21252 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform -1 0 13892 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1679235063
transform 1 0 23828 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1679235063
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1679235063
transform 1 0 21988 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1679235063
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1679235063
transform 1 0 20148 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1679235063
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1679235063
transform 1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1679235063
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1679235063
transform 1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1679235063
transform 1 0 14628 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1679235063
transform -1 0 16468 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1679235063
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1679235063
transform 1 0 16836 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1679235063
transform -1 0 3404 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1679235063
transform -1 0 3496 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1679235063
transform -1 0 3496 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1679235063
transform -1 0 6072 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1679235063
transform -1 0 6808 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1679235063
transform -1 0 8556 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1679235063
transform -1 0 6808 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1679235063
transform -1 0 8648 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1679235063
transform -1 0 6072 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1679235063
transform -1 0 9292 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1679235063
transform -1 0 8648 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1679235063
transform -1 0 3496 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1679235063
transform -1 0 9384 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1679235063
transform -1 0 11132 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1679235063
transform -1 0 8648 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1679235063
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1679235063
transform 1 0 10764 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1679235063
transform -1 0 11868 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1679235063
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1679235063
transform 1 0 11868 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1679235063
transform 1 0 12236 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1679235063
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1679235063
transform -1 0 3772 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1679235063
transform -1 0 3496 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1679235063
transform -1 0 4232 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1679235063
transform -1 0 3496 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1679235063
transform -1 0 5612 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1679235063
transform -1 0 4232 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1679235063
transform -1 0 6072 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1679235063
transform -1 0 6716 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1679235063
transform -1 0 3036 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1679235063
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1679235063
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1679235063
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1679235063
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1679235063
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1679235063
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1679235063
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1679235063
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1679235063
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1679235063
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1679235063
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1679235063
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1679235063
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1679235063
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1679235063
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1679235063
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1679235063
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1679235063
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1679235063
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1679235063
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1679235063
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1679235063
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1679235063
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1679235063
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1679235063
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1679235063
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1679235063
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1679235063
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1679235063
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1679235063
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1679235063
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1679235063
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1679235063
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1679235063
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1679235063
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1679235063
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1679235063
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1679235063
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1679235063
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1679235063
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1679235063
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1679235063
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1679235063
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1679235063
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1679235063
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1679235063
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1679235063
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1679235063
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1679235063
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1679235063
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1679235063
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1679235063
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1679235063
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1679235063
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1679235063
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1679235063
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1679235063
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1679235063
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1679235063
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1679235063
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1679235063
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1679235063
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1679235063
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1679235063
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1679235063
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1679235063
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1679235063
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1679235063
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1679235063
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1679235063
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1679235063
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1679235063
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1679235063
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1679235063
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1679235063
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1679235063
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1679235063
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1679235063
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1679235063
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1679235063
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1679235063
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1679235063
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1679235063
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1679235063
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1679235063
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1679235063
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1679235063
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1679235063
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1679235063
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1679235063
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1679235063
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1679235063
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1679235063
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1679235063
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1679235063
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1679235063
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1679235063
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1679235063
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1679235063
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1679235063
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1679235063
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1679235063
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1679235063
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1679235063
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1679235063
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1679235063
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1679235063
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1679235063
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1679235063
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1679235063
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1679235063
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 20976 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17664 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 20148 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19872 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 21896 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21252 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22908 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 24196 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 19044 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 17204 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 16376 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12788 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 13064 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15180 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 21252 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 22172 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 23460 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 24840 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 23920 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 18952 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 18768 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 17296 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 16100 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 12604 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15548 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 19872 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 17296 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 10488 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17848 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 25300 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23460 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 24748 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22264 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 25300 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 24104 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22264 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 25024 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22632 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 25392 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 25392 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22172 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 24104 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 23828 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 21528 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18676 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 21252 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 21068 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 19964 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 20884 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 19872 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 16836 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 18676 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 17480 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 15272 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 16284 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 14260 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 15088 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 14260 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11684 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 13524 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 12420 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 11500 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 11592 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9292 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 10856 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 8648 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6808 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 8372 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6808 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8188 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12788 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 16100 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 13340 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9384 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10672 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 17020 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 17388 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15916 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 18676 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18032 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 21436 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21804 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 24104 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 23552 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21068 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 21712 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18124 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 19964 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19044 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3956 0 -1 50048
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9016 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 10028 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11868 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13156 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 14168 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12696 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 11224 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 10948 0 -1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 9292 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5612 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 8648 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 7360 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4232 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 8464 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5796 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8004 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9844 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 10672 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8464 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6624 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4232 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 5428 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 8464 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6256 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7820 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11040 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14904 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 18952 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 18676 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1679235063
transform -1 0 18308 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18768 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1679235063
transform -1 0 15824 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17848 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__266
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1679235063
transform -1 0 17204 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17572 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1679235063
transform -1 0 20240 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20700 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__217
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1679235063
transform -1 0 18492 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1679235063
transform -1 0 19964 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1679235063
transform -1 0 20240 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1679235063
transform -1 0 22816 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1679235063
transform -1 0 21436 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22540 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1679235063
transform -1 0 22264 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__220
timestamp 1679235063
transform -1 0 21068 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17572 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19964 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1679235063
transform 1 0 16836 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__222
timestamp 1679235063
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1679235063
transform -1 0 16376 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17480 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1679235063
transform -1 0 16376 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15824 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18308 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1679235063
transform 1 0 15272 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__267
timestamp 1679235063
transform -1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1679235063
transform -1 0 12972 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15364 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1679235063
transform -1 0 13800 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1679235063
transform -1 0 15272 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1679235063
transform -1 0 18216 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20792 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1679235063
transform -1 0 18860 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1679235063
transform -1 0 20332 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__268
timestamp 1679235063
transform 1 0 19504 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1679235063
transform -1 0 20056 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1679235063
transform -1 0 20332 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1679235063
transform -1 0 22816 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1679235063
transform -1 0 20976 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22448 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__269
timestamp 1679235063
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22172 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1679235063
transform -1 0 21528 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21804 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1679235063
transform -1 0 17572 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20240 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18676 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17572 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__270
timestamp 1679235063
transform 1 0 20884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17480 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1679235063
transform -1 0 17204 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1679235063
transform -1 0 12788 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__218
timestamp 1679235063
transform -1 0 11868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13432 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1679235063
transform -1 0 20976 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20792 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__219
timestamp 1679235063
transform 1 0 23092 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14996 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__221
timestamp 1679235063
transform 1 0 16100 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform -1 0 21712 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform -1 0 21988 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform -1 0 22908 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform -1 0 22080 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__223
timestamp 1679235063
transform -1 0 21528 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform -1 0 23736 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23736 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform -1 0 23184 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform -1 0 22816 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1679235063
transform -1 0 21068 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__229
timestamp 1679235063
transform 1 0 23736 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform -1 0 23368 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform -1 0 24012 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 24656 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform -1 0 22632 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform -1 0 20700 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__240
timestamp 1679235063
transform -1 0 20056 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform -1 0 23000 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 23920 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform -1 0 22816 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform -1 0 22816 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1679235063
transform -1 0 20424 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform -1 0 23828 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__249
timestamp 1679235063
transform -1 0 22724 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform -1 0 24012 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 24840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform -1 0 22080 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1679235063
transform -1 0 21804 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1679235063
transform -1 0 19688 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform -1 0 22724 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22816 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__250
timestamp 1679235063
transform -1 0 22264 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1679235063
transform -1 0 23184 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 24012 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20240 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20608 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform -1 0 20424 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__224
timestamp 1679235063
transform 1 0 17296 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform -1 0 17664 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform -1 0 20884 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 22632 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19596 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__225
timestamp 1679235063
transform 1 0 18032 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1679235063
transform -1 0 18216 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1679235063
transform -1 0 20056 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23000 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform -1 0 17756 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__226
timestamp 1679235063
transform 1 0 19412 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1679235063
transform -1 0 17204 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1679235063
transform -1 0 19044 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 21528 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform -1 0 18032 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17204 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__227
timestamp 1679235063
transform 1 0 15732 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1679235063
transform -1 0 15364 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1679235063
transform -1 0 17664 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 20700 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__228
timestamp 1679235063
transform 1 0 13984 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1679235063
transform -1 0 13800 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1679235063
transform -1 0 17020 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 20976 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14628 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1679235063
transform -1 0 13156 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__230
timestamp 1679235063
transform 1 0 12788 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1679235063
transform -1 0 14904 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 18952 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1679235063
transform -1 0 13616 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__231
timestamp 1679235063
transform 1 0 11868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1679235063
transform -1 0 11224 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1679235063
transform -1 0 13432 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 18308 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__232
timestamp 1679235063
transform 1 0 11684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1679235063
transform -1 0 11684 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1679235063
transform -1 0 13432 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 17664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14812 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__233
timestamp 1679235063
transform 1 0 10488 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1679235063
transform -1 0 10120 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1679235063
transform -1 0 12420 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 17112 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12236 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__234
timestamp 1679235063
transform -1 0 7820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform -1 0 8648 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform -1 0 11408 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1679235063
transform -1 0 9936 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__235
timestamp 1679235063
transform -1 0 9016 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform -1 0 12604 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14352 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1679235063
transform -1 0 11224 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__236
timestamp 1679235063
transform 1 0 11408 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform -1 0 15088 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__237
timestamp 1679235063
transform -1 0 12512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1679235063
transform -1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform -1 0 16376 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform -1 0 9936 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__238
timestamp 1679235063
transform 1 0 7820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1679235063
transform -1 0 8188 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1679235063
transform -1 0 11224 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1679235063
transform -1 0 13432 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__239
timestamp 1679235063
transform 1 0 16376 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1679235063
transform -1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1679235063
transform -1 0 15180 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__241
timestamp 1679235063
transform 1 0 17112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1679235063
transform -1 0 17664 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform -1 0 16376 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__242
timestamp 1679235063
transform 1 0 18124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform -1 0 18584 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 23000 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform -1 0 17848 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__243
timestamp 1679235063
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform -1 0 20424 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 23460 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform -1 0 20240 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__244
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform -1 0 22816 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 24104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform -1 0 22816 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__245
timestamp 1679235063
transform -1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1679235063
transform -1 0 20240 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform -1 0 22816 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform -1 0 21436 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform -1 0 22816 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__246
timestamp 1679235063
transform -1 0 22356 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 23552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1679235063
transform -1 0 18584 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__247
timestamp 1679235063
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1679235063
transform -1 0 20056 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 21804 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1679235063
transform -1 0 18952 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__248
timestamp 1679235063
transform 1 0 23276 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1679235063
transform -1 0 21068 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform -1 0 10028 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17112 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14904 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1679235063
transform -1 0 10580 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__251
timestamp 1679235063
transform -1 0 10028 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11868 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform -1 0 11500 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 11960 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17112 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1679235063
transform -1 0 13248 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15364 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__254
timestamp 1679235063
transform 1 0 13340 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform -1 0 13800 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13340 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12788 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform -1 0 16284 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18952 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1679235063
transform 1 0 11040 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15824 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform -1 0 11776 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__258
timestamp 1679235063
transform 1 0 11684 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 11960 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform -1 0 10028 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17388 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1679235063
transform -1 0 8832 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__261
timestamp 1679235063
transform 1 0 8372 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9292 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 9108 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16100 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1679235063
transform 1 0 12604 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__252
timestamp 1679235063
transform 1 0 9108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1679235063
transform -1 0 8280 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9476 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform -1 0 8280 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 8280 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12604 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16836 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1679235063
transform 1 0 8372 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__253
timestamp 1679235063
transform -1 0 7636 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1679235063
transform -1 0 8372 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 8188 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14720 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18308 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1679235063
transform -1 0 10028 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13892 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__255
timestamp 1679235063
transform 1 0 10948 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1679235063
transform -1 0 10580 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10488 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 8648 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12696 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9476 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1679235063
transform -1 0 6072 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__256
timestamp 1679235063
transform 1 0 5796 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1679235063
transform 1 0 6532 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 6164 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform -1 0 12420 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12236 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__257
timestamp 1679235063
transform -1 0 8648 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1679235063
transform -1 0 9200 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7360 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__259
timestamp 1679235063
transform -1 0 11224 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1679235063
transform -1 0 11592 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11960 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9200 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__260
timestamp 1679235063
transform 1 0 15456 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1679235063
transform -1 0 15088 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15088 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10580 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1679235063
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1679235063
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1679235063
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1679235063
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1679235063
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1679235063
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1679235063
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1679235063
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1679235063
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1679235063
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1679235063
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1679235063
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1679235063
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1679235063
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1679235063
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1679235063
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1679235063
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1679235063
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1679235063
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1679235063
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1679235063
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1679235063
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1679235063
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1679235063
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1679235063
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1679235063
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1679235063
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1679235063
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1679235063
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1679235063
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1679235063
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1679235063
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1679235063
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1679235063
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1679235063
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1679235063
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1679235063
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1679235063
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1679235063
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1679235063
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1679235063
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1679235063
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1679235063
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1679235063
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1679235063
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1679235063
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1679235063
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1679235063
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1679235063
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1679235063
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1679235063
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1679235063
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1679235063
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1679235063
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1679235063
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1679235063
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1679235063
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1679235063
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1679235063
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1679235063
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1679235063
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1679235063
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1679235063
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1679235063
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1679235063
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1679235063
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1679235063
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1679235063
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1679235063
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1679235063
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1679235063
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1679235063
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1679235063
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1679235063
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1679235063
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1679235063
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1679235063
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1679235063
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1679235063
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1679235063
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1679235063
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1679235063
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1679235063
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1679235063
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1679235063
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1679235063
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1679235063
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1679235063
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1679235063
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1679235063
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1679235063
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1679235063
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1679235063
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1679235063
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1679235063
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1679235063
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1679235063
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1679235063
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1679235063
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1679235063
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1679235063
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1679235063
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1679235063
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1679235063
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1679235063
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1679235063
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1679235063
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1679235063
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1679235063
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1679235063
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1679235063
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1679235063
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1679235063
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1679235063
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1679235063
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1679235063
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1679235063
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1679235063
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1679235063
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1679235063
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1679235063
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1679235063
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1679235063
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1679235063
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1679235063
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1679235063
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1679235063
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1679235063
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1679235063
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1679235063
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1679235063
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1679235063
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1679235063
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1679235063
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1679235063
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1679235063
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1679235063
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1679235063
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1679235063
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1679235063
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1679235063
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1679235063
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1679235063
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1679235063
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1679235063
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1679235063
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1679235063
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1679235063
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1679235063
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1679235063
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1679235063
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1679235063
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1679235063
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1679235063
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1679235063
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1679235063
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1679235063
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1679235063
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1679235063
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1679235063
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1679235063
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1679235063
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1679235063
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1679235063
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 55360 800 55480 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1490 56200 1546 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 12898 56200 12954 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 16578 56200 16634 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 16946 56200 17002 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 17314 56200 17370 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 17682 56200 17738 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 18050 56200 18106 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 18418 56200 18474 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 18786 56200 18842 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 19154 56200 19210 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 19522 56200 19578 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 19890 56200 19946 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 13266 56200 13322 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 20626 56200 20682 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 20994 56200 21050 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 21362 56200 21418 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 22098 56200 22154 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 22466 56200 22522 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 22834 56200 22890 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 23202 56200 23258 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 23570 56200 23626 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 13634 56200 13690 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 14002 56200 14058 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 14370 56200 14426 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 14738 56200 14794 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 15474 56200 15530 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 15842 56200 15898 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1858 56200 1914 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 5538 56200 5594 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 5906 56200 5962 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 6274 56200 6330 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 6642 56200 6698 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 7010 56200 7066 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 7378 56200 7434 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 7746 56200 7802 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 8114 56200 8170 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 8482 56200 8538 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 8850 56200 8906 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 2226 56200 2282 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 9218 56200 9274 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 9586 56200 9642 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 10322 56200 10378 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 11058 56200 11114 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 11426 56200 11482 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 11794 56200 11850 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 12162 56200 12218 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 12530 56200 12586 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2594 56200 2650 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 2962 56200 3018 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 3330 56200 3386 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 3698 56200 3754 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 4434 56200 4490 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 202 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 203 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 204 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 205 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 206 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 207 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 208 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 209 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 210 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 211 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 212 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 213 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 test_enable
port 214 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal input
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 5842 24378 5842 24378 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal1 4370 24582 4370 24582 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 4370 24684 4370 24684 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 3588 20570 3588 20570 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 4186 22406 4186 22406 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal2 7130 21590 7130 21590 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 7314 7786 7314 7786 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 10442 19890 10442 19890 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 8326 19890 8326 19890 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal2 8510 14042 8510 14042 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 17204 11798 17204 11798 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13570 13804 13570 13804 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 7406 15470 7406 15470 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 6762 17850 6762 17850 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal2 15640 11628 15640 11628 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal2 9430 14280 9430 14280 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal2 7866 16898 7866 16898 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 14168 18190 14168 18190 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel via1 10994 20349 10994 20349 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal2 8280 21862 8280 21862 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 12834 14586 12834 14586 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7222 21658 7222 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 5474 24786 5474 24786 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 12834 16864 12834 16864 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12282 18734 12282 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12834 21862 12834 21862 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10396 18938 10396 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10350 16456 10350 16456 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9798 19754 9798 19754 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9568 20026 9568 20026 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 7866 21488 7866 21488 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 7452 20026 7452 20026 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15594 11866 15594 11866 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7774 16592 7774 16592 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 7084 16218 7084 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14076 14042 14076 14042 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13938 18734 13938 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14030 17952 14030 17952 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10350 15470 10350 15470 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12926 14042 12926 14042 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10718 17544 10718 17544 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9016 15674 9016 15674 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9982 17238 9982 17238 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9108 16218 9108 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15272 11322 15272 11322 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7314 18258 7314 18258 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 6026 19652 6026 19652 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13708 12954 13708 12954 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14306 19822 14306 19822 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12098 18054 12098 18054 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10350 19482 10350 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11822 15096 11822 15096 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9614 16082 9614 16082 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 7774 18598 7774 18598 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8418 17306 8418 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 8878 17306 8878 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 11914 16864 11914 16864 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6578 22746 6578 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4186 22610 4186 22610 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 12098 18530 12098 18530 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10902 19924 10902 19924 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10948 20570 10948 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9890 17034 9890 17034 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11454 20162 11454 20162 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10396 20570 10396 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8326 22610 8326 22610 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8280 22746 8280 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8280 21658 8280 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 4462 26112 4462 26112 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 3450 27506 3450 27506 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 3795 29274 3795 29274 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 4002 25670 4002 25670 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 1978 21556 1978 21556 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel via1 3519 27098 3519 27098 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 6210 21862 6210 21862 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 2530 19414 2530 19414 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 3381 26010 3381 26010 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 4094 19346 4094 19346 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel via1 4255 23834 4255 23834 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 2338 55420 2338 55420 0 ccff_head
rlabel metal2 1426 2465 1426 2465 0 ccff_head_0
rlabel metal1 23828 3706 23828 3706 0 ccff_tail
rlabel metal1 1656 49266 1656 49266 0 ccff_tail_0
rlabel metal1 21712 25874 21712 25874 0 chanx_right_in[0]
rlabel metal1 24702 34170 24702 34170 0 chanx_right_in[10]
rlabel metal2 24242 37638 24242 37638 0 chanx_right_in[11]
rlabel metal1 22310 37842 22310 37842 0 chanx_right_in[12]
rlabel via2 22218 36635 22218 36635 0 chanx_right_in[13]
rlabel metal1 24288 40494 24288 40494 0 chanx_right_in[14]
rlabel metal2 22218 38607 22218 38607 0 chanx_right_in[15]
rlabel metal1 21666 42194 21666 42194 0 chanx_right_in[16]
rlabel metal3 25906 39916 25906 39916 0 chanx_right_in[17]
rlabel metal1 24196 40902 24196 40902 0 chanx_right_in[18]
rlabel metal1 22172 40494 22172 40494 0 chanx_right_in[19]
rlabel metal1 24886 29478 24886 29478 0 chanx_right_in[1]
rlabel metal3 25446 42364 25446 42364 0 chanx_right_in[20]
rlabel metal1 24610 44302 24610 44302 0 chanx_right_in[21]
rlabel metal2 24518 44693 24518 44693 0 chanx_right_in[22]
rlabel metal2 25346 45645 25346 45645 0 chanx_right_in[23]
rlabel metal2 24518 46291 24518 46291 0 chanx_right_in[24]
rlabel metal2 25254 47209 25254 47209 0 chanx_right_in[25]
rlabel metal2 25346 47413 25346 47413 0 chanx_right_in[26]
rlabel metal1 25392 49742 25392 49742 0 chanx_right_in[27]
rlabel metal2 25346 49045 25346 49045 0 chanx_right_in[28]
rlabel metal2 25346 49997 25346 49997 0 chanx_right_in[29]
rlabel metal2 21390 27268 21390 27268 0 chanx_right_in[2]
rlabel metal2 24334 28747 24334 28747 0 chanx_right_in[3]
rlabel metal1 24058 29580 24058 29580 0 chanx_right_in[4]
rlabel metal1 23230 30260 23230 30260 0 chanx_right_in[5]
rlabel metal1 25116 32878 25116 32878 0 chanx_right_in[6]
rlabel metal1 25392 33966 25392 33966 0 chanx_right_in[7]
rlabel metal1 24748 32810 24748 32810 0 chanx_right_in[8]
rlabel metal2 25346 33983 25346 33983 0 chanx_right_in[9]
rlabel metal3 25676 9724 25676 9724 0 chanx_right_out[10]
rlabel metal2 24794 9945 24794 9945 0 chanx_right_out[11]
rlabel metal2 24794 10965 24794 10965 0 chanx_right_out[12]
rlabel metal2 25162 11985 25162 11985 0 chanx_right_out[13]
rlabel metal3 25952 12988 25952 12988 0 chanx_right_out[14]
rlabel metal2 24794 13277 24794 13277 0 chanx_right_out[15]
rlabel metal2 25162 14297 25162 14297 0 chanx_right_out[16]
rlabel metal3 25952 15436 25952 15436 0 chanx_right_out[17]
rlabel metal2 24702 15589 24702 15589 0 chanx_right_out[18]
rlabel metal3 25584 17068 25584 17068 0 chanx_right_out[19]
rlabel metal1 18906 5100 18906 5100 0 chanx_right_out[1]
rlabel metal2 25162 17561 25162 17561 0 chanx_right_out[20]
rlabel metal2 25162 18513 25162 18513 0 chanx_right_out[21]
rlabel metal1 24150 19890 24150 19890 0 chanx_right_out[22]
rlabel metal1 24104 20434 24104 20434 0 chanx_right_out[23]
rlabel metal1 24150 20978 24150 20978 0 chanx_right_out[24]
rlabel metal2 24794 21165 24794 21165 0 chanx_right_out[25]
rlabel metal2 22862 23443 22862 23443 0 chanx_right_out[26]
rlabel metal1 23276 23086 23276 23086 0 chanx_right_out[27]
rlabel metal1 22954 24684 22954 24684 0 chanx_right_out[28]
rlabel metal2 24702 24973 24702 24973 0 chanx_right_out[29]
rlabel metal1 18446 4692 18446 4692 0 chanx_right_out[2]
rlabel metal1 21022 6188 21022 6188 0 chanx_right_out[3]
rlabel metal3 24894 4828 24894 4828 0 chanx_right_out[4]
rlabel metal2 24794 5389 24794 5389 0 chanx_right_out[5]
rlabel metal1 24150 6834 24150 6834 0 chanx_right_out[6]
rlabel metal3 25584 7276 25584 7276 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal2 25162 8721 25162 8721 0 chanx_right_out[9]
rlabel metal1 1610 4998 1610 4998 0 chany_bottom_in[0]
rlabel metal1 5198 3026 5198 3026 0 chany_bottom_in[10]
rlabel metal1 5934 2346 5934 2346 0 chany_bottom_in[11]
rlabel metal1 6026 3502 6026 3502 0 chany_bottom_in[12]
rlabel metal2 6486 1792 6486 1792 0 chany_bottom_in[13]
rlabel metal2 6854 1894 6854 1894 0 chany_bottom_in[14]
rlabel metal2 7222 1588 7222 1588 0 chany_bottom_in[15]
rlabel metal1 7636 2414 7636 2414 0 chany_bottom_in[16]
rlabel metal1 7820 3366 7820 3366 0 chany_bottom_in[17]
rlabel metal1 7958 3026 7958 3026 0 chany_bottom_in[18]
rlabel metal1 8648 3026 8648 3026 0 chany_bottom_in[19]
rlabel metal1 2162 4454 2162 4454 0 chany_bottom_in[1]
rlabel metal1 9476 3026 9476 3026 0 chany_bottom_in[20]
rlabel metal2 9430 2132 9430 2132 0 chany_bottom_in[21]
rlabel metal1 9844 3502 9844 3502 0 chany_bottom_in[22]
rlabel metal1 9890 2414 9890 2414 0 chany_bottom_in[23]
rlabel metal1 10856 3026 10856 3026 0 chany_bottom_in[24]
rlabel metal1 10948 3502 10948 3502 0 chany_bottom_in[25]
rlabel metal1 11500 3026 11500 3026 0 chany_bottom_in[26]
rlabel metal1 11684 4046 11684 4046 0 chany_bottom_in[27]
rlabel metal1 11730 2448 11730 2448 0 chany_bottom_in[28]
rlabel metal2 11178 2142 11178 2142 0 chany_bottom_in[29]
rlabel metal1 2622 4590 2622 4590 0 chany_bottom_in[2]
rlabel metal1 4002 3468 4002 3468 0 chany_bottom_in[3]
rlabel metal1 3542 4046 3542 4046 0 chany_bottom_in[4]
rlabel metal1 3358 3502 3358 3502 0 chany_bottom_in[5]
rlabel metal1 4002 3026 4002 3026 0 chany_bottom_in[6]
rlabel metal2 4278 1588 4278 1588 0 chany_bottom_in[7]
rlabel metal1 5106 2414 5106 2414 0 chany_bottom_in[8]
rlabel metal1 4922 3366 4922 3366 0 chany_bottom_in[9]
rlabel metal2 12742 2098 12742 2098 0 chany_bottom_out[0]
rlabel metal1 16951 4046 16951 4046 0 chany_bottom_out[10]
rlabel metal2 16790 1792 16790 1792 0 chany_bottom_out[11]
rlabel metal2 17158 1826 17158 1826 0 chany_bottom_out[12]
rlabel metal2 17526 2404 17526 2404 0 chany_bottom_out[13]
rlabel metal2 17894 2166 17894 2166 0 chany_bottom_out[14]
rlabel metal2 18262 959 18262 959 0 chany_bottom_out[15]
rlabel metal2 18630 1928 18630 1928 0 chany_bottom_out[16]
rlabel metal2 18998 2098 18998 2098 0 chany_bottom_out[17]
rlabel metal2 19366 1962 19366 1962 0 chany_bottom_out[18]
rlabel metal2 19734 2948 19734 2948 0 chany_bottom_out[19]
rlabel metal2 13110 823 13110 823 0 chany_bottom_out[1]
rlabel metal2 20102 2608 20102 2608 0 chany_bottom_out[20]
rlabel metal2 20470 2404 20470 2404 0 chany_bottom_out[21]
rlabel metal2 20838 1792 20838 1792 0 chany_bottom_out[22]
rlabel metal2 21206 1860 21206 1860 0 chany_bottom_out[23]
rlabel metal2 21574 2370 21574 2370 0 chany_bottom_out[24]
rlabel metal2 21942 3254 21942 3254 0 chany_bottom_out[25]
rlabel metal2 22310 3492 22310 3492 0 chany_bottom_out[26]
rlabel metal2 22678 1826 22678 1826 0 chany_bottom_out[27]
rlabel metal2 23046 823 23046 823 0 chany_bottom_out[28]
rlabel metal2 23414 2064 23414 2064 0 chany_bottom_out[29]
rlabel metal2 13478 2404 13478 2404 0 chany_bottom_out[2]
rlabel metal2 13846 1554 13846 1554 0 chany_bottom_out[3]
rlabel metal2 14214 1860 14214 1860 0 chany_bottom_out[4]
rlabel metal2 14582 1622 14582 1622 0 chany_bottom_out[5]
rlabel metal2 14950 2098 14950 2098 0 chany_bottom_out[6]
rlabel metal2 15318 1622 15318 1622 0 chany_bottom_out[7]
rlabel metal2 15686 1860 15686 1860 0 chany_bottom_out[8]
rlabel metal2 16054 2166 16054 2166 0 chany_bottom_out[9]
rlabel metal1 11730 54196 11730 54196 0 chany_top_in_0[0]
rlabel metal1 16652 53550 16652 53550 0 chany_top_in_0[10]
rlabel metal1 17434 54162 17434 54162 0 chany_top_in_0[11]
rlabel metal1 17388 53550 17388 53550 0 chany_top_in_0[12]
rlabel metal2 17710 55711 17710 55711 0 chany_top_in_0[13]
rlabel metal2 18262 56236 18262 56236 0 chany_top_in_0[14]
rlabel metal2 18446 55711 18446 55711 0 chany_top_in_0[15]
rlabel metal1 18952 53074 18952 53074 0 chany_top_in_0[16]
rlabel metal1 19320 53550 19320 53550 0 chany_top_in_0[17]
rlabel metal1 20470 54196 20470 54196 0 chany_top_in_0[18]
rlabel metal1 20148 53550 20148 53550 0 chany_top_in_0[19]
rlabel metal2 13294 55711 13294 55711 0 chany_top_in_0[1]
rlabel metal1 20424 53074 20424 53074 0 chany_top_in_0[20]
rlabel metal2 20654 55711 20654 55711 0 chany_top_in_0[21]
rlabel metal1 21068 53550 21068 53550 0 chany_top_in_0[22]
rlabel metal1 21850 54162 21850 54162 0 chany_top_in_0[23]
rlabel metal1 21896 53550 21896 53550 0 chany_top_in_0[24]
rlabel metal1 22218 53210 22218 53210 0 chany_top_in_0[25]
rlabel metal1 22632 54162 22632 54162 0 chany_top_in_0[26]
rlabel metal1 23092 53550 23092 53550 0 chany_top_in_0[27]
rlabel metal2 23230 55711 23230 55711 0 chany_top_in_0[28]
rlabel metal1 23874 53074 23874 53074 0 chany_top_in_0[29]
rlabel metal1 13754 53142 13754 53142 0 chany_top_in_0[2]
rlabel metal1 14306 53550 14306 53550 0 chany_top_in_0[3]
rlabel metal1 14444 53074 14444 53074 0 chany_top_in_0[4]
rlabel metal1 14674 54298 14674 54298 0 chany_top_in_0[5]
rlabel metal1 15548 54162 15548 54162 0 chany_top_in_0[6]
rlabel metal1 15640 53550 15640 53550 0 chany_top_in_0[7]
rlabel metal2 15870 55711 15870 55711 0 chany_top_in_0[8]
rlabel metal1 16721 54162 16721 54162 0 chany_top_in_0[9]
rlabel metal1 2024 49878 2024 49878 0 chany_top_out_0[0]
rlabel metal1 5566 53516 5566 53516 0 chany_top_out_0[10]
rlabel metal1 4968 53754 4968 53754 0 chany_top_out_0[11]
rlabel metal1 5934 53006 5934 53006 0 chany_top_out_0[12]
rlabel metal1 6486 52530 6486 52530 0 chany_top_out_0[13]
rlabel metal1 7176 51442 7176 51442 0 chany_top_out_0[14]
rlabel metal1 6302 53550 6302 53550 0 chany_top_out_0[15]
rlabel metal2 7774 54376 7774 54376 0 chany_top_out_0[16]
rlabel metal2 7958 56236 7958 56236 0 chany_top_out_0[17]
rlabel metal2 8510 54070 8510 54070 0 chany_top_out_0[18]
rlabel metal1 8510 53618 8510 53618 0 chany_top_out_0[19]
rlabel metal2 2254 53288 2254 53288 0 chany_top_out_0[1]
rlabel metal1 9062 53006 9062 53006 0 chany_top_out_0[20]
rlabel metal2 9660 53550 9660 53550 0 chany_top_out_0[21]
rlabel metal2 9982 55711 9982 55711 0 chany_top_out_0[22]
rlabel metal2 10350 54614 10350 54614 0 chany_top_out_0[23]
rlabel metal1 10994 52530 10994 52530 0 chany_top_out_0[24]
rlabel metal2 11086 54920 11086 54920 0 chany_top_out_0[25]
rlabel metal1 11224 54230 11224 54230 0 chany_top_out_0[26]
rlabel metal1 12098 53006 12098 53006 0 chany_top_out_0[27]
rlabel metal1 12466 53618 12466 53618 0 chany_top_out_0[28]
rlabel metal2 12558 55711 12558 55711 0 chany_top_out_0[29]
rlabel metal2 2714 52972 2714 52972 0 chany_top_out_0[2]
rlabel metal2 2990 55711 2990 55711 0 chany_top_out_0[3]
rlabel metal1 3312 52054 3312 52054 0 chany_top_out_0[4]
rlabel metal1 3358 52666 3358 52666 0 chany_top_out_0[5]
rlabel metal2 4140 52972 4140 52972 0 chany_top_out_0[6]
rlabel metal1 4094 53006 4094 53006 0 chany_top_out_0[7]
rlabel metal2 4830 54138 4830 54138 0 chany_top_out_0[8]
rlabel metal2 5382 56236 5382 56236 0 chany_top_out_0[9]
rlabel metal1 19688 41514 19688 41514 0 clknet_0_prog_clk
rlabel metal1 8878 12274 8878 12274 0 clknet_4_0_0_prog_clk
rlabel metal2 10074 48518 10074 48518 0 clknet_4_10_0_prog_clk
rlabel metal1 14260 41582 14260 41582 0 clknet_4_11_0_prog_clk
rlabel metal1 19642 33422 19642 33422 0 clknet_4_12_0_prog_clk
rlabel metal1 25300 36686 25300 36686 0 clknet_4_13_0_prog_clk
rlabel metal1 19918 43316 19918 43316 0 clknet_4_14_0_prog_clk
rlabel metal2 22034 42194 22034 42194 0 clknet_4_15_0_prog_clk
rlabel metal2 12190 11424 12190 11424 0 clknet_4_1_0_prog_clk
rlabel metal1 8372 20434 8372 20434 0 clknet_4_2_0_prog_clk
rlabel metal1 13570 20978 13570 20978 0 clknet_4_3_0_prog_clk
rlabel metal1 17204 19890 17204 19890 0 clknet_4_4_0_prog_clk
rlabel metal1 23506 16660 23506 16660 0 clknet_4_5_0_prog_clk
rlabel metal1 16330 25908 16330 25908 0 clknet_4_6_0_prog_clk
rlabel metal2 22678 21250 22678 21250 0 clknet_4_7_0_prog_clk
rlabel metal2 8050 32096 8050 32096 0 clknet_4_8_0_prog_clk
rlabel metal2 13478 35360 13478 35360 0 clknet_4_9_0_prog_clk
rlabel metal3 820 13804 820 13804 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 16252 1004 16252 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18700 1004 18700 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 21148 1004 21148 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 1426 33490 1426 33490 0 gfpga_pad_io_soc_in[0]
rlabel metal1 1840 36142 1840 36142 0 gfpga_pad_io_soc_in[1]
rlabel metal1 1472 38318 1472 38318 0 gfpga_pad_io_soc_in[2]
rlabel metal1 1472 41106 1472 41106 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1786 23596 1786 23596 0 gfpga_pad_io_soc_out[0]
rlabel metal2 2806 24599 2806 24599 0 gfpga_pad_io_soc_out[1]
rlabel metal2 2898 26605 2898 26605 0 gfpga_pad_io_soc_out[2]
rlabel metal2 2806 29223 2806 29223 0 gfpga_pad_io_soc_out[3]
rlabel metal1 1518 43282 1518 43282 0 isol_n
rlabel metal1 3726 52462 3726 52462 0 net1
rlabel metal1 20700 42058 20700 42058 0 net10
rlabel metal1 17572 43282 17572 43282 0 net100
rlabel metal1 23368 39814 23368 39814 0 net101
rlabel metal1 17250 41446 17250 41446 0 net102
rlabel metal1 21436 42670 21436 42670 0 net103
rlabel metal1 22448 38998 22448 38998 0 net104
rlabel metal1 23368 33830 23368 33830 0 net105
rlabel via2 22218 37995 22218 37995 0 net106
rlabel metal1 22126 8432 22126 8432 0 net107
rlabel metal1 9982 37706 9982 37706 0 net108
rlabel metal2 22862 9860 22862 9860 0 net109
rlabel metal1 18124 42194 18124 42194 0 net11
rlabel metal2 23966 10030 23966 10030 0 net110
rlabel metal2 23966 12478 23966 12478 0 net111
rlabel metal1 23920 11730 23920 11730 0 net112
rlabel metal1 22448 13294 22448 13294 0 net113
rlabel metal1 23690 12818 23690 12818 0 net114
rlabel metal1 23736 13906 23736 13906 0 net115
rlabel metal2 22678 18123 22678 18123 0 net116
rlabel metal1 22310 19754 22310 19754 0 net117
rlabel metal1 24104 21930 24104 21930 0 net118
rlabel metal1 19274 5236 19274 5236 0 net119
rlabel metal2 21114 38250 21114 38250 0 net12
rlabel metal1 23828 17170 23828 17170 0 net120
rlabel metal2 23966 21692 23966 21692 0 net121
rlabel metal1 23828 19822 23828 19822 0 net122
rlabel metal2 22356 23868 22356 23868 0 net123
rlabel metal1 24288 20910 24288 20910 0 net124
rlabel metal1 25024 28458 25024 28458 0 net125
rlabel metal2 24058 24650 24058 24650 0 net126
rlabel metal1 24104 23086 24104 23086 0 net127
rlabel metal1 23644 24786 23644 24786 0 net128
rlabel metal2 21206 26384 21206 26384 0 net129
rlabel metal2 17342 40358 17342 40358 0 net13
rlabel metal1 18906 4624 18906 4624 0 net130
rlabel metal1 23046 6630 23046 6630 0 net131
rlabel metal1 23368 7378 23368 7378 0 net132
rlabel metal1 24426 7718 24426 7718 0 net133
rlabel metal1 24380 8806 24380 8806 0 net134
rlabel metal2 23966 7548 23966 7548 0 net135
rlabel metal1 23966 7310 23966 7310 0 net136
rlabel metal1 23736 8466 23736 8466 0 net137
rlabel metal1 13984 3502 13984 3502 0 net138
rlabel metal1 16146 4046 16146 4046 0 net139
rlabel metal2 17250 28322 17250 28322 0 net14
rlabel metal2 19458 5882 19458 5882 0 net140
rlabel metal1 18216 3026 18216 3026 0 net141
rlabel via3 18837 4012 18837 4012 0 net142
rlabel metal1 18906 3502 18906 3502 0 net143
rlabel metal1 18676 2482 18676 2482 0 net144
rlabel metal1 19136 11050 19136 11050 0 net145
rlabel metal1 21068 3502 21068 3502 0 net146
rlabel metal1 21528 3094 21528 3094 0 net147
rlabel metal1 20884 8330 20884 8330 0 net148
rlabel metal1 13754 3060 13754 3060 0 net149
rlabel metal1 24794 41140 24794 41140 0 net15
rlabel metal1 21068 11050 21068 11050 0 net150
rlabel metal2 22218 4063 22218 4063 0 net151
rlabel metal1 23230 3026 23230 3026 0 net152
rlabel metal1 21942 5202 21942 5202 0 net153
rlabel metal1 21206 4114 21206 4114 0 net154
rlabel metal1 21804 5678 21804 5678 0 net155
rlabel metal1 22080 6290 22080 6290 0 net156
rlabel metal1 20424 7174 20424 7174 0 net157
rlabel metal1 20608 6426 20608 6426 0 net158
rlabel metal1 20332 6630 20332 6630 0 net159
rlabel metal1 14628 38386 14628 38386 0 net16
rlabel metal2 13524 9724 13524 9724 0 net160
rlabel metal1 12236 2414 12236 2414 0 net161
rlabel metal2 14306 7038 14306 7038 0 net162
rlabel metal1 13754 2414 13754 2414 0 net163
rlabel metal1 16514 3502 16514 3502 0 net164
rlabel metal2 17066 6188 17066 6188 0 net165
rlabel metal1 16698 3026 16698 3026 0 net166
rlabel metal1 16330 12682 16330 12682 0 net167
rlabel metal2 3450 46036 3450 46036 0 net168
rlabel metal1 3956 53550 3956 53550 0 net169
rlabel metal2 23138 35972 23138 35972 0 net17
rlabel metal1 4554 54162 4554 54162 0 net170
rlabel metal1 6118 53074 6118 53074 0 net171
rlabel metal1 6808 52462 6808 52462 0 net172
rlabel metal1 8832 46070 8832 46070 0 net173
rlabel metal1 6808 50966 6808 50966 0 net174
rlabel metal1 8740 52462 8740 52462 0 net175
rlabel metal1 7590 44506 7590 44506 0 net176
rlabel metal1 8924 51986 8924 51986 0 net177
rlabel metal1 8924 50490 8924 50490 0 net178
rlabel metal1 4048 42262 4048 42262 0 net179
rlabel metal1 22402 37128 22402 37128 0 net18
rlabel metal1 8786 53074 8786 53074 0 net180
rlabel metal1 10994 44982 10994 44982 0 net181
rlabel metal1 8602 54196 8602 54196 0 net182
rlabel metal1 9660 53074 9660 53074 0 net183
rlabel metal1 10212 52462 10212 52462 0 net184
rlabel metal1 11960 53550 11960 53550 0 net185
rlabel metal1 10120 51578 10120 51578 0 net186
rlabel metal2 11914 52598 11914 52598 0 net187
rlabel metal2 12650 53108 12650 53108 0 net188
rlabel metal2 12558 53142 12558 53142 0 net189
rlabel metal1 24058 37264 24058 37264 0 net19
rlabel metal1 4140 41718 4140 41718 0 net190
rlabel metal1 3450 51340 3450 51340 0 net191
rlabel metal1 4094 51952 4094 51952 0 net192
rlabel metal1 3358 52530 3358 52530 0 net193
rlabel metal1 5612 42738 5612 42738 0 net194
rlabel metal1 4186 53074 4186 53074 0 net195
rlabel metal1 6256 51986 6256 51986 0 net196
rlabel metal2 6670 48212 6670 48212 0 net197
rlabel metal2 2806 15436 2806 15436 0 net198
rlabel metal1 1932 19210 1932 19210 0 net199
rlabel metal2 4002 4998 4002 4998 0 net2
rlabel metal1 23989 38794 23989 38794 0 net20
rlabel metal2 1702 20026 1702 20026 0 net200
rlabel metal2 1794 22474 1794 22474 0 net201
rlabel metal1 5849 7854 5849 7854 0 net202
rlabel metal1 22533 17578 22533 17578 0 net203
rlabel metal2 15134 20111 15134 20111 0 net204
rlabel metal2 12374 24344 12374 24344 0 net205
rlabel metal1 23775 21590 23775 21590 0 net206
rlabel metal1 17013 24786 17013 24786 0 net207
rlabel metal1 24334 19346 24334 19346 0 net208
rlabel metal1 13669 38998 13669 38998 0 net209
rlabel via2 22494 41123 22494 41123 0 net21
rlabel metal2 9798 35122 9798 35122 0 net210
rlabel metal2 23598 35977 23598 35977 0 net211
rlabel metal1 15042 42262 15042 42262 0 net212
rlabel metal1 24709 40086 24709 40086 0 net213
rlabel metal1 17211 44778 17211 44778 0 net214
rlabel metal1 23828 37434 23828 37434 0 net215
rlabel metal1 24564 2414 24564 2414 0 net216
rlabel metal1 18768 20842 18768 20842 0 net217
rlabel metal1 12098 28594 12098 28594 0 net218
rlabel metal1 22770 33626 22770 33626 0 net219
rlabel metal1 19412 42602 19412 42602 0 net22
rlabel metal1 21436 23018 21436 23018 0 net220
rlabel metal1 15778 37978 15778 37978 0 net221
rlabel metal1 17020 23766 17020 23766 0 net222
rlabel metal1 21574 29274 21574 29274 0 net223
rlabel metal2 17250 36992 17250 36992 0 net224
rlabel metal2 17802 39202 17802 39202 0 net225
rlabel metal1 18124 39338 18124 39338 0 net226
rlabel metal1 15364 40086 15364 40086 0 net227
rlabel metal1 13708 37230 13708 37230 0 net228
rlabel metal1 23368 40494 23368 40494 0 net229
rlabel metal1 18630 42330 18630 42330 0 net23
rlabel metal2 12834 32130 12834 32130 0 net230
rlabel metal1 11362 30294 11362 30294 0 net231
rlabel metal2 11270 26622 11270 26622 0 net232
rlabel metal1 10120 26962 10120 26962 0 net233
rlabel metal1 8004 25262 8004 25262 0 net234
rlabel metal1 9246 24922 9246 24922 0 net235
rlabel metal1 11408 23154 11408 23154 0 net236
rlabel metal1 12788 21590 12788 21590 0 net237
rlabel metal2 7774 8704 7774 8704 0 net238
rlabel metal1 15870 10710 15870 10710 0 net239
rlabel metal2 21620 47804 21620 47804 0 net24
rlabel metal1 20148 32946 20148 32946 0 net240
rlabel metal1 17204 12954 17204 12954 0 net241
rlabel metal1 18308 15130 18308 15130 0 net242
rlabel metal2 20010 16320 20010 16320 0 net243
rlabel metal1 22816 16082 22816 16082 0 net244
rlabel metal1 19504 15470 19504 15470 0 net245
rlabel metal1 22356 12274 22356 12274 0 net246
rlabel metal1 20378 10710 20378 10710 0 net247
rlabel metal1 21988 13974 21988 13974 0 net248
rlabel metal1 23138 35054 23138 35054 0 net249
rlabel metal1 14766 27098 14766 27098 0 net25
rlabel metal1 23046 41582 23046 41582 0 net250
rlabel metal1 10074 38318 10074 38318 0 net251
rlabel metal1 8510 31450 8510 31450 0 net252
rlabel metal1 7682 32334 7682 32334 0 net253
rlabel metal2 13386 42432 13386 42432 0 net254
rlabel metal1 10580 33490 10580 33490 0 net255
rlabel metal1 5750 34034 5750 34034 0 net256
rlabel metal2 8786 39168 8786 39168 0 net257
rlabel metal1 11546 38318 11546 38318 0 net258
rlabel metal2 11178 41310 11178 41310 0 net259
rlabel metal1 17066 31994 17066 31994 0 net26
rlabel metal1 15088 36074 15088 36074 0 net260
rlabel metal2 8418 33218 8418 33218 0 net261
rlabel metal1 10396 23018 10396 23018 0 net262
rlabel metal1 12512 19346 12512 19346 0 net263
rlabel metal1 9568 17306 9568 17306 0 net264
rlabel metal2 9982 23936 9982 23936 0 net265
rlabel metal2 16790 22474 16790 22474 0 net266
rlabel metal2 12558 25534 12558 25534 0 net267
rlabel metal1 19596 26010 19596 26010 0 net268
rlabel metal1 23046 25262 23046 25262 0 net269
rlabel metal1 19688 36754 19688 36754 0 net27
rlabel metal1 19412 29206 19412 29206 0 net270
rlabel metal1 2990 3162 2990 3162 0 net271
rlabel metal1 3864 6426 3864 6426 0 net272
rlabel metal1 4646 53618 4646 53618 0 net273
rlabel metal2 4002 50762 4002 50762 0 net274
rlabel metal1 21160 17578 21160 17578 0 net275
rlabel metal1 20424 12682 20424 12682 0 net276
rlabel metal2 18722 17000 18722 17000 0 net277
rlabel metal2 12834 46342 12834 46342 0 net278
rlabel metal1 25208 39610 25208 39610 0 net279
rlabel metal2 20194 32844 20194 32844 0 net28
rlabel metal2 19550 47838 19550 47838 0 net280
rlabel metal1 15078 42874 15078 42874 0 net281
rlabel metal2 21482 18258 21482 18258 0 net282
rlabel metal1 16468 19754 16468 19754 0 net283
rlabel metal2 16882 45696 16882 45696 0 net284
rlabel metal1 15870 26554 15870 26554 0 net285
rlabel metal1 11132 11050 11132 11050 0 net286
rlabel metal1 17388 13226 17388 13226 0 net287
rlabel metal2 19458 11492 19458 11492 0 net288
rlabel metal1 15134 41038 15134 41038 0 net289
rlabel metal1 25116 33082 25116 33082 0 net29
rlabel metal2 15134 33762 15134 33762 0 net290
rlabel metal1 17756 17850 17756 17850 0 net291
rlabel metal1 13202 16626 13202 16626 0 net292
rlabel metal1 14076 41990 14076 41990 0 net293
rlabel metal2 21390 44642 21390 44642 0 net294
rlabel metal2 19458 14484 19458 14484 0 net295
rlabel metal1 18446 41446 18446 41446 0 net296
rlabel metal1 5290 25976 5290 25976 0 net297
rlabel metal2 7866 20026 7866 20026 0 net298
rlabel metal1 18906 44982 18906 44982 0 net299
rlabel metal1 20010 25738 20010 25738 0 net3
rlabel metal1 25162 33864 25162 33864 0 net30
rlabel metal2 16698 46308 16698 46308 0 net300
rlabel metal1 17756 14314 17756 14314 0 net301
rlabel metal2 7498 17748 7498 17748 0 net302
rlabel via1 4639 22202 4639 22202 0 net303
rlabel metal1 8280 40698 8280 40698 0 net304
rlabel metal2 9706 25296 9706 25296 0 net305
rlabel metal1 12696 11322 12696 11322 0 net306
rlabel metal1 7958 42126 7958 42126 0 net307
rlabel metal2 11270 30396 11270 30396 0 net308
rlabel metal1 17480 46138 17480 46138 0 net309
rlabel metal2 23874 33320 23874 33320 0 net31
rlabel metal1 13846 12138 13846 12138 0 net310
rlabel metal1 23966 32538 23966 32538 0 net311
rlabel metal1 16284 15130 16284 15130 0 net312
rlabel metal2 21390 15164 21390 15164 0 net313
rlabel metal1 15916 25466 15916 25466 0 net314
rlabel metal1 13248 22678 13248 22678 0 net315
rlabel metal1 9016 13498 9016 13498 0 net316
rlabel metal1 24242 22202 24242 22202 0 net317
rlabel metal1 24978 35258 24978 35258 0 net318
rlabel metal1 19872 23290 19872 23290 0 net319
rlabel metal1 22494 32368 22494 32368 0 net32
rlabel metal2 5382 39202 5382 39202 0 net320
rlabel metal1 22402 17306 22402 17306 0 net321
rlabel metal1 21436 12138 21436 12138 0 net322
rlabel metal1 6302 25194 6302 25194 0 net323
rlabel metal1 17664 31858 17664 31858 0 net324
rlabel metal1 20838 47430 20838 47430 0 net325
rlabel metal1 24518 18666 24518 18666 0 net326
rlabel metal1 23322 16626 23322 16626 0 net327
rlabel metal2 8326 32606 8326 32606 0 net328
rlabel metal1 21528 20570 21528 20570 0 net329
rlabel metal1 3772 5066 3772 5066 0 net33
rlabel metal1 11132 28118 11132 28118 0 net330
rlabel metal1 13248 35258 13248 35258 0 net331
rlabel metal1 8372 34170 8372 34170 0 net332
rlabel metal1 12926 43350 12926 43350 0 net333
rlabel metal1 10580 39950 10580 39950 0 net334
rlabel metal1 6992 34170 6992 34170 0 net335
rlabel metal2 23874 27302 23874 27302 0 net336
rlabel metal1 23414 20842 23414 20842 0 net337
rlabel metal2 24978 43486 24978 43486 0 net338
rlabel metal1 8740 28458 8740 28458 0 net339
rlabel metal2 11730 20400 11730 20400 0 net34
rlabel metal1 18262 45594 18262 45594 0 net340
rlabel metal2 8326 38046 8326 38046 0 net341
rlabel metal2 23506 45662 23506 45662 0 net342
rlabel metal1 18308 35734 18308 35734 0 net343
rlabel metal2 10166 16456 10166 16456 0 net344
rlabel metal1 11960 34986 11960 34986 0 net345
rlabel metal2 7130 26860 7130 26860 0 net346
rlabel metal2 17250 34850 17250 34850 0 net347
rlabel metal1 7084 28118 7084 28118 0 net348
rlabel metal1 7176 35802 7176 35802 0 net349
rlabel metal2 5934 5031 5934 5031 0 net35
rlabel metal1 23966 27030 23966 27030 0 net350
rlabel metal1 20746 28594 20746 28594 0 net351
rlabel metal1 11040 14790 11040 14790 0 net352
rlabel metal1 22625 31994 22625 31994 0 net353
rlabel metal1 19320 34986 19320 34986 0 net354
rlabel metal1 15134 32198 15134 32198 0 net355
rlabel metal2 9154 19652 9154 19652 0 net356
rlabel metal1 18400 37910 18400 37910 0 net357
rlabel metal2 19642 43690 19642 43690 0 net358
rlabel metal1 20010 42126 20010 42126 0 net359
rlabel metal2 16146 3876 16146 3876 0 net36
rlabel metal1 9653 27642 9653 27642 0 net360
rlabel metal1 24518 39338 24518 39338 0 net361
rlabel metal1 24518 38522 24518 38522 0 net362
rlabel metal1 14904 41650 14904 41650 0 net363
rlabel metal2 12006 35870 12006 35870 0 net364
rlabel metal2 25070 36958 25070 36958 0 net365
rlabel metal1 9200 14314 9200 14314 0 net366
rlabel metal1 7820 15674 7820 15674 0 net367
rlabel metal1 14214 26894 14214 26894 0 net368
rlabel metal2 18446 29852 18446 29852 0 net369
rlabel metal2 6762 3808 6762 3808 0 net37
rlabel metal1 17250 24106 17250 24106 0 net370
rlabel metal1 5888 20026 5888 20026 0 net371
rlabel metal1 20010 33558 20010 33558 0 net372
rlabel metal1 11270 40358 11270 40358 0 net373
rlabel metal2 22402 27676 22402 27676 0 net374
rlabel metal1 25116 31654 25116 31654 0 net375
rlabel metal1 7222 24106 7222 24106 0 net376
rlabel metal1 25116 45050 25116 45050 0 net377
rlabel metal2 24518 26622 24518 26622 0 net378
rlabel metal1 23591 42874 23591 42874 0 net379
rlabel metal1 9200 2822 9200 2822 0 net38
rlabel metal2 7038 15198 7038 15198 0 net380
rlabel metal1 21574 43826 21574 43826 0 net381
rlabel metal1 22632 36074 22632 36074 0 net382
rlabel metal2 5382 17442 5382 17442 0 net383
rlabel metal2 11730 24344 11730 24344 0 net384
rlabel metal1 19780 30294 19780 30294 0 net385
rlabel metal1 20516 21454 20516 21454 0 net386
rlabel metal1 14214 45594 14214 45594 0 net387
rlabel metal1 2254 2448 2254 2448 0 net388
rlabel metal1 3312 2958 3312 2958 0 net389
rlabel metal2 7130 2108 7130 2108 0 net39
rlabel metal1 2668 5338 2668 5338 0 net390
rlabel metal1 4462 7514 4462 7514 0 net391
rlabel metal1 2530 51986 2530 51986 0 net392
rlabel metal2 1610 51884 1610 51884 0 net393
rlabel metal2 4646 51850 4646 51850 0 net394
rlabel metal2 4278 50014 4278 50014 0 net395
rlabel metal2 7222 52598 7222 52598 0 net396
rlabel metal2 9154 52700 9154 52700 0 net397
rlabel metal1 2392 53074 2392 53074 0 net398
rlabel metal2 2714 3162 2714 3162 0 net399
rlabel metal2 21390 34102 21390 34102 0 net4
rlabel metal2 13892 2788 13892 2788 0 net40
rlabel metal1 2254 2618 2254 2618 0 net400
rlabel metal2 1794 3196 1794 3196 0 net401
rlabel metal1 8602 3706 8602 3706 0 net41
rlabel metal1 7590 3162 7590 3162 0 net42
rlabel via2 8418 3179 8418 3179 0 net43
rlabel metal1 5152 4658 5152 4658 0 net44
rlabel metal1 11454 4998 11454 4998 0 net45
rlabel metal3 11661 7956 11661 7956 0 net46
rlabel metal3 12535 10948 12535 10948 0 net47
rlabel metal1 12144 2618 12144 2618 0 net48
rlabel metal1 12420 2890 12420 2890 0 net49
rlabel metal1 25346 37638 25346 37638 0 net5
rlabel metal1 12972 3570 12972 3570 0 net50
rlabel metal1 11500 3162 11500 3162 0 net51
rlabel metal1 13294 10574 13294 10574 0 net52
rlabel metal1 17756 12138 17756 12138 0 net53
rlabel metal1 13570 4658 13570 4658 0 net54
rlabel metal1 6026 4726 6026 4726 0 net55
rlabel metal1 4186 3604 4186 3604 0 net56
rlabel metal1 5474 4114 5474 4114 0 net57
rlabel metal2 3358 3417 3358 3417 0 net58
rlabel metal1 5750 3094 5750 3094 0 net59
rlabel metal1 20976 32470 20976 32470 0 net6
rlabel via2 4094 2635 4094 2635 0 net60
rlabel metal1 7958 2482 7958 2482 0 net61
rlabel via2 5290 3621 5290 3621 0 net62
rlabel metal2 12604 43996 12604 43996 0 net63
rlabel metal2 17342 43724 17342 43724 0 net64
rlabel metal2 16606 44183 16606 44183 0 net65
rlabel metal2 17618 50762 17618 50762 0 net66
rlabel metal1 17802 47770 17802 47770 0 net67
rlabel metal2 18354 50830 18354 50830 0 net68
rlabel metal2 19366 50592 19366 50592 0 net69
rlabel metal1 17572 37162 17572 37162 0 net7
rlabel metal1 18630 46920 18630 46920 0 net70
rlabel metal1 19044 11322 19044 11322 0 net71
rlabel metal1 20562 45866 20562 45866 0 net72
rlabel metal1 20746 47226 20746 47226 0 net73
rlabel metal1 14996 52462 14996 52462 0 net74
rlabel metal2 20102 49980 20102 49980 0 net75
rlabel via2 21390 43061 21390 43061 0 net76
rlabel via2 21850 44693 21850 44693 0 net77
rlabel metal2 22126 11849 22126 11849 0 net78
rlabel metal1 20700 46002 20700 46002 0 net79
rlabel metal2 22034 40290 22034 40290 0 net8
rlabel metal1 21758 46954 21758 46954 0 net80
rlabel metal1 21620 11118 21620 11118 0 net81
rlabel metal1 22724 53686 22724 53686 0 net82
rlabel metal1 22954 44506 22954 44506 0 net83
rlabel metal1 23690 52870 23690 52870 0 net84
rlabel via3 14053 52564 14053 52564 0 net85
rlabel metal1 14536 53414 14536 53414 0 net86
rlabel metal1 15456 43418 15456 43418 0 net87
rlabel metal1 14490 11186 14490 11186 0 net88
rlabel metal1 15732 53958 15732 53958 0 net89
rlabel metal1 19458 36652 19458 36652 0 net9
rlabel metal2 15916 45540 15916 45540 0 net90
rlabel metal2 16146 50320 16146 50320 0 net91
rlabel metal3 17135 53924 17135 53924 0 net92
rlabel metal1 2852 33286 2852 33286 0 net93
rlabel metal1 2990 36006 2990 36006 0 net94
rlabel metal1 2944 38182 2944 38182 0 net95
rlabel metal1 2760 40902 2760 40902 0 net96
rlabel metal1 5842 19278 5842 19278 0 net97
rlabel metal2 24610 11169 24610 11169 0 net98
rlabel metal1 22954 40392 22954 40392 0 net99
rlabel metal2 23782 2115 23782 2115 0 prog_clk
rlabel metal1 24472 2346 24472 2346 0 prog_reset
rlabel metal2 25346 50711 25346 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 25346 51357 25346 51357 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 25346 52309 25346 52309 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25346 53023 25346 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25346 53975 25346 53975 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 25024 53550 25024 53550 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25538 55420 25538 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal3 25446 56236 25446 56236 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 2384 4012 2384 4012 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1924 6460 1924 6460 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1786 8908 1786 8908 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1740 11356 1740 11356 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 20792 15130 20792 15130 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel via1 18446 22066 18446 22066 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 19090 19482 19090 19482 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal2 19458 24208 19458 24208 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal1 15732 24038 15732 24038 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 14812 26758 14812 26758 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 18814 34442 18814 34442 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 14444 27846 14444 27846 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal2 20378 26792 20378 26792 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 19872 29138 19872 29138 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal2 19458 27761 19458 27761 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal1 20930 24684 20930 24684 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal2 22448 32436 22448 32436 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal1 24472 27438 24472 27438 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 17342 29818 17342 29818 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 20654 36686 20654 36686 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 17664 32334 17664 32334 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal1 19734 20774 19734 20774 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 19826 27506 19826 27506 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 17894 20944 17894 20944 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 14260 31110 14260 31110 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 15732 32810 15732 32810 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 14260 32742 14260 32742 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal1 18538 33286 18538 33286 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 18262 35088 18262 35088 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 22586 33456 22586 33456 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 23782 21318 23782 21318 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal2 22126 30209 22126 30209 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 21666 23188 21666 23188 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal2 15686 36822 15686 36822 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal1 20056 31926 20056 31926 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 18078 24174 18078 24174 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal1 16698 37978 16698 37978 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 23322 30770 23322 30770 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal2 22034 34714 22034 34714 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal2 24058 32130 24058 32130 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 22678 41038 22678 41038 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal1 20332 41990 20332 41990 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 21988 45254 21988 45254 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 19734 42806 19734 42806 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal1 18538 43078 18538 43078 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal1 19826 45050 19826 45050 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 19136 44370 19136 44370 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 18492 44166 18492 44166 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal2 18814 47600 18814 47600 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal2 17158 43758 17158 43758 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 17204 45934 17204 45934 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal1 17250 46342 17250 46342 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 17802 43894 17802 43894 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal2 16606 41922 16606 41922 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 17480 45458 17480 45458 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal2 16698 43078 16698 43078 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 23736 38862 23736 38862 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal1 22172 39950 22172 39950 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 22632 40562 22632 40562 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal2 13478 33422 13478 33422 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal1 14306 42194 14306 42194 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal1 12604 37230 12604 37230 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal1 10948 31314 10948 31314 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 12052 36142 12052 36142 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal2 11730 34476 11730 34476 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal1 12742 25840 12742 25840 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal1 14858 28628 14858 28628 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal2 7682 28322 7682 28322 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal1 9430 27982 9430 27982 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 7498 27404 7498 27404 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal2 12834 28390 12834 28390 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 11500 25874 11500 25874 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 12995 27506 12995 27506 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal2 13846 23868 13846 23868 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal1 13110 24786 13110 24786 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal1 15916 21114 15916 21114 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal1 14536 20842 14536 20842 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal1 10902 12070 10902 12070 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 14490 20026 14490 20026 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal1 9568 8398 9568 8398 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 14582 11526 14582 11526 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal1 12604 11186 12604 11186 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal1 24288 36006 24288 36006 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 24610 40460 24610 40460 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal1 22494 37230 22494 37230 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal1 17434 12750 17434 12750 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal2 16054 13430 16054 13430 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal1 18124 15674 18124 15674 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal2 15686 16048 15686 16048 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal2 19826 17034 19826 17034 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal1 17020 17646 17020 17646 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 24104 17850 24104 17850 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal1 19688 17510 19688 17510 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal2 23782 18394 23782 18394 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal2 22310 19737 22310 19737 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal1 22494 13906 22494 13906 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal2 20838 16252 20838 16252 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal2 19918 11084 19918 11084 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal1 18952 12342 18952 12342 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal2 18814 14722 18814 14722 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 24150 36890 24150 36890 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal1 22862 37774 22862 37774 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal2 24426 38148 24426 38148 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal1 23598 40018 23598 40018 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal1 22448 43826 22448 43826 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 11822 46444 11822 46444 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal1 17296 42126 17296 42126 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal1 12466 44268 12466 44268 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 8096 38318 8096 38318 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal2 6026 36448 6026 36448 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal2 15962 36992 15962 36992 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal1 9660 34034 9660 34034 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal2 7590 34102 7590 34102 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal2 12558 35054 12558 35054 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 6624 32946 6624 32946 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 12972 44846 12972 44846 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 17802 42772 17802 42772 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 14858 44166 14858 44166 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal1 9108 34714 9108 34714 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal1 14996 32742 14996 32742 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 13386 34408 13386 34408 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal1 6026 38964 6026 38964 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 12466 34782 12466 34782 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal1 5520 34510 5520 34510 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal2 8602 42228 8602 42228 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 9752 40494 9752 40494 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal2 8602 39338 8602 39338 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 10074 42228 10074 42228 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 14904 43146 14904 43146 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal2 13478 40324 13478 40324 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 13478 43826 13478 43826 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal1 13386 39848 13386 39848 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal1 19228 41582 19228 41582 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 17618 39406 17618 39406 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal1 14858 31892 14858 31892 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal1 10028 35122 10028 35122 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 18446 6766 18446 6766 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal2 18354 26928 18354 26928 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18998 32198 18998 32198 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16238 22406 16238 22406 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18216 22134 18216 22134 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17158 21896 17158 21896 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17480 21862 17480 21862 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16974 7446 16974 7446 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal2 15870 30056 15870 30056 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17710 34646 17710 34646 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13984 26418 13984 26418 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13156 25466 13156 25466 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15088 25194 15088 25194 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14766 25262 14766 25262 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15364 25126 15364 25126 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 19964 8942 19964 8942 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal2 19826 29886 19826 29886 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 29614 20378 29614 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19504 25874 19504 25874 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20010 27132 20010 27132 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19918 25296 19918 25296 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19044 19822 19044 19822 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 21436 8534 21436 8534 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal2 22954 29750 22954 29750 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22816 29614 22816 29614 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22586 25330 22586 25330 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21022 27268 21022 27268 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22310 25024 22310 25024 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 21528 19686 21528 19686 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16698 8942 16698 8942 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 17802 32538 17802 32538 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18768 32470 18768 32470 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18354 29274 18354 29274 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17158 28594 17158 28594 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17158 28526 17158 28526 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17112 28390 17112 28390 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19596 6358 19596 6358 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal1 20056 25262 20056 25262 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20286 25194 20286 25194 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19734 20502 19734 20502 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19550 20808 19550 20808 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19642 17306 19642 17306 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13616 9622 13616 9622 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal1 16744 33626 16744 33626 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16836 33558 16836 33558 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14766 29274 14766 29274 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13294 29274 13294 29274 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12834 20910 12834 20910 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17940 10030 17940 10030 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal1 21114 36210 21114 36210 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20884 36006 20884 36006 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21390 33286 21390 33286 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19320 19890 19320 19890 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15594 11186 15594 11186 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal2 20654 27200 20654 27200 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 26350 22862 26350 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21758 24140 21758 24140 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22540 21658 22540 21658 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22310 21658 22310 21658 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 21574 14994 21574 14994 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10764 10778 10764 10778 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal2 14582 38318 14582 38318 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14766 38080 14766 38080 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11684 37638 11684 37638 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17756 7786 17756 7786 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 17802 27506 17802 27506 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 32198 19688 32198 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15870 24956 15870 24956 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16238 23834 16238 23834 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17434 23834 17434 23834 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16928 23834 16928 23834 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16238 18734 16238 18734 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 22310 28118 22310 28118 0 sb_0__1_.mux_right_track_0.out
rlabel metal2 22402 32164 22402 32164 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22494 32623 22494 32623 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23046 30702 23046 30702 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23322 30192 23322 30192 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23966 29852 23966 29852 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23368 32810 23368 32810 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 20102 42738 20102 42738 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20332 41242 20332 41242 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20378 40800 20378 40800 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18676 36890 18676 36890 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22402 33728 22402 33728 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22678 33014 22678 33014 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 19780 47158 19780 47158 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19504 40154 19504 40154 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18262 38522 18262 38522 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22862 33745 22862 33745 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22839 32470 22839 32470 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 17388 43418 17388 43418 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18078 43146 18078 43146 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17894 39610 17894 39610 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20746 32402 20746 32402 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21390 33014 21390 33014 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 17848 47974 17848 47974 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17204 41242 17204 41242 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15640 40154 15640 40154 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19044 32878 19044 32878 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21114 27166 21114 27166 0 sb_0__1_.mux_right_track_18.out
rlabel metal1 16928 47430 16928 47430 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16468 41446 16468 41446 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13800 37094 13800 37094 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17572 37298 17572 37298 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24702 34714 24702 34714 0 sb_0__1_.mux_right_track_2.out
rlabel metal2 25070 43996 25070 43996 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23874 40154 23874 40154 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 37944 21022 37944 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24058 38998 24058 38998 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23460 39066 23460 39066 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24150 38726 24150 38726 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 22862 21760 22862 21760 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 15088 43078 15088 43078 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14398 34510 14398 34510 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13800 32538 13800 32538 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15824 27302 15824 27302 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21988 19822 21988 19822 0 sb_0__1_.mux_right_track_22.out
rlabel metal1 13524 33898 13524 33898 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12880 33830 12880 33830 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11178 30158 11178 30158 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17296 25262 17296 25262 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19412 19754 19412 19754 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 13248 25942 13248 25942 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13018 26248 13018 26248 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14490 21930 14490 21930 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23322 18190 23322 18190 0 sb_0__1_.mux_right_track_26.out
rlabel metal1 13938 31144 13938 31144 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11040 27098 11040 27098 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12742 24854 12742 24854 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23230 17136 23230 17136 0 sb_0__1_.mux_right_track_28.out
rlabel metal2 10902 26860 10902 26860 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9798 25194 9798 25194 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15088 20502 15088 20502 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21068 16558 21068 16558 0 sb_0__1_.mux_right_track_30.out
rlabel metal1 12190 23698 12190 23698 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12144 23834 12144 23834 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16698 19822 16698 19822 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22425 14994 22425 14994 0 sb_0__1_.mux_right_track_32.out
rlabel metal2 14582 24820 14582 24820 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14214 23086 14214 23086 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17848 19346 17848 19346 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23138 14382 23138 14382 0 sb_0__1_.mux_right_track_34.out
rlabel metal1 16376 21658 16376 21658 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13570 21318 13570 21318 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19734 17170 19734 17170 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22034 10574 22034 10574 0 sb_0__1_.mux_right_track_36.out
rlabel metal1 14306 22066 14306 22066 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10304 11866 10304 11866 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8004 8602 8004 8602 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16146 10574 16146 10574 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21298 9554 21298 9554 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 15318 10574 15318 10574 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17595 10642 17595 10642 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24426 26350 24426 26350 0 sb_0__1_.mux_right_track_4.out
rlabel metal2 22126 41276 22126 41276 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22034 38522 22034 38522 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22540 34714 22540 34714 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22586 34612 22586 34612 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23322 34510 23322 34510 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22724 10642 22724 10642 0 sb_0__1_.mux_right_track_40.out
rlabel metal1 16790 12818 16790 12818 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19044 12614 19044 12614 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23598 8942 23598 8942 0 sb_0__1_.mux_right_track_44.out
rlabel metal1 18354 14926 18354 14926 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 11730 21988 11730 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24978 8942 24978 8942 0 sb_0__1_.mux_right_track_46.out
rlabel metal2 19918 17544 19918 17544 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22494 12206 22494 12206 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24886 9962 24886 9962 0 sb_0__1_.mux_right_track_48.out
rlabel metal2 20194 17408 20194 17408 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23874 12240 23874 12240 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23874 9962 23874 9962 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 22540 18258 22540 18258 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20562 15674 20562 15674 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23046 18054 23046 18054 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24702 6766 24702 6766 0 sb_0__1_.mux_right_track_52.out
rlabel metal2 21758 14144 21758 14144 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 11084 23322 11084 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22494 4590 22494 4590 0 sb_0__1_.mux_right_track_54.out
rlabel metal2 19550 11424 19550 11424 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 7854 21528 7854 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23506 5678 23506 5678 0 sb_0__1_.mux_right_track_56.out
rlabel metal1 20056 14042 20056 14042 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 14042 21528 14042 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24886 27914 24886 27914 0 sb_0__1_.mux_right_track_6.out
rlabel metal1 23368 38386 23368 38386 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23092 36890 23092 36890 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 34170 20746 34170 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24472 36142 24472 36142 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24472 36074 24472 36074 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 24610 33354 24610 33354 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24196 34714 24196 34714 0 sb_0__1_.mux_right_track_8.out
rlabel metal1 22356 43622 22356 43622 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22218 43146 22218 43146 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20608 38794 20608 38794 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22678 42432 22678 42432 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22816 41242 22816 41242 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 24104 37332 24104 37332 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12144 49946 12144 49946 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 11178 43962 11178 43962 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14398 43418 14398 43418 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14352 37638 14352 37638 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10626 38522 10626 38522 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 11914 45186 11914 45186 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11684 40970 11684 40970 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11454 47974 11454 47974 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8050 45050 8050 45050 0 sb_0__1_.mux_top_track_10.out
rlabel metal1 10212 37978 10212 37978 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16146 37570 16146 37570 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10902 33898 10902 33898 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8694 33830 8694 33830 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8372 37230 8372 37230 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 9154 35632 9154 35632 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7958 37434 7958 37434 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7958 43418 7958 43418 0 sb_0__1_.mux_top_track_12.out
rlabel metal1 12236 33626 12236 33626 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16790 31178 16790 31178 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8418 29920 8418 29920 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11730 33592 11730 33592 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 8418 33660 8418 33660 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7820 35258 7820 35258 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 12834 50932 12834 50932 0 sb_0__1_.mux_top_track_2.out
rlabel metal1 17158 42568 17158 42568 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18906 43894 18906 43894 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13340 42126 13340 42126 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14628 43962 14628 43962 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 13754 43894 13754 43894 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13478 45322 13478 45322 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9016 43962 9016 43962 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 14582 34714 14582 34714 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18124 34442 18124 34442 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10028 33422 10028 33422 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13800 34714 13800 34714 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10718 33626 10718 33626 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10396 37094 10396 37094 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 6118 47974 6118 47974 0 sb_0__1_.mux_top_track_28.out
rlabel metal1 10534 36142 10534 36142 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14306 35122 14306 35122 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8280 36346 8280 36346 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 6072 34714 6072 34714 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 6256 39066 6256 39066 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7452 47226 7452 47226 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 12742 39474 12742 39474 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12282 39304 12282 39304 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9292 39066 9292 39066 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9062 42534 9062 42534 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11822 47770 11822 47770 0 sb_0__1_.mux_top_track_4.out
rlabel metal2 16330 40732 16330 40732 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18998 38488 18998 38488 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11178 34170 11178 34170 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15318 40698 15318 40698 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11776 38522 11776 38522 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11730 44982 11730 44982 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9292 47770 9292 47770 0 sb_0__1_.mux_top_track_44.out
rlabel metal1 14674 43690 14674 43690 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11960 39610 11960 39610 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11500 43894 11500 43894 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9936 46682 9936 46682 0 sb_0__1_.mux_top_track_52.out
rlabel metal2 19550 39168 19550 39168 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18078 37978 18078 37978 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15272 36346 15272 36346 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14628 39542 14628 39542 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9752 51374 9752 51374 0 sb_0__1_.mux_top_track_6.out
rlabel metal1 10626 38930 10626 38930 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12558 39032 12558 39032 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 31994 13478 31994 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9246 33626 9246 33626 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10028 39066 10028 39066 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9430 35258 9430 35258 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9016 46546 9016 46546 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9430 40358 9430 40358 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 17204 42670 17204 42670 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1211 50524 1211 50524 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1832 52972 1832 52972 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
