magic
tech sky130A
magscale 1 2
timestamp 1679320555
<< obsli1 >>
rect 1104 2159 49864 54417
<< obsm1 >>
rect 934 2048 49864 54664
<< metal2 >>
rect 1582 56200 1638 57000
rect 2226 56200 2282 57000
rect 2870 56200 2926 57000
rect 3514 56200 3570 57000
rect 4158 56200 4214 57000
rect 4802 56200 4858 57000
rect 5446 56200 5502 57000
rect 6090 56200 6146 57000
rect 6734 56200 6790 57000
rect 7378 56200 7434 57000
rect 8022 56200 8078 57000
rect 8666 56200 8722 57000
rect 9310 56200 9366 57000
rect 9954 56200 10010 57000
rect 10598 56200 10654 57000
rect 11242 56200 11298 57000
rect 11886 56200 11942 57000
rect 12530 56200 12586 57000
rect 13174 56200 13230 57000
rect 13818 56200 13874 57000
rect 14462 56200 14518 57000
rect 15106 56200 15162 57000
rect 15750 56200 15806 57000
rect 16394 56200 16450 57000
rect 17038 56200 17094 57000
rect 17682 56200 17738 57000
rect 18326 56200 18382 57000
rect 18970 56200 19026 57000
rect 19614 56200 19670 57000
rect 20258 56200 20314 57000
rect 20902 56200 20958 57000
rect 21546 56200 21602 57000
rect 22190 56200 22246 57000
rect 22834 56200 22890 57000
rect 23478 56200 23534 57000
rect 24122 56200 24178 57000
rect 24766 56200 24822 57000
rect 25410 56200 25466 57000
rect 26054 56200 26110 57000
rect 26698 56200 26754 57000
rect 27342 56200 27398 57000
rect 27986 56200 28042 57000
rect 28630 56200 28686 57000
rect 29274 56200 29330 57000
rect 29918 56200 29974 57000
rect 30562 56200 30618 57000
rect 31206 56200 31262 57000
rect 31850 56200 31906 57000
rect 32494 56200 32550 57000
rect 33138 56200 33194 57000
rect 33782 56200 33838 57000
rect 34426 56200 34482 57000
rect 35070 56200 35126 57000
rect 35714 56200 35770 57000
rect 36358 56200 36414 57000
rect 37002 56200 37058 57000
rect 37646 56200 37702 57000
rect 38290 56200 38346 57000
rect 38934 56200 38990 57000
rect 39578 56200 39634 57000
rect 40222 56200 40278 57000
rect 42154 56200 42210 57000
rect 42798 56200 42854 57000
rect 43442 56200 43498 57000
rect 44086 56200 44142 57000
rect 44730 56200 44786 57000
rect 45374 56200 45430 57000
rect 46018 56200 46074 57000
rect 46662 56200 46718 57000
rect 47306 56200 47362 57000
rect 47950 56200 48006 57000
rect 48594 56200 48650 57000
rect 49238 56200 49294 57000
rect 2226 0 2282 800
rect 5538 0 5594 800
rect 8850 0 8906 800
rect 12162 0 12218 800
rect 15474 0 15530 800
rect 18786 0 18842 800
rect 22098 0 22154 800
rect 25410 0 25466 800
rect 28722 0 28778 800
rect 32034 0 32090 800
rect 35346 0 35402 800
rect 38658 0 38714 800
rect 41970 0 42026 800
rect 45282 0 45338 800
rect 48594 0 48650 800
<< obsm2 >>
rect 938 56144 1526 56250
rect 1694 56144 2170 56250
rect 2338 56144 2814 56250
rect 2982 56144 3458 56250
rect 3626 56144 4102 56250
rect 4270 56144 4746 56250
rect 4914 56144 5390 56250
rect 5558 56144 6034 56250
rect 6202 56144 6678 56250
rect 6846 56144 7322 56250
rect 7490 56144 7966 56250
rect 8134 56144 8610 56250
rect 8778 56144 9254 56250
rect 9422 56144 9898 56250
rect 10066 56144 10542 56250
rect 10710 56144 11186 56250
rect 11354 56144 11830 56250
rect 11998 56144 12474 56250
rect 12642 56144 13118 56250
rect 13286 56144 13762 56250
rect 13930 56144 14406 56250
rect 14574 56144 15050 56250
rect 15218 56144 15694 56250
rect 15862 56144 16338 56250
rect 16506 56144 16982 56250
rect 17150 56144 17626 56250
rect 17794 56144 18270 56250
rect 18438 56144 18914 56250
rect 19082 56144 19558 56250
rect 19726 56144 20202 56250
rect 20370 56144 20846 56250
rect 21014 56144 21490 56250
rect 21658 56144 22134 56250
rect 22302 56144 22778 56250
rect 22946 56144 23422 56250
rect 23590 56144 24066 56250
rect 24234 56144 24710 56250
rect 24878 56144 25354 56250
rect 25522 56144 25998 56250
rect 26166 56144 26642 56250
rect 26810 56144 27286 56250
rect 27454 56144 27930 56250
rect 28098 56144 28574 56250
rect 28742 56144 29218 56250
rect 29386 56144 29862 56250
rect 30030 56144 30506 56250
rect 30674 56144 31150 56250
rect 31318 56144 31794 56250
rect 31962 56144 32438 56250
rect 32606 56144 33082 56250
rect 33250 56144 33726 56250
rect 33894 56144 34370 56250
rect 34538 56144 35014 56250
rect 35182 56144 35658 56250
rect 35826 56144 36302 56250
rect 36470 56144 36946 56250
rect 37114 56144 37590 56250
rect 37758 56144 38234 56250
rect 38402 56144 38878 56250
rect 39046 56144 39522 56250
rect 39690 56144 40166 56250
rect 40334 56144 42098 56250
rect 42266 56144 42742 56250
rect 42910 56144 43386 56250
rect 43554 56144 44030 56250
rect 44198 56144 44674 56250
rect 44842 56144 45318 56250
rect 45486 56144 45962 56250
rect 46130 56144 46606 56250
rect 46774 56144 47250 56250
rect 47418 56144 47894 56250
rect 48062 56144 48538 56250
rect 48706 56144 49182 56250
rect 49350 56144 49386 56250
rect 938 856 49386 56144
rect 938 800 2170 856
rect 2338 800 5482 856
rect 5650 800 8794 856
rect 8962 800 12106 856
rect 12274 800 15418 856
rect 15586 800 18730 856
rect 18898 800 22042 856
rect 22210 800 25354 856
rect 25522 800 28666 856
rect 28834 800 31978 856
rect 32146 800 35290 856
rect 35458 800 38602 856
rect 38770 800 41914 856
rect 42082 800 45226 856
rect 45394 800 48538 856
rect 48706 800 49386 856
<< metal3 >>
rect 0 54544 800 54664
rect 50200 54544 51000 54664
rect 0 53728 800 53848
rect 50200 53728 51000 53848
rect 0 52912 800 53032
rect 50200 52912 51000 53032
rect 0 52096 800 52216
rect 50200 52096 51000 52216
rect 0 51280 800 51400
rect 50200 51280 51000 51400
rect 0 50464 800 50584
rect 50200 50464 51000 50584
rect 0 49648 800 49768
rect 50200 49648 51000 49768
rect 0 48832 800 48952
rect 50200 48832 51000 48952
rect 0 48016 800 48136
rect 50200 48016 51000 48136
rect 0 47200 800 47320
rect 50200 47200 51000 47320
rect 0 46384 800 46504
rect 50200 46384 51000 46504
rect 0 45568 800 45688
rect 50200 45568 51000 45688
rect 0 44752 800 44872
rect 50200 44752 51000 44872
rect 0 43936 800 44056
rect 50200 43936 51000 44056
rect 0 43120 800 43240
rect 50200 43120 51000 43240
rect 0 42304 800 42424
rect 50200 42304 51000 42424
rect 0 41488 800 41608
rect 50200 41488 51000 41608
rect 0 40672 800 40792
rect 50200 40672 51000 40792
rect 0 39856 800 39976
rect 50200 39856 51000 39976
rect 0 39040 800 39160
rect 50200 39040 51000 39160
rect 0 38224 800 38344
rect 50200 38224 51000 38344
rect 0 37408 800 37528
rect 50200 37408 51000 37528
rect 0 36592 800 36712
rect 50200 36592 51000 36712
rect 0 35776 800 35896
rect 50200 35776 51000 35896
rect 0 34960 800 35080
rect 50200 34960 51000 35080
rect 0 34144 800 34264
rect 50200 34144 51000 34264
rect 0 33328 800 33448
rect 50200 33328 51000 33448
rect 0 32512 800 32632
rect 50200 32512 51000 32632
rect 0 31696 800 31816
rect 50200 31696 51000 31816
rect 0 30880 800 31000
rect 50200 30880 51000 31000
rect 0 30064 800 30184
rect 50200 30064 51000 30184
rect 0 29248 800 29368
rect 50200 29248 51000 29368
rect 0 28432 800 28552
rect 50200 28432 51000 28552
rect 0 27616 800 27736
rect 50200 27616 51000 27736
rect 0 26800 800 26920
rect 50200 26800 51000 26920
rect 0 25984 800 26104
rect 50200 25984 51000 26104
rect 0 25168 800 25288
rect 50200 25168 51000 25288
rect 0 24352 800 24472
rect 50200 24352 51000 24472
rect 0 23536 800 23656
rect 50200 23536 51000 23656
rect 0 22720 800 22840
rect 50200 22720 51000 22840
rect 0 21904 800 22024
rect 50200 21904 51000 22024
rect 0 21088 800 21208
rect 50200 21088 51000 21208
rect 0 20272 800 20392
rect 50200 20272 51000 20392
rect 0 19456 800 19576
rect 50200 19456 51000 19576
rect 0 18640 800 18760
rect 50200 18640 51000 18760
rect 0 17824 800 17944
rect 50200 17824 51000 17944
rect 0 17008 800 17128
rect 50200 17008 51000 17128
rect 0 16192 800 16312
rect 50200 16192 51000 16312
rect 0 15376 800 15496
rect 50200 15376 51000 15496
rect 0 14560 800 14680
rect 50200 14560 51000 14680
rect 0 13744 800 13864
rect 50200 13744 51000 13864
rect 0 12928 800 13048
rect 50200 12928 51000 13048
rect 0 12112 800 12232
rect 50200 12112 51000 12232
rect 0 11296 800 11416
rect 50200 11296 51000 11416
rect 0 10480 800 10600
rect 50200 10480 51000 10600
rect 0 9664 800 9784
rect 50200 9664 51000 9784
rect 0 8848 800 8968
rect 50200 8848 51000 8968
rect 0 8032 800 8152
rect 50200 8032 51000 8152
rect 0 7216 800 7336
rect 50200 7216 51000 7336
rect 0 6400 800 6520
rect 50200 6400 51000 6520
rect 0 5584 800 5704
rect 50200 5584 51000 5704
rect 0 4768 800 4888
rect 50200 4768 51000 4888
rect 0 3952 800 4072
rect 50200 3952 51000 4072
rect 0 3136 800 3256
rect 50200 3136 51000 3256
rect 50200 2320 51000 2440
<< obsm3 >>
rect 880 54464 50120 54637
rect 800 53928 50200 54464
rect 880 53648 50120 53928
rect 800 53112 50200 53648
rect 880 52832 50120 53112
rect 800 52296 50200 52832
rect 880 52016 50120 52296
rect 800 51480 50200 52016
rect 880 51200 50120 51480
rect 800 50664 50200 51200
rect 880 50384 50120 50664
rect 800 49848 50200 50384
rect 880 49568 50120 49848
rect 800 49032 50200 49568
rect 880 48752 50120 49032
rect 800 48216 50200 48752
rect 880 47936 50120 48216
rect 800 47400 50200 47936
rect 880 47120 50120 47400
rect 800 46584 50200 47120
rect 880 46304 50120 46584
rect 800 45768 50200 46304
rect 880 45488 50120 45768
rect 800 44952 50200 45488
rect 880 44672 50120 44952
rect 800 44136 50200 44672
rect 880 43856 50120 44136
rect 800 43320 50200 43856
rect 880 43040 50120 43320
rect 800 42504 50200 43040
rect 880 42224 50120 42504
rect 800 41688 50200 42224
rect 880 41408 50120 41688
rect 800 40872 50200 41408
rect 880 40592 50120 40872
rect 800 40056 50200 40592
rect 880 39776 50120 40056
rect 800 39240 50200 39776
rect 880 38960 50120 39240
rect 800 38424 50200 38960
rect 880 38144 50120 38424
rect 800 37608 50200 38144
rect 880 37328 50120 37608
rect 800 36792 50200 37328
rect 880 36512 50120 36792
rect 800 35976 50200 36512
rect 880 35696 50120 35976
rect 800 35160 50200 35696
rect 880 34880 50120 35160
rect 800 34344 50200 34880
rect 880 34064 50120 34344
rect 800 33528 50200 34064
rect 880 33248 50120 33528
rect 800 32712 50200 33248
rect 880 32432 50120 32712
rect 800 31896 50200 32432
rect 880 31616 50120 31896
rect 800 31080 50200 31616
rect 880 30800 50120 31080
rect 800 30264 50200 30800
rect 880 29984 50120 30264
rect 800 29448 50200 29984
rect 880 29168 50120 29448
rect 800 28632 50200 29168
rect 880 28352 50120 28632
rect 800 27816 50200 28352
rect 880 27536 50120 27816
rect 800 27000 50200 27536
rect 880 26720 50120 27000
rect 800 26184 50200 26720
rect 880 25904 50120 26184
rect 800 25368 50200 25904
rect 880 25088 50120 25368
rect 800 24552 50200 25088
rect 880 24272 50120 24552
rect 800 23736 50200 24272
rect 880 23456 50120 23736
rect 800 22920 50200 23456
rect 880 22640 50120 22920
rect 800 22104 50200 22640
rect 880 21824 50120 22104
rect 800 21288 50200 21824
rect 880 21008 50120 21288
rect 800 20472 50200 21008
rect 880 20192 50120 20472
rect 800 19656 50200 20192
rect 880 19376 50120 19656
rect 800 18840 50200 19376
rect 880 18560 50120 18840
rect 800 18024 50200 18560
rect 880 17744 50120 18024
rect 800 17208 50200 17744
rect 880 16928 50120 17208
rect 800 16392 50200 16928
rect 880 16112 50120 16392
rect 800 15576 50200 16112
rect 880 15296 50120 15576
rect 800 14760 50200 15296
rect 880 14480 50120 14760
rect 800 13944 50200 14480
rect 880 13664 50120 13944
rect 800 13128 50200 13664
rect 880 12848 50120 13128
rect 800 12312 50200 12848
rect 880 12032 50120 12312
rect 800 11496 50200 12032
rect 880 11216 50120 11496
rect 800 10680 50200 11216
rect 880 10400 50120 10680
rect 800 9864 50200 10400
rect 880 9584 50120 9864
rect 800 9048 50200 9584
rect 880 8768 50120 9048
rect 800 8232 50200 8768
rect 880 7952 50120 8232
rect 800 7416 50200 7952
rect 880 7136 50120 7416
rect 800 6600 50200 7136
rect 880 6320 50120 6600
rect 800 5784 50200 6320
rect 880 5504 50120 5784
rect 800 4968 50200 5504
rect 880 4688 50120 4968
rect 800 4152 50200 4688
rect 880 3872 50120 4152
rect 800 3336 50200 3872
rect 880 3056 50120 3336
rect 800 2520 50200 3056
rect 800 2240 50120 2520
rect 800 2143 50200 2240
<< metal4 >>
rect 2944 2128 3264 54448
rect 7944 2128 8264 54448
rect 12944 2128 13264 54448
rect 17944 2128 18264 54448
rect 22944 2128 23264 54448
rect 27944 2128 28264 54448
rect 32944 2128 33264 54448
rect 37944 2128 38264 54448
rect 42944 2128 43264 54448
rect 47944 2128 48264 54448
<< obsm4 >>
rect 18459 14315 22864 52053
rect 23344 14315 27864 52053
rect 28344 14315 32864 52053
rect 33344 14315 34165 52053
<< labels >>
rlabel metal4 s 7944 2128 8264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27944 2128 28264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37944 2128 38264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47944 2128 48264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 32944 2128 33264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 42944 2128 43264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 2226 0 2282 800 6 ccff_head
port 3 nsew signal input
rlabel metal2 s 49238 56200 49294 57000 6 ccff_head_1
port 4 nsew signal input
rlabel metal3 s 50200 2320 51000 2440 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 1582 56200 1638 57000 6 ccff_tail_0
port 6 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 chanx_left_in[0]
port 7 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[10]
port 8 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[11]
port 9 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[12]
port 10 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_in[13]
port 11 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 chanx_left_in[14]
port 12 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 chanx_left_in[15]
port 13 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 chanx_left_in[16]
port 14 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 chanx_left_in[17]
port 15 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 chanx_left_in[18]
port 16 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 chanx_left_in[19]
port 17 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[1]
port 18 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 chanx_left_in[20]
port 19 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 chanx_left_in[21]
port 20 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 chanx_left_in[22]
port 21 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 chanx_left_in[23]
port 22 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 chanx_left_in[24]
port 23 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 chanx_left_in[25]
port 24 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 chanx_left_in[26]
port 25 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 chanx_left_in[27]
port 26 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 chanx_left_in[28]
port 27 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 chanx_left_in[29]
port 28 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 29 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[3]
port 30 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 chanx_left_in[4]
port 31 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[5]
port 32 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[6]
port 33 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[7]
port 34 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[8]
port 35 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[9]
port 36 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 chanx_left_out[0]
port 37 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 chanx_left_out[10]
port 38 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 chanx_left_out[11]
port 39 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 chanx_left_out[12]
port 40 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 chanx_left_out[13]
port 41 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 chanx_left_out[14]
port 42 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 chanx_left_out[15]
port 43 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 chanx_left_out[16]
port 44 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 chanx_left_out[17]
port 45 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 chanx_left_out[18]
port 46 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 chanx_left_out[19]
port 47 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 chanx_left_out[1]
port 48 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 chanx_left_out[20]
port 49 nsew signal output
rlabel metal3 s 0 44752 800 44872 6 chanx_left_out[21]
port 50 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 chanx_left_out[22]
port 51 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 chanx_left_out[23]
port 52 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 chanx_left_out[24]
port 53 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 chanx_left_out[25]
port 54 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 chanx_left_out[26]
port 55 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 chanx_left_out[27]
port 56 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 chanx_left_out[28]
port 57 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 chanx_left_out[29]
port 58 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 chanx_left_out[2]
port 59 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 chanx_left_out[3]
port 60 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 chanx_left_out[4]
port 61 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 chanx_left_out[5]
port 62 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 chanx_left_out[6]
port 63 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 chanx_left_out[7]
port 64 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 chanx_left_out[8]
port 65 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 chanx_left_out[9]
port 66 nsew signal output
rlabel metal3 s 50200 27616 51000 27736 6 chanx_right_in_0[0]
port 67 nsew signal input
rlabel metal3 s 50200 35776 51000 35896 6 chanx_right_in_0[10]
port 68 nsew signal input
rlabel metal3 s 50200 36592 51000 36712 6 chanx_right_in_0[11]
port 69 nsew signal input
rlabel metal3 s 50200 37408 51000 37528 6 chanx_right_in_0[12]
port 70 nsew signal input
rlabel metal3 s 50200 38224 51000 38344 6 chanx_right_in_0[13]
port 71 nsew signal input
rlabel metal3 s 50200 39040 51000 39160 6 chanx_right_in_0[14]
port 72 nsew signal input
rlabel metal3 s 50200 39856 51000 39976 6 chanx_right_in_0[15]
port 73 nsew signal input
rlabel metal3 s 50200 40672 51000 40792 6 chanx_right_in_0[16]
port 74 nsew signal input
rlabel metal3 s 50200 41488 51000 41608 6 chanx_right_in_0[17]
port 75 nsew signal input
rlabel metal3 s 50200 42304 51000 42424 6 chanx_right_in_0[18]
port 76 nsew signal input
rlabel metal3 s 50200 43120 51000 43240 6 chanx_right_in_0[19]
port 77 nsew signal input
rlabel metal3 s 50200 28432 51000 28552 6 chanx_right_in_0[1]
port 78 nsew signal input
rlabel metal3 s 50200 43936 51000 44056 6 chanx_right_in_0[20]
port 79 nsew signal input
rlabel metal3 s 50200 44752 51000 44872 6 chanx_right_in_0[21]
port 80 nsew signal input
rlabel metal3 s 50200 45568 51000 45688 6 chanx_right_in_0[22]
port 81 nsew signal input
rlabel metal3 s 50200 46384 51000 46504 6 chanx_right_in_0[23]
port 82 nsew signal input
rlabel metal3 s 50200 47200 51000 47320 6 chanx_right_in_0[24]
port 83 nsew signal input
rlabel metal3 s 50200 48016 51000 48136 6 chanx_right_in_0[25]
port 84 nsew signal input
rlabel metal3 s 50200 48832 51000 48952 6 chanx_right_in_0[26]
port 85 nsew signal input
rlabel metal3 s 50200 49648 51000 49768 6 chanx_right_in_0[27]
port 86 nsew signal input
rlabel metal3 s 50200 50464 51000 50584 6 chanx_right_in_0[28]
port 87 nsew signal input
rlabel metal3 s 50200 51280 51000 51400 6 chanx_right_in_0[29]
port 88 nsew signal input
rlabel metal3 s 50200 29248 51000 29368 6 chanx_right_in_0[2]
port 89 nsew signal input
rlabel metal3 s 50200 30064 51000 30184 6 chanx_right_in_0[3]
port 90 nsew signal input
rlabel metal3 s 50200 30880 51000 31000 6 chanx_right_in_0[4]
port 91 nsew signal input
rlabel metal3 s 50200 31696 51000 31816 6 chanx_right_in_0[5]
port 92 nsew signal input
rlabel metal3 s 50200 32512 51000 32632 6 chanx_right_in_0[6]
port 93 nsew signal input
rlabel metal3 s 50200 33328 51000 33448 6 chanx_right_in_0[7]
port 94 nsew signal input
rlabel metal3 s 50200 34144 51000 34264 6 chanx_right_in_0[8]
port 95 nsew signal input
rlabel metal3 s 50200 34960 51000 35080 6 chanx_right_in_0[9]
port 96 nsew signal input
rlabel metal3 s 50200 3136 51000 3256 6 chanx_right_out_0[0]
port 97 nsew signal output
rlabel metal3 s 50200 11296 51000 11416 6 chanx_right_out_0[10]
port 98 nsew signal output
rlabel metal3 s 50200 12112 51000 12232 6 chanx_right_out_0[11]
port 99 nsew signal output
rlabel metal3 s 50200 12928 51000 13048 6 chanx_right_out_0[12]
port 100 nsew signal output
rlabel metal3 s 50200 13744 51000 13864 6 chanx_right_out_0[13]
port 101 nsew signal output
rlabel metal3 s 50200 14560 51000 14680 6 chanx_right_out_0[14]
port 102 nsew signal output
rlabel metal3 s 50200 15376 51000 15496 6 chanx_right_out_0[15]
port 103 nsew signal output
rlabel metal3 s 50200 16192 51000 16312 6 chanx_right_out_0[16]
port 104 nsew signal output
rlabel metal3 s 50200 17008 51000 17128 6 chanx_right_out_0[17]
port 105 nsew signal output
rlabel metal3 s 50200 17824 51000 17944 6 chanx_right_out_0[18]
port 106 nsew signal output
rlabel metal3 s 50200 18640 51000 18760 6 chanx_right_out_0[19]
port 107 nsew signal output
rlabel metal3 s 50200 3952 51000 4072 6 chanx_right_out_0[1]
port 108 nsew signal output
rlabel metal3 s 50200 19456 51000 19576 6 chanx_right_out_0[20]
port 109 nsew signal output
rlabel metal3 s 50200 20272 51000 20392 6 chanx_right_out_0[21]
port 110 nsew signal output
rlabel metal3 s 50200 21088 51000 21208 6 chanx_right_out_0[22]
port 111 nsew signal output
rlabel metal3 s 50200 21904 51000 22024 6 chanx_right_out_0[23]
port 112 nsew signal output
rlabel metal3 s 50200 22720 51000 22840 6 chanx_right_out_0[24]
port 113 nsew signal output
rlabel metal3 s 50200 23536 51000 23656 6 chanx_right_out_0[25]
port 114 nsew signal output
rlabel metal3 s 50200 24352 51000 24472 6 chanx_right_out_0[26]
port 115 nsew signal output
rlabel metal3 s 50200 25168 51000 25288 6 chanx_right_out_0[27]
port 116 nsew signal output
rlabel metal3 s 50200 25984 51000 26104 6 chanx_right_out_0[28]
port 117 nsew signal output
rlabel metal3 s 50200 26800 51000 26920 6 chanx_right_out_0[29]
port 118 nsew signal output
rlabel metal3 s 50200 4768 51000 4888 6 chanx_right_out_0[2]
port 119 nsew signal output
rlabel metal3 s 50200 5584 51000 5704 6 chanx_right_out_0[3]
port 120 nsew signal output
rlabel metal3 s 50200 6400 51000 6520 6 chanx_right_out_0[4]
port 121 nsew signal output
rlabel metal3 s 50200 7216 51000 7336 6 chanx_right_out_0[5]
port 122 nsew signal output
rlabel metal3 s 50200 8032 51000 8152 6 chanx_right_out_0[6]
port 123 nsew signal output
rlabel metal3 s 50200 8848 51000 8968 6 chanx_right_out_0[7]
port 124 nsew signal output
rlabel metal3 s 50200 9664 51000 9784 6 chanx_right_out_0[8]
port 125 nsew signal output
rlabel metal3 s 50200 10480 51000 10600 6 chanx_right_out_0[9]
port 126 nsew signal output
rlabel metal2 s 21546 56200 21602 57000 6 chany_top_in[0]
port 127 nsew signal input
rlabel metal2 s 27986 56200 28042 57000 6 chany_top_in[10]
port 128 nsew signal input
rlabel metal2 s 28630 56200 28686 57000 6 chany_top_in[11]
port 129 nsew signal input
rlabel metal2 s 29274 56200 29330 57000 6 chany_top_in[12]
port 130 nsew signal input
rlabel metal2 s 29918 56200 29974 57000 6 chany_top_in[13]
port 131 nsew signal input
rlabel metal2 s 30562 56200 30618 57000 6 chany_top_in[14]
port 132 nsew signal input
rlabel metal2 s 31206 56200 31262 57000 6 chany_top_in[15]
port 133 nsew signal input
rlabel metal2 s 31850 56200 31906 57000 6 chany_top_in[16]
port 134 nsew signal input
rlabel metal2 s 32494 56200 32550 57000 6 chany_top_in[17]
port 135 nsew signal input
rlabel metal2 s 33138 56200 33194 57000 6 chany_top_in[18]
port 136 nsew signal input
rlabel metal2 s 33782 56200 33838 57000 6 chany_top_in[19]
port 137 nsew signal input
rlabel metal2 s 22190 56200 22246 57000 6 chany_top_in[1]
port 138 nsew signal input
rlabel metal2 s 34426 56200 34482 57000 6 chany_top_in[20]
port 139 nsew signal input
rlabel metal2 s 35070 56200 35126 57000 6 chany_top_in[21]
port 140 nsew signal input
rlabel metal2 s 35714 56200 35770 57000 6 chany_top_in[22]
port 141 nsew signal input
rlabel metal2 s 36358 56200 36414 57000 6 chany_top_in[23]
port 142 nsew signal input
rlabel metal2 s 37002 56200 37058 57000 6 chany_top_in[24]
port 143 nsew signal input
rlabel metal2 s 37646 56200 37702 57000 6 chany_top_in[25]
port 144 nsew signal input
rlabel metal2 s 38290 56200 38346 57000 6 chany_top_in[26]
port 145 nsew signal input
rlabel metal2 s 38934 56200 38990 57000 6 chany_top_in[27]
port 146 nsew signal input
rlabel metal2 s 39578 56200 39634 57000 6 chany_top_in[28]
port 147 nsew signal input
rlabel metal2 s 40222 56200 40278 57000 6 chany_top_in[29]
port 148 nsew signal input
rlabel metal2 s 22834 56200 22890 57000 6 chany_top_in[2]
port 149 nsew signal input
rlabel metal2 s 23478 56200 23534 57000 6 chany_top_in[3]
port 150 nsew signal input
rlabel metal2 s 24122 56200 24178 57000 6 chany_top_in[4]
port 151 nsew signal input
rlabel metal2 s 24766 56200 24822 57000 6 chany_top_in[5]
port 152 nsew signal input
rlabel metal2 s 25410 56200 25466 57000 6 chany_top_in[6]
port 153 nsew signal input
rlabel metal2 s 26054 56200 26110 57000 6 chany_top_in[7]
port 154 nsew signal input
rlabel metal2 s 26698 56200 26754 57000 6 chany_top_in[8]
port 155 nsew signal input
rlabel metal2 s 27342 56200 27398 57000 6 chany_top_in[9]
port 156 nsew signal input
rlabel metal2 s 2226 56200 2282 57000 6 chany_top_out[0]
port 157 nsew signal output
rlabel metal2 s 8666 56200 8722 57000 6 chany_top_out[10]
port 158 nsew signal output
rlabel metal2 s 9310 56200 9366 57000 6 chany_top_out[11]
port 159 nsew signal output
rlabel metal2 s 9954 56200 10010 57000 6 chany_top_out[12]
port 160 nsew signal output
rlabel metal2 s 10598 56200 10654 57000 6 chany_top_out[13]
port 161 nsew signal output
rlabel metal2 s 11242 56200 11298 57000 6 chany_top_out[14]
port 162 nsew signal output
rlabel metal2 s 11886 56200 11942 57000 6 chany_top_out[15]
port 163 nsew signal output
rlabel metal2 s 12530 56200 12586 57000 6 chany_top_out[16]
port 164 nsew signal output
rlabel metal2 s 13174 56200 13230 57000 6 chany_top_out[17]
port 165 nsew signal output
rlabel metal2 s 13818 56200 13874 57000 6 chany_top_out[18]
port 166 nsew signal output
rlabel metal2 s 14462 56200 14518 57000 6 chany_top_out[19]
port 167 nsew signal output
rlabel metal2 s 2870 56200 2926 57000 6 chany_top_out[1]
port 168 nsew signal output
rlabel metal2 s 15106 56200 15162 57000 6 chany_top_out[20]
port 169 nsew signal output
rlabel metal2 s 15750 56200 15806 57000 6 chany_top_out[21]
port 170 nsew signal output
rlabel metal2 s 16394 56200 16450 57000 6 chany_top_out[22]
port 171 nsew signal output
rlabel metal2 s 17038 56200 17094 57000 6 chany_top_out[23]
port 172 nsew signal output
rlabel metal2 s 17682 56200 17738 57000 6 chany_top_out[24]
port 173 nsew signal output
rlabel metal2 s 18326 56200 18382 57000 6 chany_top_out[25]
port 174 nsew signal output
rlabel metal2 s 18970 56200 19026 57000 6 chany_top_out[26]
port 175 nsew signal output
rlabel metal2 s 19614 56200 19670 57000 6 chany_top_out[27]
port 176 nsew signal output
rlabel metal2 s 20258 56200 20314 57000 6 chany_top_out[28]
port 177 nsew signal output
rlabel metal2 s 20902 56200 20958 57000 6 chany_top_out[29]
port 178 nsew signal output
rlabel metal2 s 3514 56200 3570 57000 6 chany_top_out[2]
port 179 nsew signal output
rlabel metal2 s 4158 56200 4214 57000 6 chany_top_out[3]
port 180 nsew signal output
rlabel metal2 s 4802 56200 4858 57000 6 chany_top_out[4]
port 181 nsew signal output
rlabel metal2 s 5446 56200 5502 57000 6 chany_top_out[5]
port 182 nsew signal output
rlabel metal2 s 6090 56200 6146 57000 6 chany_top_out[6]
port 183 nsew signal output
rlabel metal2 s 6734 56200 6790 57000 6 chany_top_out[7]
port 184 nsew signal output
rlabel metal2 s 7378 56200 7434 57000 6 chany_top_out[8]
port 185 nsew signal output
rlabel metal2 s 8022 56200 8078 57000 6 chany_top_out[9]
port 186 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 gfpga_pad_io_soc_dir[0]
port 187 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 gfpga_pad_io_soc_dir[1]
port 188 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 gfpga_pad_io_soc_dir[2]
port 189 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 gfpga_pad_io_soc_dir[3]
port 190 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 gfpga_pad_io_soc_in[0]
port 191 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 gfpga_pad_io_soc_in[1]
port 192 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 gfpga_pad_io_soc_in[2]
port 193 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 gfpga_pad_io_soc_in[3]
port 194 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 gfpga_pad_io_soc_out[0]
port 195 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 gfpga_pad_io_soc_out[1]
port 196 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 gfpga_pad_io_soc_out[2]
port 197 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 gfpga_pad_io_soc_out[3]
port 198 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 isol_n
port 199 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 prog_clk
port 200 nsew signal input
rlabel metal2 s 42154 56200 42210 57000 6 prog_reset_top_in
port 201 nsew signal input
rlabel metal2 s 42798 56200 42854 57000 6 reset_top_in
port 202 nsew signal input
rlabel metal3 s 50200 52096 51000 52216 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 203 nsew signal input
rlabel metal3 s 50200 52912 51000 53032 6 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 204 nsew signal input
rlabel metal3 s 50200 53728 51000 53848 6 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 205 nsew signal input
rlabel metal3 s 50200 54544 51000 54664 6 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 206 nsew signal input
rlabel metal2 s 43442 56200 43498 57000 6 test_enable_top_in
port 207 nsew signal input
rlabel metal2 s 45374 56200 45430 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 208 nsew signal input
rlabel metal2 s 46018 56200 46074 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 209 nsew signal input
rlabel metal2 s 46662 56200 46718 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 210 nsew signal input
rlabel metal2 s 47306 56200 47362 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 211 nsew signal input
rlabel metal2 s 47950 56200 48006 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 212 nsew signal input
rlabel metal2 s 48594 56200 48650 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 213 nsew signal input
rlabel metal2 s 44086 56200 44142 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 214 nsew signal input
rlabel metal2 s 44730 56200 44786 57000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 215 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 top_width_0_height_0_subtile_0__pin_inpad_0_
port 216 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 top_width_0_height_0_subtile_1__pin_inpad_0_
port 217 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 top_width_0_height_0_subtile_2__pin_inpad_0_
port 218 nsew signal output
rlabel metal3 s 0 54544 800 54664 6 top_width_0_height_0_subtile_3__pin_inpad_0_
port 219 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 51000 57000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3050952
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/bottom_tile/runs/23_03_20_06_54/results/signoff/bottom_tile.magic.gds
string GDS_START 175904
<< end >>

