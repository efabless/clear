magic
tech sky130A
magscale 1 2
timestamp 1681685389
<< viali >>
rect 26433 24361 26467 24395
rect 29745 24361 29779 24395
rect 39313 24361 39347 24395
rect 42625 24361 42659 24395
rect 47593 24361 47627 24395
rect 24593 24293 24627 24327
rect 25789 24293 25823 24327
rect 27169 24293 27203 24327
rect 32965 24293 32999 24327
rect 38209 24293 38243 24327
rect 2973 24225 3007 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10701 24225 10735 24259
rect 13277 24225 13311 24259
rect 15853 24225 15887 24259
rect 18429 24225 18463 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25237 24225 25271 24259
rect 26617 24225 26651 24259
rect 29193 24225 29227 24259
rect 31493 24225 31527 24259
rect 31953 24225 31987 24259
rect 34253 24225 34287 24259
rect 34989 24225 35023 24259
rect 35173 24225 35207 24259
rect 36553 24225 36587 24259
rect 36737 24225 36771 24259
rect 37565 24225 37599 24259
rect 40601 24225 40635 24259
rect 45845 24225 45879 24259
rect 47225 24225 47259 24259
rect 3433 24157 3467 24191
rect 3985 24157 4019 24191
rect 4629 24157 4663 24191
rect 6561 24157 6595 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 11161 24157 11195 24191
rect 11897 24157 11931 24191
rect 13737 24157 13771 24191
rect 14473 24157 14507 24191
rect 16313 24157 16347 24191
rect 18889 24157 18923 24191
rect 19625 24157 19659 24191
rect 21373 24157 21407 24191
rect 22017 24157 22051 24191
rect 23857 24157 23891 24191
rect 27905 24157 27939 24191
rect 28549 24157 28583 24191
rect 29929 24157 29963 24191
rect 30389 24157 30423 24191
rect 31033 24157 31067 24191
rect 31677 24157 31711 24191
rect 32505 24157 32539 24191
rect 33149 24157 33183 24191
rect 37749 24157 37783 24191
rect 38853 24157 38887 24191
rect 39497 24157 39531 24191
rect 40417 24157 40451 24191
rect 42073 24157 42107 24191
rect 42809 24157 42843 24191
rect 43453 24157 43487 24191
rect 44373 24157 44407 24191
rect 45201 24157 45235 24191
rect 46949 24157 46983 24191
rect 48237 24157 48271 24191
rect 48973 24157 49007 24191
rect 49433 24157 49467 24191
rect 24961 24089 24995 24123
rect 25973 24089 26007 24123
rect 26801 24089 26835 24123
rect 27353 24089 27387 24123
rect 29009 24089 29043 24123
rect 33977 24089 34011 24123
rect 41061 24089 41095 24123
rect 43729 24089 43763 24123
rect 49249 24089 49283 24123
rect 4169 24021 4203 24055
rect 6745 24021 6779 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 14289 24021 14323 24055
rect 17049 24021 17083 24055
rect 19441 24021 19475 24055
rect 24041 24021 24075 24055
rect 25053 24021 25087 24055
rect 28089 24021 28123 24055
rect 28733 24021 28767 24055
rect 30573 24021 30607 24055
rect 31217 24021 31251 24055
rect 32321 24021 32355 24055
rect 33609 24021 33643 24055
rect 34069 24021 34103 24055
rect 35265 24021 35299 24055
rect 35633 24021 35667 24055
rect 36093 24021 36127 24055
rect 36461 24021 36495 24055
rect 37841 24021 37875 24055
rect 38669 24021 38703 24055
rect 40049 24021 40083 24055
rect 40509 24021 40543 24055
rect 41429 24021 41463 24055
rect 43269 24021 43303 24055
rect 44189 24021 44223 24055
rect 44649 24021 44683 24055
rect 46305 24021 46339 24055
rect 48053 24021 48087 24055
rect 48789 24021 48823 24055
rect 2329 23817 2363 23851
rect 7481 23817 7515 23851
rect 21465 23817 21499 23851
rect 28457 23817 28491 23851
rect 32321 23817 32355 23851
rect 32781 23817 32815 23851
rect 37473 23817 37507 23851
rect 37841 23817 37875 23851
rect 44649 23817 44683 23851
rect 47593 23817 47627 23851
rect 49157 23817 49191 23851
rect 49525 23817 49559 23851
rect 14289 23749 14323 23783
rect 20269 23749 20303 23783
rect 24501 23749 24535 23783
rect 26341 23749 26375 23783
rect 31493 23749 31527 23783
rect 37933 23749 37967 23783
rect 39221 23749 39255 23783
rect 39313 23749 39347 23783
rect 42441 23749 42475 23783
rect 43361 23749 43395 23783
rect 2145 23681 2179 23715
rect 4077 23681 4111 23715
rect 4721 23681 4755 23715
rect 6837 23681 6871 23715
rect 7297 23681 7331 23715
rect 9321 23681 9355 23715
rect 11161 23681 11195 23715
rect 13093 23681 13127 23715
rect 16313 23681 16347 23715
rect 18245 23681 18279 23715
rect 21281 23681 21315 23715
rect 22845 23681 22879 23715
rect 23673 23681 23707 23715
rect 24409 23681 24443 23715
rect 27353 23681 27387 23715
rect 27813 23681 27847 23715
rect 28641 23681 28675 23715
rect 29101 23681 29135 23715
rect 29561 23681 29595 23715
rect 32689 23681 32723 23715
rect 36277 23681 36311 23715
rect 42073 23681 42107 23715
rect 44189 23681 44223 23715
rect 44833 23681 44867 23715
rect 45937 23681 45971 23715
rect 46397 23681 46431 23715
rect 47317 23681 47351 23715
rect 48789 23681 48823 23715
rect 3709 23613 3743 23647
rect 5457 23613 5491 23647
rect 8861 23613 8895 23647
rect 10609 23613 10643 23647
rect 12357 23613 12391 23647
rect 12633 23613 12667 23647
rect 15853 23613 15887 23647
rect 17877 23613 17911 23647
rect 20545 23613 20579 23647
rect 22569 23613 22603 23647
rect 23765 23613 23799 23647
rect 23857 23613 23891 23647
rect 26617 23613 26651 23647
rect 31769 23613 31803 23647
rect 32965 23613 32999 23647
rect 35357 23613 35391 23647
rect 36369 23613 36403 23647
rect 36461 23613 36495 23647
rect 38025 23613 38059 23647
rect 39405 23613 39439 23647
rect 39957 23613 39991 23647
rect 40325 23613 40359 23647
rect 43177 23613 43211 23647
rect 47041 23613 47075 23647
rect 35909 23545 35943 23579
rect 36921 23545 36955 23579
rect 38853 23545 38887 23579
rect 42993 23545 43027 23579
rect 43545 23545 43579 23579
rect 44005 23545 44039 23579
rect 48145 23545 48179 23579
rect 6653 23477 6687 23511
rect 18797 23477 18831 23511
rect 20913 23477 20947 23511
rect 23305 23477 23339 23511
rect 24869 23477 24903 23511
rect 27169 23477 27203 23511
rect 27997 23477 28031 23511
rect 29285 23477 29319 23511
rect 30021 23477 30055 23511
rect 33609 23477 33643 23511
rect 35099 23477 35133 23511
rect 38577 23477 38611 23511
rect 42625 23477 42659 23511
rect 42901 23477 42935 23511
rect 45293 23477 45327 23511
rect 47869 23477 47903 23511
rect 49341 23477 49375 23511
rect 4721 23273 4755 23307
rect 27905 23273 27939 23307
rect 29009 23273 29043 23307
rect 29193 23273 29227 23307
rect 29745 23273 29779 23307
rect 34161 23273 34195 23307
rect 39313 23273 39347 23307
rect 44649 23273 44683 23307
rect 48237 23273 48271 23307
rect 19625 23205 19659 23239
rect 20361 23205 20395 23239
rect 24593 23205 24627 23239
rect 25237 23205 25271 23239
rect 34345 23205 34379 23239
rect 45937 23205 45971 23239
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 10057 23137 10091 23171
rect 11253 23137 11287 23171
rect 13277 23137 13311 23171
rect 15761 23137 15795 23171
rect 18613 23137 18647 23171
rect 19349 23137 19383 23171
rect 22109 23137 22143 23171
rect 23949 23137 23983 23171
rect 25973 23137 26007 23171
rect 28457 23137 28491 23171
rect 30205 23137 30239 23171
rect 30297 23137 30331 23171
rect 30849 23137 30883 23171
rect 31401 23137 31435 23171
rect 33149 23137 33183 23171
rect 35357 23137 35391 23171
rect 37289 23137 37323 23171
rect 39037 23137 39071 23171
rect 39497 23137 39531 23171
rect 40601 23137 40635 23171
rect 41061 23137 41095 23171
rect 43545 23137 43579 23171
rect 45753 23137 45787 23171
rect 2973 23069 3007 23103
rect 4261 23069 4295 23103
rect 4905 23069 4939 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9321 23069 9355 23103
rect 11897 23069 11931 23103
rect 13737 23069 13771 23103
rect 14841 23069 14875 23103
rect 16681 23069 16715 23103
rect 18889 23069 18923 23103
rect 23765 23069 23799 23103
rect 25697 23069 25731 23103
rect 28273 23069 28307 23103
rect 33885 23069 33919 23103
rect 35081 23069 35115 23103
rect 41521 23069 41555 23103
rect 44005 23069 44039 23103
rect 45201 23069 45235 23103
rect 45385 23069 45419 23103
rect 47133 23069 47167 23103
rect 47593 23069 47627 23103
rect 49341 23069 49375 23103
rect 1777 23001 1811 23035
rect 19809 23001 19843 23035
rect 21833 23001 21867 23035
rect 22569 23001 22603 23035
rect 22753 23001 22787 23035
rect 24777 23001 24811 23035
rect 28365 23001 28399 23035
rect 31677 23001 31711 23035
rect 38761 23001 38795 23035
rect 40417 23001 40451 23035
rect 43269 23001 43303 23035
rect 46121 23001 46155 23035
rect 4077 22933 4111 22967
rect 9229 22933 9263 22967
rect 14197 22933 14231 22967
rect 14381 22933 14415 22967
rect 14657 22933 14691 22967
rect 17141 22933 17175 22967
rect 23305 22933 23339 22967
rect 23673 22933 23707 22967
rect 25329 22933 25363 22967
rect 27445 22933 27479 22967
rect 29377 22933 29411 22967
rect 30113 22933 30147 22967
rect 31033 22933 31067 22967
rect 33701 22933 33735 22967
rect 34713 22933 34747 22967
rect 36829 22933 36863 22967
rect 40049 22933 40083 22967
rect 40509 22933 40543 22967
rect 46489 22933 46523 22967
rect 48697 22933 48731 22967
rect 9505 22729 9539 22763
rect 14565 22729 14599 22763
rect 19073 22729 19107 22763
rect 21189 22729 21223 22763
rect 27353 22729 27387 22763
rect 32321 22729 32355 22763
rect 32689 22729 32723 22763
rect 35449 22729 35483 22763
rect 35817 22729 35851 22763
rect 37473 22729 37507 22763
rect 43269 22729 43303 22763
rect 46581 22729 46615 22763
rect 4813 22661 4847 22695
rect 9965 22661 9999 22695
rect 12817 22661 12851 22695
rect 15117 22661 15151 22695
rect 18981 22661 19015 22695
rect 22293 22661 22327 22695
rect 24133 22661 24167 22695
rect 26341 22661 26375 22695
rect 29561 22661 29595 22695
rect 33977 22661 34011 22695
rect 45201 22661 45235 22695
rect 45753 22661 45787 22695
rect 45937 22661 45971 22695
rect 47961 22661 47995 22695
rect 2973 22593 3007 22627
rect 3985 22593 4019 22627
rect 6009 22593 6043 22627
rect 6653 22593 6687 22627
rect 7481 22593 7515 22627
rect 11161 22593 11195 22627
rect 11897 22593 11931 22627
rect 14013 22593 14047 22627
rect 16313 22593 16347 22627
rect 16865 22593 16899 22627
rect 19441 22593 19475 22627
rect 22017 22593 22051 22627
rect 24409 22593 24443 22627
rect 27169 22593 27203 22627
rect 27721 22593 27755 22627
rect 30665 22593 30699 22627
rect 30757 22593 30791 22627
rect 31677 22593 31711 22627
rect 32781 22593 32815 22627
rect 33701 22593 33735 22627
rect 36461 22593 36495 22627
rect 39221 22593 39255 22627
rect 39497 22593 39531 22627
rect 39773 22593 39807 22627
rect 40417 22593 40451 22627
rect 40509 22593 40543 22627
rect 41429 22593 41463 22627
rect 42073 22593 42107 22627
rect 42625 22593 42659 22627
rect 47225 22593 47259 22627
rect 49341 22593 49375 22627
rect 2513 22525 2547 22559
rect 7113 22525 7147 22559
rect 7941 22525 7975 22559
rect 17141 22525 17175 22559
rect 19717 22525 19751 22559
rect 26617 22525 26651 22559
rect 29837 22525 29871 22559
rect 30849 22525 30883 22559
rect 32873 22525 32907 22559
rect 36553 22525 36587 22559
rect 36737 22525 36771 22559
rect 38945 22525 38979 22559
rect 40601 22525 40635 22559
rect 43729 22525 43763 22559
rect 44005 22525 44039 22559
rect 48697 22525 48731 22559
rect 4169 22457 4203 22491
rect 6837 22457 6871 22491
rect 11713 22457 11747 22491
rect 24869 22457 24903 22491
rect 28089 22457 28123 22491
rect 36093 22457 36127 22491
rect 41245 22457 41279 22491
rect 45017 22457 45051 22491
rect 48329 22457 48363 22491
rect 9321 22389 9355 22423
rect 12265 22389 12299 22423
rect 14473 22389 14507 22423
rect 18613 22389 18647 22423
rect 21649 22389 21683 22423
rect 23765 22389 23799 22423
rect 24593 22389 24627 22423
rect 30297 22389 30331 22423
rect 31493 22389 31527 22423
rect 33425 22389 33459 22423
rect 40049 22389 40083 22423
rect 41889 22389 41923 22423
rect 47869 22389 47903 22423
rect 12357 22185 12391 22219
rect 15209 22185 15243 22219
rect 28365 22185 28399 22219
rect 34253 22185 34287 22219
rect 39405 22185 39439 22219
rect 39589 22185 39623 22219
rect 40233 22185 40267 22219
rect 44741 22185 44775 22219
rect 47225 22185 47259 22219
rect 14197 22117 14231 22151
rect 29745 22117 29779 22151
rect 36829 22117 36863 22151
rect 39865 22117 39899 22151
rect 6009 22049 6043 22083
rect 9781 22049 9815 22083
rect 11897 22049 11931 22083
rect 13645 22049 13679 22083
rect 17601 22049 17635 22083
rect 19901 22049 19935 22083
rect 22017 22049 22051 22083
rect 23213 22049 23247 22083
rect 25145 22049 25179 22083
rect 26525 22049 26559 22083
rect 27721 22049 27755 22083
rect 28917 22049 28951 22083
rect 33517 22049 33551 22083
rect 33701 22049 33735 22083
rect 35081 22049 35115 22083
rect 36277 22049 36311 22083
rect 39129 22049 39163 22083
rect 40693 22049 40727 22083
rect 40877 22049 40911 22083
rect 42073 22049 42107 22083
rect 42533 22049 42567 22083
rect 43085 22049 43119 22083
rect 44373 22049 44407 22083
rect 44557 22049 44591 22083
rect 45201 22049 45235 22083
rect 47041 22049 47075 22083
rect 47593 22049 47627 22083
rect 2973 21981 3007 22015
rect 5365 21981 5399 22015
rect 7205 21981 7239 22015
rect 7849 21981 7883 22015
rect 8585 21981 8619 22015
rect 9137 21981 9171 22015
rect 11621 21981 11655 22015
rect 12541 21981 12575 22015
rect 14473 21981 14507 22015
rect 16957 21981 16991 22015
rect 18797 21981 18831 22015
rect 19441 21981 19475 22015
rect 21189 21981 21223 22015
rect 23029 21981 23063 22015
rect 24041 21981 24075 22015
rect 25697 21981 25731 22015
rect 26433 21981 26467 22015
rect 29929 21981 29963 22015
rect 30849 21981 30883 22015
rect 36461 21981 36495 22015
rect 43361 21981 43395 22015
rect 44189 21981 44223 22015
rect 45477 21981 45511 22015
rect 46765 21981 46799 22015
rect 48237 21981 48271 22015
rect 49341 21981 49375 22015
rect 1777 21913 1811 21947
rect 4169 21913 4203 21947
rect 7665 21913 7699 21947
rect 14657 21913 14691 21947
rect 16681 21913 16715 21947
rect 21833 21913 21867 21947
rect 21925 21913 21959 21947
rect 24961 21913 24995 21947
rect 26341 21913 26375 21947
rect 27537 21913 27571 21947
rect 28733 21913 28767 21947
rect 28825 21913 28859 21947
rect 31125 21913 31159 21947
rect 34069 21913 34103 21947
rect 34437 21913 34471 21947
rect 38853 21913 38887 21947
rect 41797 21913 41831 21947
rect 8401 21845 8435 21879
rect 13001 21845 13035 21879
rect 13369 21845 13403 21879
rect 13461 21845 13495 21879
rect 21465 21845 21499 21879
rect 22661 21845 22695 21879
rect 23121 21845 23155 21879
rect 23857 21845 23891 21879
rect 24593 21845 24627 21879
rect 25053 21845 25087 21879
rect 25973 21845 26007 21879
rect 27169 21845 27203 21879
rect 27629 21845 27663 21879
rect 30205 21845 30239 21879
rect 30389 21845 30423 21879
rect 32597 21845 32631 21879
rect 33057 21845 33091 21879
rect 33425 21845 33459 21879
rect 35173 21845 35207 21879
rect 35265 21845 35299 21879
rect 35633 21845 35667 21879
rect 36369 21845 36403 21879
rect 37381 21845 37415 21879
rect 40601 21845 40635 21879
rect 41429 21845 41463 21879
rect 41889 21845 41923 21879
rect 42717 21845 42751 21879
rect 46581 21845 46615 21879
rect 48697 21845 48731 21879
rect 10517 21641 10551 21675
rect 11713 21641 11747 21675
rect 13185 21641 13219 21675
rect 13921 21641 13955 21675
rect 17417 21641 17451 21675
rect 17877 21641 17911 21675
rect 26433 21641 26467 21675
rect 28365 21641 28399 21675
rect 31125 21641 31159 21675
rect 32781 21641 32815 21675
rect 33609 21641 33643 21675
rect 34805 21641 34839 21675
rect 36093 21641 36127 21675
rect 42625 21641 42659 21675
rect 3617 21573 3651 21607
rect 14841 21573 14875 21607
rect 16773 21573 16807 21607
rect 21189 21573 21223 21607
rect 21373 21573 21407 21607
rect 27537 21573 27571 21607
rect 37289 21573 37323 21607
rect 40325 21573 40359 21607
rect 40417 21573 40451 21607
rect 40601 21573 40635 21607
rect 45293 21573 45327 21607
rect 45477 21573 45511 21607
rect 47133 21573 47167 21607
rect 2973 21505 3007 21539
rect 4629 21505 4663 21539
rect 5733 21505 5767 21539
rect 6561 21505 6595 21539
rect 8401 21505 8435 21539
rect 10701 21505 10735 21539
rect 12355 21505 12389 21539
rect 13277 21505 13311 21539
rect 14105 21505 14139 21539
rect 17785 21505 17819 21539
rect 25145 21505 25179 21539
rect 26617 21505 26651 21539
rect 28733 21505 28767 21539
rect 29929 21505 29963 21539
rect 30021 21505 30055 21539
rect 31217 21505 31251 21539
rect 33517 21505 33551 21539
rect 34713 21505 34747 21539
rect 37565 21505 37599 21539
rect 42809 21505 42843 21539
rect 43453 21505 43487 21539
rect 43913 21505 43947 21539
rect 45845 21505 45879 21539
rect 46397 21505 46431 21539
rect 47961 21505 47995 21539
rect 49341 21505 49375 21539
rect 1777 21437 1811 21471
rect 7021 21437 7055 21471
rect 8861 21437 8895 21471
rect 10241 21437 10275 21471
rect 12173 21437 12207 21471
rect 14565 21437 14599 21471
rect 18061 21437 18095 21471
rect 18613 21437 18647 21471
rect 18889 21437 18923 21471
rect 22477 21437 22511 21471
rect 22753 21437 22787 21471
rect 25237 21437 25271 21471
rect 25421 21437 25455 21471
rect 26065 21437 26099 21471
rect 27629 21437 27663 21471
rect 27721 21437 27755 21471
rect 28825 21437 28859 21471
rect 28917 21437 28951 21471
rect 30205 21437 30239 21471
rect 31401 21437 31435 21471
rect 31769 21437 31803 21471
rect 33333 21437 33367 21471
rect 34621 21437 34655 21471
rect 36185 21437 36219 21471
rect 36277 21437 36311 21471
rect 37013 21437 37047 21471
rect 38025 21437 38059 21471
rect 38301 21437 38335 21471
rect 39773 21437 39807 21471
rect 41245 21437 41279 21471
rect 41521 21437 41555 21471
rect 44189 21437 44223 21471
rect 46213 21437 46247 21471
rect 47777 21437 47811 21471
rect 5917 21369 5951 21403
rect 11161 21369 11195 21403
rect 11897 21369 11931 21403
rect 17141 21369 17175 21403
rect 20361 21369 20395 21403
rect 24777 21369 24811 21403
rect 40049 21369 40083 21403
rect 46949 21369 46983 21403
rect 48697 21369 48731 21403
rect 11345 21301 11379 21335
rect 12817 21301 12851 21335
rect 16313 21301 16347 21335
rect 16957 21301 16991 21335
rect 20637 21301 20671 21335
rect 20821 21301 20855 21335
rect 21925 21301 21959 21335
rect 22201 21301 22235 21335
rect 24225 21301 24259 21335
rect 25881 21301 25915 21335
rect 27169 21301 27203 21335
rect 29561 21301 29595 21335
rect 30757 21301 30791 21335
rect 33977 21301 34011 21335
rect 35173 21301 35207 21335
rect 35725 21301 35759 21335
rect 36737 21301 36771 21335
rect 37657 21301 37691 21335
rect 40877 21301 40911 21335
rect 43269 21301 43303 21335
rect 48329 21301 48363 21335
rect 14289 21097 14323 21131
rect 19993 21097 20027 21131
rect 24041 21097 24075 21131
rect 24777 21097 24811 21131
rect 29745 21097 29779 21131
rect 30849 21097 30883 21131
rect 37657 21097 37691 21131
rect 42809 21097 42843 21131
rect 44097 21097 44131 21131
rect 44465 21097 44499 21131
rect 45201 21097 45235 21131
rect 45845 21097 45879 21131
rect 9229 21029 9263 21063
rect 12725 21029 12759 21063
rect 21189 21029 21223 21063
rect 23397 21029 23431 21063
rect 29101 21029 29135 21063
rect 30297 21029 30331 21063
rect 42625 21029 42659 21063
rect 43913 21029 43947 21063
rect 44741 21029 44775 21063
rect 46581 21029 46615 21063
rect 2513 20961 2547 20995
rect 4169 20961 4203 20995
rect 6009 20961 6043 20995
rect 10057 20961 10091 20995
rect 16681 20961 16715 20995
rect 18613 20961 18647 20995
rect 20545 20961 20579 20995
rect 22661 20961 22695 20995
rect 25329 20961 25363 20995
rect 26157 20961 26191 20995
rect 26249 20961 26283 20995
rect 26709 20961 26743 20995
rect 27905 20961 27939 20995
rect 28549 20961 28583 20995
rect 31309 20961 31343 20995
rect 31493 20961 31527 20995
rect 32781 20961 32815 20995
rect 34253 20961 34287 20995
rect 36369 20961 36403 20995
rect 39405 20961 39439 20995
rect 40601 20961 40635 20995
rect 41797 20961 41831 20995
rect 42441 20961 42475 20995
rect 2973 20893 3007 20927
rect 5365 20893 5399 20927
rect 7205 20893 7239 20927
rect 8033 20893 8067 20927
rect 8401 20893 8435 20927
rect 9413 20893 9447 20927
rect 11345 20893 11379 20927
rect 11989 20893 12023 20927
rect 13737 20893 13771 20927
rect 16037 20893 16071 20927
rect 18889 20893 18923 20927
rect 20361 20893 20395 20927
rect 22937 20893 22971 20927
rect 24593 20893 24627 20927
rect 26065 20893 26099 20927
rect 26893 20893 26927 20927
rect 28641 20893 28675 20927
rect 28733 20893 28767 20927
rect 29929 20893 29963 20927
rect 32505 20893 32539 20927
rect 36645 20893 36679 20927
rect 40509 20893 40543 20927
rect 43453 20893 43487 20927
rect 43729 20893 43763 20927
rect 45385 20893 45419 20927
rect 46029 20893 46063 20927
rect 46765 20893 46799 20927
rect 47501 20893 47535 20927
rect 48237 20893 48271 20927
rect 48697 20893 48731 20927
rect 49341 20893 49375 20927
rect 12357 20825 12391 20859
rect 12909 20825 12943 20859
rect 15761 20825 15795 20859
rect 20453 20825 20487 20859
rect 23581 20825 23615 20859
rect 24225 20825 24259 20859
rect 25145 20825 25179 20859
rect 27353 20825 27387 20859
rect 31953 20825 31987 20859
rect 37197 20825 37231 20859
rect 39129 20825 39163 20859
rect 40417 20825 40451 20859
rect 41613 20825 41647 20859
rect 44649 20825 44683 20859
rect 7481 20757 7515 20791
rect 7849 20757 7883 20791
rect 10701 20757 10735 20791
rect 11161 20757 11195 20791
rect 11897 20757 11931 20791
rect 13553 20757 13587 20791
rect 17141 20757 17175 20791
rect 19349 20757 19383 20791
rect 19533 20757 19567 20791
rect 19625 20757 19659 20791
rect 25697 20757 25731 20791
rect 30389 20757 30423 20791
rect 31217 20757 31251 20791
rect 34897 20757 34931 20791
rect 36921 20757 36955 20791
rect 37289 20757 37323 20791
rect 40049 20757 40083 20791
rect 41245 20757 41279 20791
rect 41705 20757 41739 20791
rect 42257 20757 42291 20791
rect 43269 20757 43303 20791
rect 47317 20757 47351 20791
rect 48053 20757 48087 20791
rect 5457 20553 5491 20587
rect 9689 20553 9723 20587
rect 10333 20553 10367 20587
rect 14105 20553 14139 20587
rect 14933 20553 14967 20587
rect 15577 20553 15611 20587
rect 15945 20553 15979 20587
rect 16037 20553 16071 20587
rect 18797 20553 18831 20587
rect 19717 20553 19751 20587
rect 35265 20553 35299 20587
rect 40233 20553 40267 20587
rect 41797 20553 41831 20587
rect 45201 20553 45235 20587
rect 46305 20553 46339 20587
rect 46489 20553 46523 20587
rect 47685 20553 47719 20587
rect 3617 20485 3651 20519
rect 11161 20485 11195 20519
rect 22385 20485 22419 20519
rect 24133 20485 24167 20519
rect 29745 20485 29779 20519
rect 31033 20485 31067 20519
rect 36553 20485 36587 20519
rect 41153 20485 41187 20519
rect 47961 20485 47995 20519
rect 2973 20417 3007 20451
rect 4813 20417 4847 20451
rect 5273 20417 5307 20451
rect 6561 20417 6595 20451
rect 9229 20417 9263 20451
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 11897 20417 11931 20451
rect 12633 20417 12667 20451
rect 13093 20417 13127 20451
rect 13277 20417 13311 20451
rect 15117 20417 15151 20451
rect 17049 20417 17083 20451
rect 19073 20417 19107 20451
rect 21465 20417 21499 20451
rect 23397 20417 23431 20451
rect 23857 20417 23891 20451
rect 26065 20417 26099 20451
rect 27261 20417 27295 20451
rect 29837 20417 29871 20451
rect 31125 20417 31159 20451
rect 34897 20417 34931 20451
rect 36461 20417 36495 20451
rect 39497 20417 39531 20451
rect 40325 20417 40359 20451
rect 41613 20417 41647 20451
rect 45385 20417 45419 20451
rect 46029 20417 46063 20451
rect 47225 20417 47259 20451
rect 48145 20417 48179 20451
rect 48697 20417 48731 20451
rect 49341 20417 49375 20451
rect 2513 20349 2547 20383
rect 7021 20349 7055 20383
rect 14197 20349 14231 20383
rect 14289 20349 14323 20383
rect 16221 20349 16255 20383
rect 17325 20349 17359 20383
rect 21189 20349 21223 20383
rect 22477 20349 22511 20383
rect 22569 20349 22603 20383
rect 25605 20349 25639 20383
rect 27537 20349 27571 20383
rect 29561 20349 29595 20383
rect 31217 20349 31251 20383
rect 31953 20349 31987 20383
rect 32321 20349 32355 20383
rect 33793 20349 33827 20383
rect 34069 20349 34103 20383
rect 34713 20349 34747 20383
rect 34805 20349 34839 20383
rect 35725 20349 35759 20383
rect 36737 20349 36771 20383
rect 39221 20349 39255 20383
rect 40141 20349 40175 20383
rect 13737 20281 13771 20315
rect 23213 20281 23247 20315
rect 26617 20281 26651 20315
rect 29009 20281 29043 20315
rect 44925 20281 44959 20315
rect 9045 20213 9079 20247
rect 11805 20213 11839 20247
rect 12541 20213 12575 20247
rect 13461 20213 13495 20247
rect 16773 20213 16807 20247
rect 19349 20213 19383 20247
rect 22017 20213 22051 20247
rect 26249 20213 26283 20247
rect 30205 20213 30239 20247
rect 30665 20213 30699 20247
rect 31769 20213 31803 20247
rect 35541 20213 35575 20247
rect 36093 20213 36127 20247
rect 37381 20213 37415 20247
rect 37749 20213 37783 20247
rect 40693 20213 40727 20247
rect 45845 20213 45879 20247
rect 47041 20213 47075 20247
rect 14473 20009 14507 20043
rect 16865 20009 16899 20043
rect 18153 20009 18187 20043
rect 19349 20009 19383 20043
rect 20269 20009 20303 20043
rect 24041 20009 24075 20043
rect 25237 20009 25271 20043
rect 25605 20009 25639 20043
rect 31677 20009 31711 20043
rect 39589 20009 39623 20043
rect 41061 20009 41095 20043
rect 46213 20009 46247 20043
rect 47317 20009 47351 20043
rect 11253 19941 11287 19975
rect 14933 19941 14967 19975
rect 22753 19941 22787 19975
rect 25145 19941 25179 19975
rect 29377 19941 29411 19975
rect 34161 19941 34195 19975
rect 46673 19941 46707 19975
rect 4261 19873 4295 19907
rect 6009 19873 6043 19907
rect 11989 19873 12023 19907
rect 16313 19873 16347 19907
rect 17509 19873 17543 19907
rect 18797 19873 18831 19907
rect 22293 19873 22327 19907
rect 23489 19873 23523 19907
rect 24593 19873 24627 19907
rect 26065 19873 26099 19907
rect 26249 19873 26283 19907
rect 27353 19873 27387 19907
rect 28549 19873 28583 19907
rect 30297 19873 30331 19907
rect 31125 19873 31159 19907
rect 32689 19873 32723 19907
rect 33609 19873 33643 19907
rect 33701 19873 33735 19907
rect 35081 19873 35115 19907
rect 35173 19873 35207 19907
rect 36645 19873 36679 19907
rect 37933 19873 37967 19907
rect 39037 19873 39071 19907
rect 40141 19873 40175 19907
rect 40325 19873 40359 19907
rect 41245 19873 41279 19907
rect 45753 19873 45787 19907
rect 2973 19805 3007 19839
rect 5365 19805 5399 19839
rect 7205 19805 7239 19839
rect 7941 19805 7975 19839
rect 10149 19805 10183 19839
rect 10793 19805 10827 19839
rect 14289 19805 14323 19839
rect 16129 19805 16163 19839
rect 18521 19805 18555 19839
rect 23673 19805 23707 19839
rect 25973 19805 26007 19839
rect 27261 19805 27295 19839
rect 28365 19805 28399 19839
rect 30113 19805 30147 19839
rect 31217 19805 31251 19839
rect 32505 19805 32539 19839
rect 33793 19805 33827 19839
rect 35265 19805 35299 19839
rect 38117 19805 38151 19839
rect 38209 19805 38243 19839
rect 38853 19805 38887 19839
rect 40417 19805 40451 19839
rect 46029 19805 46063 19839
rect 46857 19805 46891 19839
rect 47501 19805 47535 19839
rect 49341 19805 49375 19839
rect 1777 19737 1811 19771
rect 9689 19737 9723 19771
rect 11437 19737 11471 19771
rect 12265 19737 12299 19771
rect 15117 19737 15151 19771
rect 16037 19737 16071 19771
rect 19809 19737 19843 19771
rect 22017 19737 22051 19771
rect 29009 19737 29043 19771
rect 32597 19737 32631 19771
rect 36461 19737 36495 19771
rect 47961 19737 47995 19771
rect 48145 19737 48179 19771
rect 48697 19737 48731 19771
rect 7757 19669 7791 19703
rect 9965 19669 9999 19703
rect 10609 19669 10643 19703
rect 13737 19669 13771 19703
rect 15669 19669 15703 19703
rect 17233 19669 17267 19703
rect 17325 19669 17359 19703
rect 18613 19669 18647 19703
rect 19717 19669 19751 19703
rect 20545 19669 20579 19703
rect 22661 19669 22695 19703
rect 23029 19669 23063 19703
rect 23581 19669 23615 19703
rect 26801 19669 26835 19703
rect 27169 19669 27203 19703
rect 27997 19669 28031 19703
rect 28457 19669 28491 19703
rect 29745 19669 29779 19703
rect 30205 19669 30239 19703
rect 31309 19669 31343 19703
rect 32137 19669 32171 19703
rect 34437 19669 34471 19703
rect 35633 19669 35667 19703
rect 36093 19669 36127 19703
rect 36553 19669 36587 19703
rect 37197 19669 37231 19703
rect 37381 19669 37415 19703
rect 37565 19669 37599 19703
rect 38577 19669 38611 19703
rect 40785 19669 40819 19703
rect 10977 19465 11011 19499
rect 15393 19465 15427 19499
rect 16865 19465 16899 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 28457 19465 28491 19499
rect 32689 19465 32723 19499
rect 33057 19465 33091 19499
rect 34253 19465 34287 19499
rect 35081 19465 35115 19499
rect 35449 19465 35483 19499
rect 37289 19465 37323 19499
rect 40141 19465 40175 19499
rect 40509 19465 40543 19499
rect 47041 19465 47075 19499
rect 47685 19465 47719 19499
rect 3617 19397 3651 19431
rect 10517 19397 10551 19431
rect 18061 19397 18095 19431
rect 22109 19397 22143 19431
rect 22937 19397 22971 19431
rect 26157 19397 26191 19431
rect 31493 19397 31527 19431
rect 32597 19397 32631 19431
rect 33793 19397 33827 19431
rect 36185 19397 36219 19431
rect 46397 19397 46431 19431
rect 1777 19329 1811 19363
rect 2973 19329 3007 19363
rect 4813 19329 4847 19363
rect 5457 19329 5491 19363
rect 11161 19329 11195 19363
rect 11713 19329 11747 19363
rect 12173 19329 12207 19363
rect 14473 19329 14507 19363
rect 15485 19329 15519 19363
rect 16221 19329 16255 19363
rect 17233 19329 17267 19363
rect 17325 19329 17359 19363
rect 21097 19329 21131 19363
rect 25237 19329 25271 19363
rect 26249 19329 26283 19363
rect 27629 19329 27663 19363
rect 28825 19329 28859 19363
rect 29745 19329 29779 19363
rect 30757 19329 30791 19363
rect 33885 19329 33919 19363
rect 36277 19329 36311 19363
rect 40601 19329 40635 19363
rect 41337 19329 41371 19363
rect 47225 19329 47259 19363
rect 48145 19329 48179 19363
rect 48697 19329 48731 19363
rect 49341 19329 49375 19363
rect 5273 19261 5307 19295
rect 9873 19261 9907 19295
rect 14197 19261 14231 19295
rect 14841 19261 14875 19295
rect 17417 19261 17451 19295
rect 19809 19261 19843 19295
rect 20085 19261 20119 19295
rect 21373 19261 21407 19295
rect 24961 19261 24995 19295
rect 26341 19261 26375 19295
rect 27721 19261 27755 19295
rect 27813 19261 27847 19295
rect 28917 19261 28951 19295
rect 29101 19261 29135 19295
rect 30389 19261 30423 19295
rect 32413 19261 32447 19295
rect 33701 19261 33735 19295
rect 34897 19261 34931 19295
rect 34989 19261 35023 19295
rect 36001 19261 36035 19295
rect 37565 19261 37599 19295
rect 39405 19261 39439 19295
rect 39681 19261 39715 19295
rect 40693 19261 40727 19295
rect 46581 19261 46615 19295
rect 11989 19193 12023 19227
rect 16037 19193 16071 19227
rect 30205 19193 30239 19227
rect 47961 19193 47995 19227
rect 5825 19125 5859 19159
rect 12725 19125 12759 19159
rect 15025 19125 15059 19159
rect 20453 19125 20487 19159
rect 23489 19125 23523 19159
rect 25789 19125 25823 19159
rect 27261 19125 27295 19159
rect 36645 19125 36679 19159
rect 36921 19125 36955 19159
rect 37933 19125 37967 19159
rect 41153 19125 41187 19159
rect 46673 19125 46707 19159
rect 9229 18921 9263 18955
rect 12541 18921 12575 18955
rect 13645 18921 13679 18955
rect 13829 18921 13863 18955
rect 16037 18921 16071 18955
rect 18153 18921 18187 18955
rect 19901 18921 19935 18955
rect 22293 18921 22327 18955
rect 28089 18921 28123 18955
rect 30941 18921 30975 18955
rect 33793 18921 33827 18955
rect 37381 18921 37415 18955
rect 42073 18921 42107 18955
rect 46857 18921 46891 18955
rect 11897 18853 11931 18887
rect 16957 18853 16991 18887
rect 21097 18853 21131 18887
rect 31493 18853 31527 18887
rect 48053 18853 48087 18887
rect 4169 18785 4203 18819
rect 10977 18785 11011 18819
rect 13093 18785 13127 18819
rect 14289 18785 14323 18819
rect 17509 18785 17543 18819
rect 18797 18785 18831 18819
rect 20361 18785 20395 18819
rect 20453 18785 20487 18819
rect 21649 18785 21683 18819
rect 25237 18785 25271 18819
rect 25789 18785 25823 18819
rect 27537 18785 27571 18819
rect 29929 18785 29963 18819
rect 31953 18785 31987 18819
rect 32137 18785 32171 18819
rect 32873 18785 32907 18819
rect 32965 18785 32999 18819
rect 34161 18785 34195 18819
rect 35633 18785 35667 18819
rect 38577 18785 38611 18819
rect 41797 18785 41831 18819
rect 2973 18717 3007 18751
rect 5365 18717 5399 18751
rect 8309 18717 8343 18751
rect 12081 18717 12115 18751
rect 18521 18717 18555 18751
rect 18613 18717 18647 18751
rect 24041 18717 24075 18751
rect 27813 18717 27847 18751
rect 28181 18717 28215 18751
rect 29193 18717 29227 18751
rect 34253 18717 34287 18751
rect 34437 18717 34471 18751
rect 35173 18717 35207 18751
rect 38393 18717 38427 18751
rect 47501 18717 47535 18751
rect 48237 18717 48271 18751
rect 48697 18717 48731 18751
rect 49341 18717 49375 18751
rect 1777 18649 1811 18683
rect 8125 18649 8159 18683
rect 10701 18649 10735 18683
rect 12909 18649 12943 18683
rect 13001 18649 13035 18683
rect 14565 18649 14599 18683
rect 16681 18649 16715 18683
rect 19441 18649 19475 18683
rect 20269 18649 20303 18683
rect 23765 18649 23799 18683
rect 26065 18649 26099 18683
rect 30113 18649 30147 18683
rect 30757 18649 30791 18683
rect 35909 18649 35943 18683
rect 39589 18649 39623 18683
rect 41521 18649 41555 18683
rect 47041 18649 47075 18683
rect 11345 18581 11379 18615
rect 11621 18581 11655 18615
rect 16405 18581 16439 18615
rect 17325 18581 17359 18615
rect 17417 18581 17451 18615
rect 19533 18581 19567 18615
rect 21465 18581 21499 18615
rect 21557 18581 21591 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 25053 18581 25087 18615
rect 28365 18581 28399 18615
rect 28641 18581 28675 18615
rect 29009 18581 29043 18615
rect 30021 18581 30055 18615
rect 30481 18581 30515 18615
rect 31125 18581 31159 18615
rect 31861 18581 31895 18615
rect 33057 18581 33091 18615
rect 33425 18581 33459 18615
rect 33885 18581 33919 18615
rect 37657 18581 37691 18615
rect 38025 18581 38059 18615
rect 38485 18581 38519 18615
rect 40049 18581 40083 18615
rect 47317 18581 47351 18615
rect 3617 18377 3651 18411
rect 9781 18377 9815 18411
rect 10793 18377 10827 18411
rect 17969 18377 18003 18411
rect 18429 18377 18463 18411
rect 22109 18377 22143 18411
rect 22477 18377 22511 18411
rect 26249 18377 26283 18411
rect 27629 18377 27663 18411
rect 28733 18377 28767 18411
rect 30849 18377 30883 18411
rect 32597 18377 32631 18411
rect 35357 18377 35391 18411
rect 35909 18377 35943 18411
rect 40417 18377 40451 18411
rect 40877 18377 40911 18411
rect 47685 18377 47719 18411
rect 7665 18309 7699 18343
rect 13185 18309 13219 18343
rect 14289 18309 14323 18343
rect 14381 18309 14415 18343
rect 16957 18309 16991 18343
rect 19901 18309 19935 18343
rect 24133 18309 24167 18343
rect 28825 18309 28859 18343
rect 40785 18309 40819 18343
rect 2973 18241 3007 18275
rect 3433 18241 3467 18275
rect 4445 18241 4479 18275
rect 7849 18241 7883 18275
rect 9965 18241 9999 18275
rect 10885 18241 10919 18275
rect 13461 18241 13495 18275
rect 16313 18241 16347 18275
rect 17233 18241 17267 18275
rect 17417 18241 17451 18275
rect 18337 18241 18371 18275
rect 22569 18241 22603 18275
rect 23305 18241 23339 18275
rect 25053 18241 25087 18275
rect 25145 18241 25179 18275
rect 26341 18241 26375 18275
rect 27537 18241 27571 18275
rect 30389 18241 30423 18275
rect 30481 18241 30515 18275
rect 31309 18241 31343 18275
rect 32689 18241 32723 18275
rect 36277 18241 36311 18275
rect 36369 18241 36403 18275
rect 37473 18241 37507 18275
rect 39773 18241 39807 18275
rect 48237 18241 48271 18275
rect 48697 18241 48731 18275
rect 49341 18241 49375 18275
rect 1777 18173 1811 18207
rect 4169 18173 4203 18207
rect 10977 18173 11011 18207
rect 14565 18173 14599 18207
rect 14933 18173 14967 18207
rect 15669 18173 15703 18207
rect 16773 18173 16807 18207
rect 18613 18173 18647 18207
rect 19349 18173 19383 18207
rect 19625 18173 19659 18207
rect 22661 18173 22695 18207
rect 25329 18173 25363 18207
rect 26433 18173 26467 18207
rect 27721 18173 27755 18207
rect 28917 18173 28951 18207
rect 30297 18173 30331 18207
rect 32505 18173 32539 18207
rect 33609 18173 33643 18207
rect 33885 18173 33919 18207
rect 36553 18173 36587 18207
rect 39497 18173 39531 18207
rect 40969 18173 41003 18207
rect 47409 18173 47443 18207
rect 13921 18105 13955 18139
rect 16129 18105 16163 18139
rect 24685 18105 24719 18139
rect 28365 18105 28399 18139
rect 37013 18105 37047 18139
rect 37381 18105 37415 18139
rect 38025 18105 38059 18139
rect 10425 18037 10459 18071
rect 11713 18037 11747 18071
rect 15209 18037 15243 18071
rect 18981 18037 19015 18071
rect 21373 18037 21407 18071
rect 25881 18037 25915 18071
rect 27169 18037 27203 18071
rect 29745 18037 29779 18071
rect 33057 18037 33091 18071
rect 37657 18037 37691 18071
rect 40049 18037 40083 18071
rect 48053 18037 48087 18071
rect 10149 17833 10183 17867
rect 10609 17833 10643 17867
rect 12909 17833 12943 17867
rect 14289 17833 14323 17867
rect 17509 17833 17543 17867
rect 19441 17833 19475 17867
rect 23305 17833 23339 17867
rect 25789 17833 25823 17867
rect 29561 17833 29595 17867
rect 34437 17833 34471 17867
rect 37307 17833 37341 17867
rect 40509 17833 40543 17867
rect 24593 17765 24627 17799
rect 33977 17765 34011 17799
rect 48053 17765 48087 17799
rect 12357 17697 12391 17731
rect 16037 17697 16071 17731
rect 16957 17697 16991 17731
rect 18797 17697 18831 17731
rect 21741 17697 21775 17731
rect 22017 17697 22051 17731
rect 23765 17697 23799 17731
rect 23949 17697 23983 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 31493 17697 31527 17731
rect 32965 17697 32999 17731
rect 33057 17697 33091 17731
rect 33885 17697 33919 17731
rect 38117 17697 38151 17731
rect 40969 17697 41003 17731
rect 41061 17697 41095 17731
rect 2973 17629 3007 17663
rect 13093 17629 13127 17663
rect 13737 17629 13771 17663
rect 17141 17629 17175 17663
rect 19625 17629 19659 17663
rect 22293 17629 22327 17663
rect 25973 17629 26007 17663
rect 26249 17629 26283 17663
rect 28825 17629 28859 17663
rect 30665 17629 30699 17663
rect 31585 17629 31619 17663
rect 37565 17629 37599 17663
rect 48237 17629 48271 17663
rect 48697 17629 48731 17663
rect 49341 17629 49375 17663
rect 1777 17561 1811 17595
rect 12081 17561 12115 17595
rect 15761 17561 15795 17595
rect 17049 17561 17083 17595
rect 17969 17561 18003 17595
rect 22845 17561 22879 17595
rect 23673 17561 23707 17595
rect 28549 17561 28583 17595
rect 29377 17561 29411 17595
rect 29929 17561 29963 17595
rect 31677 17561 31711 17595
rect 40877 17561 40911 17595
rect 47501 17561 47535 17595
rect 10333 17493 10367 17527
rect 13553 17493 13587 17527
rect 16497 17493 16531 17527
rect 20269 17493 20303 17527
rect 24961 17493 24995 17527
rect 26433 17493 26467 17527
rect 27077 17493 27111 17527
rect 29101 17493 29135 17527
rect 32045 17493 32079 17527
rect 32321 17493 32355 17527
rect 33149 17493 33183 17527
rect 33517 17493 33551 17527
rect 34345 17493 34379 17527
rect 35081 17493 35115 17527
rect 35449 17493 35483 17527
rect 35817 17493 35851 17527
rect 38301 17493 38335 17527
rect 38393 17493 38427 17527
rect 38761 17493 38795 17527
rect 39037 17493 39071 17527
rect 39221 17493 39255 17527
rect 47685 17493 47719 17527
rect 11805 17289 11839 17323
rect 14197 17289 14231 17323
rect 17417 17289 17451 17323
rect 19165 17289 19199 17323
rect 22661 17289 22695 17323
rect 24869 17289 24903 17323
rect 25329 17289 25363 17323
rect 27353 17289 27387 17323
rect 29009 17289 29043 17323
rect 37841 17289 37875 17323
rect 38485 17289 38519 17323
rect 40969 17289 41003 17323
rect 47041 17289 47075 17323
rect 11897 17221 11931 17255
rect 13001 17221 13035 17255
rect 13093 17221 13127 17255
rect 14289 17221 14323 17255
rect 17969 17221 18003 17255
rect 20637 17221 20671 17255
rect 21925 17221 21959 17255
rect 25973 17221 26007 17255
rect 28917 17221 28951 17255
rect 30205 17221 30239 17255
rect 35541 17221 35575 17255
rect 37013 17221 37047 17255
rect 40417 17221 40451 17255
rect 2973 17153 3007 17187
rect 9873 17153 9907 17187
rect 10793 17153 10827 17187
rect 15117 17153 15151 17187
rect 15945 17153 15979 17187
rect 17049 17153 17083 17187
rect 18705 17153 18739 17187
rect 20913 17153 20947 17187
rect 24409 17153 24443 17187
rect 25237 17153 25271 17187
rect 27721 17153 27755 17187
rect 31309 17153 31343 17187
rect 31401 17153 31435 17187
rect 32321 17153 32355 17187
rect 36277 17153 36311 17187
rect 36369 17153 36403 17187
rect 37933 17153 37967 17187
rect 47225 17153 47259 17187
rect 48145 17153 48179 17187
rect 48697 17153 48731 17187
rect 49341 17153 49375 17187
rect 1777 17085 1811 17119
rect 9505 17085 9539 17119
rect 10517 17085 10551 17119
rect 10701 17085 10735 17119
rect 12817 17085 12851 17119
rect 16037 17085 16071 17119
rect 16129 17085 16163 17119
rect 24133 17085 24167 17119
rect 25513 17085 25547 17119
rect 27813 17085 27847 17119
rect 27905 17085 27939 17119
rect 28733 17085 28767 17119
rect 30021 17085 30055 17119
rect 30113 17085 30147 17119
rect 31125 17085 31159 17119
rect 32597 17085 32631 17119
rect 34069 17085 34103 17119
rect 34805 17085 34839 17119
rect 36093 17085 36127 17119
rect 38025 17085 38059 17119
rect 40693 17085 40727 17119
rect 47961 17085 47995 17119
rect 9781 17017 9815 17051
rect 10057 17017 10091 17051
rect 11161 17017 11195 17051
rect 12449 17017 12483 17051
rect 14933 17017 14967 17051
rect 15577 17017 15611 17051
rect 21281 17017 21315 17051
rect 21649 17017 21683 17051
rect 29377 17017 29411 17051
rect 30573 17017 30607 17051
rect 13461 16949 13495 16983
rect 13737 16949 13771 16983
rect 16957 16949 16991 16983
rect 31769 16949 31803 16983
rect 36737 16949 36771 16983
rect 37473 16949 37507 16983
rect 38945 16949 38979 16983
rect 47685 16949 47719 16983
rect 10425 16745 10459 16779
rect 16681 16745 16715 16779
rect 24685 16745 24719 16779
rect 28273 16745 28307 16779
rect 29377 16745 29411 16779
rect 34529 16745 34563 16779
rect 36277 16745 36311 16779
rect 41061 16745 41095 16779
rect 41245 16745 41279 16779
rect 21005 16677 21039 16711
rect 28825 16677 28859 16711
rect 29193 16677 29227 16711
rect 41521 16677 41555 16711
rect 7941 16609 7975 16643
rect 11161 16609 11195 16643
rect 13185 16609 13219 16643
rect 13277 16609 13311 16643
rect 14197 16609 14231 16643
rect 14657 16609 14691 16643
rect 16129 16609 16163 16643
rect 16221 16609 16255 16643
rect 18613 16609 18647 16643
rect 18889 16609 18923 16643
rect 22477 16609 22511 16643
rect 22753 16609 22787 16643
rect 23765 16609 23799 16643
rect 23949 16609 23983 16643
rect 25605 16609 25639 16643
rect 27077 16609 27111 16643
rect 27629 16609 27663 16643
rect 29837 16609 29871 16643
rect 30021 16609 30055 16643
rect 31125 16609 31159 16643
rect 31217 16609 31251 16643
rect 32229 16609 32263 16643
rect 32505 16609 32539 16643
rect 35081 16609 35115 16643
rect 36921 16609 36955 16643
rect 39221 16609 39255 16643
rect 40233 16609 40267 16643
rect 47685 16609 47719 16643
rect 2973 16541 3007 16575
rect 8125 16541 8159 16575
rect 12357 16541 12391 16575
rect 13369 16541 13403 16575
rect 14841 16541 14875 16575
rect 20269 16541 20303 16575
rect 24593 16541 24627 16575
rect 27353 16541 27387 16575
rect 30113 16541 30147 16575
rect 35817 16541 35851 16575
rect 36737 16541 36771 16575
rect 37289 16541 37323 16575
rect 39497 16541 39531 16575
rect 48237 16541 48271 16575
rect 48697 16541 48731 16575
rect 49341 16541 49375 16575
rect 1777 16473 1811 16507
rect 8033 16473 8067 16507
rect 10057 16473 10091 16507
rect 10517 16473 10551 16507
rect 11437 16473 11471 16507
rect 28457 16473 28491 16507
rect 40325 16473 40359 16507
rect 40417 16473 40451 16507
rect 8493 16405 8527 16439
rect 9045 16405 9079 16439
rect 11345 16405 11379 16439
rect 11805 16405 11839 16439
rect 12541 16405 12575 16439
rect 13737 16405 13771 16439
rect 14749 16405 14783 16439
rect 15209 16405 15243 16439
rect 15669 16405 15703 16439
rect 16037 16405 16071 16439
rect 17141 16405 17175 16439
rect 19441 16405 19475 16439
rect 20085 16405 20119 16439
rect 20637 16405 20671 16439
rect 23305 16405 23339 16439
rect 23673 16405 23707 16439
rect 27997 16405 28031 16439
rect 28549 16405 28583 16439
rect 30481 16405 30515 16439
rect 31309 16405 31343 16439
rect 31677 16405 31711 16439
rect 33977 16405 34011 16439
rect 34345 16405 34379 16439
rect 36645 16405 36679 16439
rect 37749 16405 37783 16439
rect 40785 16405 40819 16439
rect 48053 16405 48087 16439
rect 8309 16201 8343 16235
rect 9229 16201 9263 16235
rect 10977 16201 11011 16235
rect 11989 16201 12023 16235
rect 12449 16201 12483 16235
rect 13185 16201 13219 16235
rect 14749 16201 14783 16235
rect 17417 16201 17451 16235
rect 17785 16201 17819 16235
rect 30941 16201 30975 16235
rect 33793 16201 33827 16235
rect 40509 16201 40543 16235
rect 40969 16201 41003 16235
rect 13553 16133 13587 16167
rect 19441 16133 19475 16167
rect 30849 16133 30883 16167
rect 32597 16133 32631 16167
rect 34529 16133 34563 16167
rect 38485 16133 38519 16167
rect 2973 16065 3007 16099
rect 8217 16065 8251 16099
rect 9321 16065 9355 16099
rect 10425 16065 10459 16099
rect 11069 16065 11103 16099
rect 12357 16065 12391 16099
rect 15853 16065 15887 16099
rect 15945 16065 15979 16099
rect 17049 16065 17083 16099
rect 19165 16065 19199 16099
rect 23489 16065 23523 16099
rect 26341 16065 26375 16099
rect 27537 16065 27571 16099
rect 27629 16065 27663 16099
rect 28365 16065 28399 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 36921 16065 36955 16099
rect 38209 16065 38243 16099
rect 40877 16065 40911 16099
rect 48421 16065 48455 16099
rect 48697 16065 48731 16099
rect 1777 15997 1811 16031
rect 8125 15997 8159 16031
rect 12633 15997 12667 16031
rect 13645 15997 13679 16031
rect 13737 15997 13771 16031
rect 14841 15997 14875 16031
rect 14933 15997 14967 16031
rect 15761 15997 15795 16031
rect 16957 15997 16991 16031
rect 17877 15997 17911 16031
rect 17969 15997 18003 16031
rect 20913 15997 20947 16031
rect 23305 15997 23339 16031
rect 23397 15997 23431 16031
rect 24593 15997 24627 16031
rect 26065 15997 26099 16031
rect 27721 15997 27755 16031
rect 28641 15997 28675 16031
rect 30665 15997 30699 16031
rect 31861 15997 31895 16031
rect 32413 15997 32447 16031
rect 33609 15997 33643 16031
rect 36645 15997 36679 16031
rect 37473 15997 37507 16031
rect 41061 15997 41095 16031
rect 8677 15929 8711 15963
rect 14381 15929 14415 15963
rect 16313 15929 16347 15963
rect 18889 15929 18923 15963
rect 23857 15929 23891 15963
rect 26709 15929 26743 15963
rect 34253 15929 34287 15963
rect 10517 15861 10551 15895
rect 11621 15861 11655 15895
rect 16773 15861 16807 15895
rect 21281 15861 21315 15895
rect 21557 15861 21591 15895
rect 22753 15861 22787 15895
rect 27169 15861 27203 15895
rect 30113 15861 30147 15895
rect 31309 15861 31343 15895
rect 31677 15861 31711 15895
rect 33057 15861 33091 15895
rect 34713 15861 34747 15895
rect 35173 15861 35207 15895
rect 39957 15861 39991 15895
rect 41613 15861 41647 15895
rect 49341 15861 49375 15895
rect 10793 15657 10827 15691
rect 16773 15657 16807 15691
rect 17877 15657 17911 15691
rect 18061 15657 18095 15691
rect 18981 15657 19015 15691
rect 19349 15657 19383 15691
rect 19901 15657 19935 15691
rect 21189 15657 21223 15691
rect 26985 15657 27019 15691
rect 28549 15657 28583 15691
rect 29285 15657 29319 15691
rect 34437 15657 34471 15691
rect 36645 15657 36679 15691
rect 37749 15657 37783 15691
rect 42073 15657 42107 15691
rect 48421 15657 48455 15691
rect 49157 15657 49191 15691
rect 18429 15589 18463 15623
rect 22293 15589 22327 15623
rect 32229 15589 32263 15623
rect 41797 15589 41831 15623
rect 10517 15521 10551 15555
rect 12265 15521 12299 15555
rect 12541 15521 12575 15555
rect 13185 15521 13219 15555
rect 14841 15521 14875 15555
rect 16129 15521 16163 15555
rect 17325 15521 17359 15555
rect 20545 15521 20579 15555
rect 21741 15521 21775 15555
rect 23673 15521 23707 15555
rect 25237 15521 25271 15555
rect 26433 15521 26467 15555
rect 27997 15521 28031 15555
rect 30481 15521 30515 15555
rect 32873 15521 32907 15555
rect 32965 15521 32999 15555
rect 34897 15521 34931 15555
rect 35173 15521 35207 15555
rect 39497 15521 39531 15555
rect 40049 15521 40083 15555
rect 40325 15521 40359 15555
rect 2973 15453 3007 15487
rect 15945 15453 15979 15487
rect 18613 15453 18647 15487
rect 21649 15453 21683 15487
rect 23581 15453 23615 15487
rect 27905 15453 27939 15487
rect 28641 15453 28675 15487
rect 29193 15453 29227 15487
rect 48145 15453 48179 15487
rect 48605 15453 48639 15487
rect 49341 15453 49375 15487
rect 1777 15385 1811 15419
rect 6377 15385 6411 15419
rect 6561 15385 6595 15419
rect 13277 15385 13311 15419
rect 13369 15385 13403 15419
rect 14749 15385 14783 15419
rect 20361 15385 20395 15419
rect 23489 15385 23523 15419
rect 25053 15385 25087 15419
rect 26249 15385 26283 15419
rect 26341 15385 26375 15419
rect 27813 15385 27847 15419
rect 29009 15385 29043 15419
rect 30757 15385 30791 15419
rect 39221 15385 39255 15419
rect 9045 15317 9079 15351
rect 13737 15317 13771 15351
rect 14289 15317 14323 15351
rect 14657 15317 14691 15351
rect 15577 15317 15611 15351
rect 16037 15317 16071 15351
rect 17141 15317 17175 15351
rect 17233 15317 17267 15351
rect 19533 15317 19567 15351
rect 20269 15317 20303 15351
rect 21557 15317 21591 15351
rect 23121 15317 23155 15351
rect 24133 15317 24167 15351
rect 24685 15317 24719 15351
rect 25145 15317 25179 15351
rect 25881 15317 25915 15351
rect 27077 15317 27111 15351
rect 27445 15317 27479 15351
rect 30021 15317 30055 15351
rect 33057 15317 33091 15351
rect 33425 15317 33459 15351
rect 33885 15317 33919 15351
rect 37105 15317 37139 15351
rect 9689 15113 9723 15147
rect 9781 15113 9815 15147
rect 11897 15113 11931 15147
rect 13001 15113 13035 15147
rect 13369 15113 13403 15147
rect 15577 15113 15611 15147
rect 15945 15113 15979 15147
rect 18337 15113 18371 15147
rect 18797 15113 18831 15147
rect 19533 15113 19567 15147
rect 22937 15113 22971 15147
rect 24133 15113 24167 15147
rect 25329 15113 25363 15147
rect 25605 15113 25639 15147
rect 26341 15113 26375 15147
rect 27445 15113 27479 15147
rect 29745 15113 29779 15147
rect 30573 15113 30607 15147
rect 31401 15113 31435 15147
rect 33885 15113 33919 15147
rect 35081 15113 35115 15147
rect 39681 15113 39715 15147
rect 40141 15113 40175 15147
rect 10885 15045 10919 15079
rect 11069 15045 11103 15079
rect 16037 15045 16071 15079
rect 19901 15045 19935 15079
rect 21097 15045 21131 15079
rect 21833 15045 21867 15079
rect 23397 15045 23431 15079
rect 27077 15045 27111 15079
rect 31861 15045 31895 15079
rect 36185 15045 36219 15079
rect 36277 15045 36311 15079
rect 37749 15045 37783 15079
rect 1777 14977 1811 15011
rect 2973 14977 3007 15011
rect 12265 14977 12299 15011
rect 12357 14977 12391 15011
rect 15117 14977 15151 15011
rect 17233 14977 17267 15011
rect 18705 14977 18739 15011
rect 19993 14977 20027 15011
rect 22017 14977 22051 15011
rect 23305 14977 23339 15011
rect 24501 14977 24535 15011
rect 24593 14977 24627 15011
rect 25237 14977 25271 15011
rect 26249 14977 26283 15011
rect 27261 14977 27295 15011
rect 27997 14977 28031 15011
rect 30665 14977 30699 15011
rect 32689 14977 32723 15011
rect 32781 14977 32815 15011
rect 37473 14977 37507 15011
rect 40049 14977 40083 15011
rect 40877 14977 40911 15011
rect 48237 14977 48271 15011
rect 48697 14977 48731 15011
rect 49341 14977 49375 15011
rect 9597 14909 9631 14943
rect 11621 14909 11655 14943
rect 12449 14909 12483 14943
rect 14841 14909 14875 14943
rect 16129 14909 16163 14943
rect 17325 14909 17359 14943
rect 17417 14909 17451 14943
rect 18889 14909 18923 14943
rect 20177 14909 20211 14943
rect 21189 14909 21223 14943
rect 21373 14909 21407 14943
rect 23581 14909 23615 14943
rect 24685 14909 24719 14943
rect 26433 14909 26467 14943
rect 28273 14909 28307 14943
rect 30757 14909 30791 14943
rect 32873 14909 32907 14943
rect 33701 14909 33735 14943
rect 33793 14909 33827 14943
rect 34897 14909 34931 14943
rect 34989 14909 35023 14943
rect 36093 14909 36127 14943
rect 39221 14909 39255 14943
rect 40233 14909 40267 14943
rect 47685 14909 47719 14943
rect 10149 14841 10183 14875
rect 18061 14841 18095 14875
rect 20729 14841 20763 14875
rect 32321 14841 32355 14875
rect 36645 14841 36679 14875
rect 48053 14841 48087 14875
rect 10609 14773 10643 14807
rect 16865 14773 16899 14807
rect 25881 14773 25915 14807
rect 27537 14773 27571 14807
rect 30205 14773 30239 14807
rect 34253 14773 34287 14807
rect 35449 14773 35483 14807
rect 36921 14773 36955 14807
rect 41061 14773 41095 14807
rect 11805 14569 11839 14603
rect 13001 14569 13035 14603
rect 14473 14569 14507 14603
rect 18153 14569 18187 14603
rect 22845 14569 22879 14603
rect 25605 14569 25639 14603
rect 36645 14569 36679 14603
rect 38589 14569 38623 14603
rect 39865 14569 39899 14603
rect 40049 14569 40083 14603
rect 10241 14501 10275 14535
rect 20729 14501 20763 14535
rect 30481 14501 30515 14535
rect 34069 14501 34103 14535
rect 1777 14433 1811 14467
rect 12449 14433 12483 14467
rect 13553 14433 13587 14467
rect 14197 14433 14231 14467
rect 15117 14433 15151 14467
rect 16957 14433 16991 14467
rect 17509 14433 17543 14467
rect 18705 14433 18739 14467
rect 20085 14433 20119 14467
rect 21097 14433 21131 14467
rect 21373 14433 21407 14467
rect 27077 14433 27111 14467
rect 27905 14433 27939 14467
rect 29929 14433 29963 14467
rect 31033 14433 31067 14467
rect 32229 14433 32263 14467
rect 33425 14433 33459 14467
rect 34897 14433 34931 14467
rect 38853 14433 38887 14467
rect 47685 14433 47719 14467
rect 2973 14365 3007 14399
rect 9505 14365 9539 14399
rect 11253 14365 11287 14399
rect 14841 14365 14875 14399
rect 17601 14365 17635 14399
rect 18521 14365 18555 14399
rect 19901 14365 19935 14399
rect 23489 14365 23523 14399
rect 24685 14365 24719 14399
rect 27353 14365 27387 14399
rect 28089 14365 28123 14399
rect 31309 14365 31343 14399
rect 32413 14365 32447 14399
rect 33609 14365 33643 14399
rect 33701 14365 33735 14399
rect 39313 14365 39347 14399
rect 47961 14365 47995 14399
rect 49341 14365 49375 14399
rect 9689 14297 9723 14331
rect 10425 14297 10459 14331
rect 12173 14297 12207 14331
rect 13369 14297 13403 14331
rect 15945 14297 15979 14331
rect 16773 14297 16807 14331
rect 20545 14297 20579 14331
rect 28181 14297 28215 14331
rect 31217 14297 31251 14331
rect 35173 14297 35207 14331
rect 48145 14297 48179 14331
rect 48697 14297 48731 14331
rect 11161 14229 11195 14263
rect 12265 14229 12299 14263
rect 13461 14229 13495 14263
rect 14933 14229 14967 14263
rect 16405 14229 16439 14263
rect 16865 14229 16899 14263
rect 17877 14229 17911 14263
rect 18613 14229 18647 14263
rect 19533 14229 19567 14263
rect 19993 14229 20027 14263
rect 23213 14229 23247 14263
rect 23857 14229 23891 14263
rect 24409 14229 24443 14263
rect 25145 14229 25179 14263
rect 28549 14229 28583 14263
rect 29009 14229 29043 14263
rect 30021 14229 30055 14263
rect 30113 14229 30147 14263
rect 31677 14229 31711 14263
rect 32505 14229 32539 14263
rect 32873 14229 32907 14263
rect 34345 14229 34379 14263
rect 37105 14229 37139 14263
rect 39497 14229 39531 14263
rect 3617 14025 3651 14059
rect 9965 14025 9999 14059
rect 10701 14025 10735 14059
rect 11989 14025 12023 14059
rect 15577 14025 15611 14059
rect 16773 14025 16807 14059
rect 17141 14025 17175 14059
rect 17509 14025 17543 14059
rect 17601 14025 17635 14059
rect 18337 14025 18371 14059
rect 18705 14025 18739 14059
rect 21465 14025 21499 14059
rect 22017 14025 22051 14059
rect 24869 14025 24903 14059
rect 27629 14025 27663 14059
rect 29377 14025 29411 14059
rect 31769 14025 31803 14059
rect 36093 14025 36127 14059
rect 36461 14025 36495 14059
rect 37841 14025 37875 14059
rect 38209 14025 38243 14059
rect 45845 14025 45879 14059
rect 1777 13957 1811 13991
rect 13277 13957 13311 13991
rect 15025 13957 15059 13991
rect 16037 13957 16071 13991
rect 26341 13957 26375 13991
rect 34805 13957 34839 13991
rect 34897 13957 34931 13991
rect 36921 13957 36955 13991
rect 37749 13957 37783 13991
rect 38577 13957 38611 13991
rect 38945 13957 38979 13991
rect 45017 13957 45051 13991
rect 47961 13957 47995 13991
rect 2973 13889 3007 13923
rect 3525 13889 3559 13923
rect 3985 13889 4019 13923
rect 11161 13889 11195 13923
rect 12081 13889 12115 13923
rect 15209 13889 15243 13923
rect 15945 13889 15979 13923
rect 19441 13889 19475 13923
rect 23765 13889 23799 13923
rect 28917 13889 28951 13923
rect 31125 13889 31159 13923
rect 36001 13889 36035 13923
rect 45661 13889 45695 13923
rect 47225 13889 47259 13923
rect 48145 13889 48179 13923
rect 48697 13889 48731 13923
rect 49341 13889 49375 13923
rect 10517 13821 10551 13855
rect 11897 13821 11931 13855
rect 13001 13821 13035 13855
rect 16129 13821 16163 13855
rect 17785 13821 17819 13855
rect 18797 13821 18831 13855
rect 18889 13821 18923 13855
rect 19717 13821 19751 13855
rect 23489 13821 23523 13855
rect 24225 13821 24259 13855
rect 26617 13821 26651 13855
rect 30849 13821 30883 13855
rect 32321 13821 32355 13855
rect 34069 13821 34103 13855
rect 34621 13821 34655 13855
rect 35909 13821 35943 13855
rect 37657 13821 37691 13855
rect 45201 13821 45235 13855
rect 47685 13821 47719 13855
rect 35265 13753 35299 13787
rect 36737 13753 36771 13787
rect 47041 13753 47075 13787
rect 12449 13685 12483 13719
rect 14749 13685 14783 13719
rect 19980 13685 20014 13719
rect 33811 13685 33845 13719
rect 13645 13481 13679 13515
rect 13921 13481 13955 13515
rect 18153 13481 18187 13515
rect 19441 13481 19475 13515
rect 20453 13481 20487 13515
rect 20913 13481 20947 13515
rect 24041 13481 24075 13515
rect 25605 13481 25639 13515
rect 28181 13481 28215 13515
rect 29193 13481 29227 13515
rect 35633 13481 35667 13515
rect 38209 13481 38243 13515
rect 38577 13481 38611 13515
rect 39589 13481 39623 13515
rect 47685 13481 47719 13515
rect 14289 13413 14323 13447
rect 22109 13413 22143 13447
rect 33333 13413 33367 13447
rect 36185 13413 36219 13447
rect 1777 13345 1811 13379
rect 10793 13345 10827 13379
rect 12541 13345 12575 13379
rect 13093 13345 13127 13379
rect 15393 13345 15427 13379
rect 15485 13345 15519 13379
rect 16405 13345 16439 13379
rect 19901 13345 19935 13379
rect 21373 13345 21407 13379
rect 21557 13345 21591 13379
rect 22569 13345 22603 13379
rect 22753 13345 22787 13379
rect 23489 13345 23523 13379
rect 25053 13345 25087 13379
rect 28549 13345 28583 13379
rect 29837 13345 29871 13379
rect 30021 13345 30055 13379
rect 31125 13345 31159 13379
rect 33885 13345 33919 13379
rect 34345 13345 34379 13379
rect 35081 13345 35115 13379
rect 2973 13277 3007 13311
rect 14473 13277 14507 13311
rect 15577 13277 15611 13311
rect 22477 13277 22511 13311
rect 23673 13277 23707 13311
rect 25237 13277 25271 13311
rect 28825 13277 28859 13311
rect 30113 13277 30147 13311
rect 32873 13277 32907 13311
rect 36461 13277 36495 13311
rect 41337 13277 41371 13311
rect 47961 13277 47995 13311
rect 49157 13277 49191 13311
rect 10517 13209 10551 13243
rect 11069 13209 11103 13243
rect 14841 13209 14875 13243
rect 16681 13209 16715 13243
rect 18889 13209 18923 13243
rect 20085 13209 20119 13243
rect 26801 13209 26835 13243
rect 27537 13209 27571 13243
rect 32597 13209 32631 13243
rect 35265 13209 35299 13243
rect 36737 13209 36771 13243
rect 15945 13141 15979 13175
rect 19993 13141 20027 13175
rect 21281 13141 21315 13175
rect 23581 13141 23615 13175
rect 24501 13141 24535 13175
rect 25145 13141 25179 13175
rect 26065 13141 26099 13175
rect 27721 13141 27755 13175
rect 27905 13141 27939 13175
rect 28733 13141 28767 13175
rect 30481 13141 30515 13175
rect 33701 13141 33735 13175
rect 33793 13141 33827 13175
rect 35173 13141 35207 13175
rect 36001 13141 36035 13175
rect 41521 13141 41555 13175
rect 1777 12937 1811 12971
rect 11345 12937 11379 12971
rect 11989 12937 12023 12971
rect 12817 12937 12851 12971
rect 13093 12937 13127 12971
rect 15853 12937 15887 12971
rect 20729 12937 20763 12971
rect 21189 12937 21223 12971
rect 23397 12937 23431 12971
rect 26709 12937 26743 12971
rect 32597 12937 32631 12971
rect 35817 12937 35851 12971
rect 36645 12937 36679 12971
rect 1685 12869 1719 12903
rect 2145 12869 2179 12903
rect 11161 12869 11195 12903
rect 14565 12869 14599 12903
rect 15945 12869 15979 12903
rect 16681 12869 16715 12903
rect 18705 12869 18739 12903
rect 25329 12869 25363 12903
rect 26157 12869 26191 12903
rect 27169 12869 27203 12903
rect 28917 12869 28951 12903
rect 29561 12869 29595 12903
rect 33425 12869 33459 12903
rect 34805 12869 34839 12903
rect 37013 12869 37047 12903
rect 2881 12801 2915 12835
rect 12081 12801 12115 12835
rect 14841 12801 14875 12835
rect 16957 12801 16991 12835
rect 17877 12801 17911 12835
rect 19625 12801 19659 12835
rect 20361 12801 20395 12835
rect 21097 12801 21131 12835
rect 23029 12801 23063 12835
rect 25605 12801 25639 12835
rect 29193 12801 29227 12835
rect 30021 12801 30055 12835
rect 32689 12801 32723 12835
rect 34069 12801 34103 12835
rect 36829 12801 36863 12835
rect 37473 12801 37507 12835
rect 40049 12801 40083 12835
rect 40509 12801 40543 12835
rect 45937 12801 45971 12835
rect 47961 12801 47995 12835
rect 49157 12801 49191 12835
rect 11805 12733 11839 12767
rect 15669 12733 15703 12767
rect 17417 12733 17451 12767
rect 19717 12733 19751 12767
rect 19901 12733 19935 12767
rect 21281 12733 21315 12767
rect 22017 12733 22051 12767
rect 22753 12733 22787 12767
rect 22937 12733 22971 12767
rect 30297 12733 30331 12767
rect 32413 12733 32447 12767
rect 35541 12733 35575 12767
rect 35725 12733 35759 12767
rect 36461 12733 36495 12767
rect 37749 12733 37783 12767
rect 39497 12733 39531 12767
rect 2513 12665 2547 12699
rect 15301 12665 15335 12699
rect 19257 12665 19291 12699
rect 23857 12665 23891 12699
rect 33057 12665 33091 12699
rect 36185 12665 36219 12699
rect 40233 12665 40267 12699
rect 2329 12597 2363 12631
rect 3525 12597 3559 12631
rect 12449 12597 12483 12631
rect 16313 12597 16347 12631
rect 25973 12597 26007 12631
rect 31769 12597 31803 12631
rect 33517 12597 33551 12631
rect 33701 12597 33735 12631
rect 46121 12597 46155 12631
rect 3065 12393 3099 12427
rect 11253 12393 11287 12427
rect 14381 12393 14415 12427
rect 15865 12393 15899 12427
rect 19441 12393 19475 12427
rect 26341 12393 26375 12427
rect 27721 12393 27755 12427
rect 39313 12393 39347 12427
rect 39497 12393 39531 12427
rect 21649 12325 21683 12359
rect 26709 12325 26743 12359
rect 39037 12325 39071 12359
rect 40325 12325 40359 12359
rect 2145 12257 2179 12291
rect 9505 12257 9539 12291
rect 11713 12257 11747 12291
rect 16129 12257 16163 12291
rect 16497 12257 16531 12291
rect 17325 12257 17359 12291
rect 19993 12257 20027 12291
rect 20637 12257 20671 12291
rect 21005 12257 21039 12291
rect 22293 12257 22327 12291
rect 22385 12257 22419 12291
rect 23949 12257 23983 12291
rect 24869 12257 24903 12291
rect 27169 12257 27203 12291
rect 28365 12257 28399 12291
rect 29745 12257 29779 12291
rect 31769 12257 31803 12291
rect 33885 12257 33919 12291
rect 37197 12257 37231 12291
rect 38393 12257 38427 12291
rect 38577 12257 38611 12291
rect 49157 12257 49191 12291
rect 2421 12189 2455 12223
rect 2881 12189 2915 12223
rect 17141 12189 17175 12223
rect 19809 12189 19843 12223
rect 21281 12189 21315 12223
rect 24593 12189 24627 12223
rect 29193 12189 29227 12223
rect 32137 12189 32171 12223
rect 34345 12189 34379 12223
rect 34897 12189 34931 12223
rect 37381 12189 37415 12223
rect 40785 12189 40819 12223
rect 41429 12189 41463 12223
rect 45937 12189 45971 12223
rect 47961 12189 47995 12223
rect 9781 12121 9815 12155
rect 11989 12121 12023 12155
rect 13737 12121 13771 12155
rect 18153 12121 18187 12155
rect 18889 12121 18923 12155
rect 22477 12121 22511 12155
rect 23673 12121 23707 12155
rect 27261 12121 27295 12155
rect 30021 12121 30055 12155
rect 32413 12121 32447 12155
rect 35173 12121 35207 12155
rect 40141 12121 40175 12155
rect 16773 12053 16807 12087
rect 17233 12053 17267 12087
rect 19901 12053 19935 12087
rect 21189 12053 21223 12087
rect 22845 12053 22879 12087
rect 23305 12053 23339 12087
rect 23765 12053 23799 12087
rect 27353 12053 27387 12087
rect 31493 12053 31527 12087
rect 34161 12053 34195 12087
rect 36645 12053 36679 12087
rect 37473 12053 37507 12087
rect 37841 12053 37875 12087
rect 38669 12053 38703 12087
rect 40969 12053 41003 12087
rect 41613 12053 41647 12087
rect 46121 12053 46155 12087
rect 2237 11849 2271 11883
rect 3985 11849 4019 11883
rect 11621 11849 11655 11883
rect 12725 11849 12759 11883
rect 13553 11849 13587 11883
rect 14197 11849 14231 11883
rect 14289 11849 14323 11883
rect 16865 11849 16899 11883
rect 19901 11849 19935 11883
rect 20269 11849 20303 11883
rect 20729 11849 20763 11883
rect 21097 11849 21131 11883
rect 22109 11849 22143 11883
rect 25697 11849 25731 11883
rect 26617 11849 26651 11883
rect 27905 11849 27939 11883
rect 31493 11849 31527 11883
rect 32597 11849 32631 11883
rect 32689 11849 32723 11883
rect 33057 11849 33091 11883
rect 33885 11849 33919 11883
rect 34713 11849 34747 11883
rect 37749 11849 37783 11883
rect 38669 11849 38703 11883
rect 39129 11849 39163 11883
rect 12817 11781 12851 11815
rect 15577 11781 15611 11815
rect 18337 11781 18371 11815
rect 23397 11781 23431 11815
rect 26157 11781 26191 11815
rect 27537 11781 27571 11815
rect 30021 11781 30055 11815
rect 39957 11781 39991 11815
rect 40417 11781 40451 11815
rect 45109 11781 45143 11815
rect 49157 11781 49191 11815
rect 1593 11713 1627 11747
rect 2697 11713 2731 11747
rect 3341 11713 3375 11747
rect 3801 11713 3835 11747
rect 15485 11713 15519 11747
rect 16405 11713 16439 11747
rect 19809 11713 19843 11747
rect 22569 11713 22603 11747
rect 23949 11713 23983 11747
rect 31125 11713 31159 11747
rect 33793 11713 33827 11747
rect 37841 11713 37875 11747
rect 39037 11713 39071 11747
rect 40601 11713 40635 11747
rect 47961 11713 47995 11747
rect 12909 11645 12943 11679
rect 14105 11645 14139 11679
rect 15669 11645 15703 11679
rect 18613 11645 18647 11679
rect 19073 11645 19107 11679
rect 19717 11645 19751 11679
rect 21189 11645 21223 11679
rect 21373 11645 21407 11679
rect 24225 11645 24259 11679
rect 27353 11645 27387 11679
rect 27445 11645 27479 11679
rect 30297 11645 30331 11679
rect 30849 11645 30883 11679
rect 31033 11645 31067 11679
rect 32505 11645 32539 11679
rect 33609 11645 33643 11679
rect 35173 11645 35207 11679
rect 35449 11645 35483 11679
rect 37565 11645 37599 11679
rect 39221 11645 39255 11679
rect 14657 11577 14691 11611
rect 36921 11577 36955 11611
rect 40141 11577 40175 11611
rect 45293 11577 45327 11611
rect 11989 11509 12023 11543
rect 12357 11509 12391 11543
rect 13369 11509 13403 11543
rect 15117 11509 15151 11543
rect 16221 11509 16255 11543
rect 19165 11509 19199 11543
rect 21833 11509 21867 11543
rect 22293 11509 22327 11543
rect 28549 11509 28583 11543
rect 31769 11509 31803 11543
rect 34253 11509 34287 11543
rect 34529 11509 34563 11543
rect 38209 11509 38243 11543
rect 2881 11305 2915 11339
rect 13277 11305 13311 11339
rect 14381 11305 14415 11339
rect 16773 11305 16807 11339
rect 19073 11305 19107 11339
rect 19349 11305 19383 11339
rect 23305 11305 23339 11339
rect 26341 11305 26375 11339
rect 28641 11305 28675 11339
rect 29009 11305 29043 11339
rect 30481 11305 30515 11339
rect 34713 11305 34747 11339
rect 38761 11305 38795 11339
rect 39589 11305 39623 11339
rect 3249 11237 3283 11271
rect 4169 11237 4203 11271
rect 16313 11237 16347 11271
rect 19533 11237 19567 11271
rect 20453 11237 20487 11271
rect 32873 11237 32907 11271
rect 38393 11237 38427 11271
rect 40969 11237 41003 11271
rect 3433 11169 3467 11203
rect 10977 11169 11011 11203
rect 12449 11169 12483 11203
rect 13093 11169 13127 11203
rect 14841 11169 14875 11203
rect 15025 11169 15059 11203
rect 15761 11169 15795 11203
rect 15853 11169 15887 11203
rect 17417 11169 17451 11203
rect 18613 11169 18647 11203
rect 19993 11169 20027 11203
rect 23765 11169 23799 11203
rect 23949 11169 23983 11203
rect 24869 11169 24903 11203
rect 29929 11169 29963 11203
rect 34069 11169 34103 11203
rect 37749 11169 37783 11203
rect 49157 11169 49191 11203
rect 1593 11101 1627 11135
rect 2237 11101 2271 11135
rect 2697 11101 2731 11135
rect 3985 11101 4019 11135
rect 12725 11101 12759 11135
rect 15945 11101 15979 11135
rect 17141 11101 17175 11135
rect 22201 11101 22235 11135
rect 22661 11101 22695 11135
rect 24593 11101 24627 11135
rect 26893 11101 26927 11135
rect 30021 11101 30055 11135
rect 31125 11101 31159 11135
rect 33333 11101 33367 11135
rect 38209 11101 38243 11135
rect 40141 11101 40175 11135
rect 40785 11101 40819 11135
rect 45661 11101 45695 11135
rect 47961 11101 47995 11135
rect 13737 11033 13771 11067
rect 14749 11033 14783 11067
rect 18337 11033 18371 11067
rect 21925 11033 21959 11067
rect 23673 11033 23707 11067
rect 27169 11033 27203 11067
rect 30113 11033 30147 11067
rect 31401 11033 31435 11067
rect 35725 11033 35759 11067
rect 37473 11033 37507 11067
rect 40325 11033 40359 11067
rect 45845 11033 45879 11067
rect 17233 10965 17267 10999
rect 17969 10965 18003 10999
rect 18429 10965 18463 10999
rect 29101 10965 29135 10999
rect 29285 10965 29319 10999
rect 30757 10965 30791 10999
rect 2237 10761 2271 10795
rect 3985 10761 4019 10795
rect 12265 10761 12299 10795
rect 13185 10761 13219 10795
rect 14381 10761 14415 10795
rect 14749 10761 14783 10795
rect 15945 10761 15979 10795
rect 17141 10761 17175 10795
rect 17509 10761 17543 10795
rect 18337 10761 18371 10795
rect 19533 10761 19567 10795
rect 20729 10761 20763 10795
rect 21097 10761 21131 10795
rect 24225 10761 24259 10795
rect 26341 10761 26375 10795
rect 27537 10761 27571 10795
rect 28549 10761 28583 10795
rect 30573 10761 30607 10795
rect 31401 10761 31435 10795
rect 33057 10761 33091 10795
rect 36829 10761 36863 10795
rect 14841 10693 14875 10727
rect 17601 10693 17635 10727
rect 21189 10693 21223 10727
rect 28827 10693 28861 10727
rect 33333 10693 33367 10727
rect 35357 10693 35391 10727
rect 49157 10693 49191 10727
rect 1593 10625 1627 10659
rect 2697 10625 2731 10659
rect 3801 10625 3835 10659
rect 13553 10625 13587 10659
rect 13645 10625 13679 10659
rect 18705 10625 18739 10659
rect 19901 10625 19935 10659
rect 24593 10625 24627 10659
rect 25421 10625 25455 10659
rect 25973 10625 26007 10659
rect 32689 10625 32723 10659
rect 35633 10625 35667 10659
rect 36461 10625 36495 10659
rect 39773 10625 39807 10659
rect 40233 10625 40267 10659
rect 47961 10625 47995 10659
rect 12541 10557 12575 10591
rect 13829 10557 13863 10591
rect 14933 10557 14967 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 17693 10557 17727 10591
rect 18797 10557 18831 10591
rect 18981 10557 19015 10591
rect 19993 10557 20027 10591
rect 20177 10557 20211 10591
rect 21373 10557 21407 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24685 10557 24719 10591
rect 24869 10557 24903 10591
rect 27353 10557 27387 10591
rect 27445 10557 27479 10591
rect 29561 10557 29595 10591
rect 30389 10557 30423 10591
rect 30481 10557 30515 10591
rect 32413 10557 32447 10591
rect 32597 10557 32631 10591
rect 36185 10557 36219 10591
rect 36369 10557 36403 10591
rect 12725 10489 12759 10523
rect 16865 10489 16899 10523
rect 23765 10489 23799 10523
rect 27905 10489 27939 10523
rect 33885 10489 33919 10523
rect 39957 10489 39991 10523
rect 3341 10421 3375 10455
rect 12081 10421 12115 10455
rect 12909 10421 12943 10455
rect 15577 10421 15611 10455
rect 26065 10421 26099 10455
rect 26525 10421 26559 10455
rect 26801 10421 26835 10455
rect 30941 10421 30975 10455
rect 31861 10421 31895 10455
rect 37289 10421 37323 10455
rect 37473 10421 37507 10455
rect 2191 10217 2225 10251
rect 13461 10217 13495 10251
rect 16681 10217 16715 10251
rect 18153 10217 18187 10251
rect 20269 10217 20303 10251
rect 23765 10217 23799 10251
rect 24593 10217 24627 10251
rect 28733 10217 28767 10251
rect 30389 10217 30423 10251
rect 36645 10217 36679 10251
rect 3801 10149 3835 10183
rect 29009 10149 29043 10183
rect 29377 10149 29411 10183
rect 2421 10081 2455 10115
rect 3985 10081 4019 10115
rect 12909 10081 12943 10115
rect 13001 10081 13035 10115
rect 17417 10081 17451 10115
rect 17601 10081 17635 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 19717 10081 19751 10115
rect 21741 10081 21775 10115
rect 26065 10081 26099 10115
rect 26341 10081 26375 10115
rect 26985 10081 27019 10115
rect 29929 10081 29963 10115
rect 32137 10081 32171 10115
rect 32689 10081 32723 10115
rect 32873 10081 32907 10115
rect 35173 10081 35207 10115
rect 38485 10081 38519 10115
rect 49157 10081 49191 10115
rect 3157 10013 3191 10047
rect 3433 10013 3467 10047
rect 12449 10013 12483 10047
rect 13093 10013 13127 10047
rect 13829 10013 13863 10047
rect 16037 10013 16071 10047
rect 16497 10013 16531 10047
rect 22017 10013 22051 10047
rect 23213 10013 23247 10047
rect 34897 10013 34931 10047
rect 38301 10013 38335 10047
rect 38761 10013 38795 10047
rect 40141 10013 40175 10047
rect 40325 10013 40359 10047
rect 46121 10013 46155 10047
rect 47961 10013 47995 10047
rect 15761 9945 15795 9979
rect 22477 9945 22511 9979
rect 23857 9945 23891 9979
rect 27261 9945 27295 9979
rect 31861 9945 31895 9979
rect 33793 9945 33827 9979
rect 40601 9945 40635 9979
rect 44373 9945 44407 9979
rect 44557 9945 44591 9979
rect 47317 9945 47351 9979
rect 2973 9877 3007 9911
rect 14289 9877 14323 9911
rect 16957 9877 16991 9911
rect 17325 9877 17359 9911
rect 18521 9877 18555 9911
rect 24041 9877 24075 9911
rect 26709 9877 26743 9911
rect 32965 9877 32999 9911
rect 33333 9877 33367 9911
rect 36921 9877 36955 9911
rect 21097 9673 21131 9707
rect 32965 9673 32999 9707
rect 35633 9673 35667 9707
rect 36185 9673 36219 9707
rect 2237 9605 2271 9639
rect 12449 9605 12483 9639
rect 13369 9605 13403 9639
rect 16221 9605 16255 9639
rect 16865 9605 16899 9639
rect 21557 9605 21591 9639
rect 22753 9605 22787 9639
rect 29009 9605 29043 9639
rect 49157 9605 49191 9639
rect 1593 9537 1627 9571
rect 2973 9537 3007 9571
rect 3525 9537 3559 9571
rect 12541 9537 12575 9571
rect 15393 9537 15427 9571
rect 15761 9537 15795 9571
rect 16497 9537 16531 9571
rect 22661 9537 22695 9571
rect 25237 9537 25271 9571
rect 26065 9537 26099 9571
rect 32873 9537 32907 9571
rect 33885 9537 33919 9571
rect 47961 9537 47995 9571
rect 3709 9469 3743 9503
rect 12265 9469 12299 9503
rect 15117 9469 15151 9503
rect 15945 9469 15979 9503
rect 18613 9469 18647 9503
rect 18889 9469 18923 9503
rect 19349 9469 19383 9503
rect 19625 9469 19659 9503
rect 22937 9469 22971 9503
rect 24961 9469 24995 9503
rect 25881 9469 25915 9503
rect 25973 9469 26007 9503
rect 27537 9469 27571 9503
rect 29285 9469 29319 9503
rect 29745 9469 29779 9503
rect 30021 9469 30055 9503
rect 31493 9469 31527 9503
rect 31769 9469 31803 9503
rect 32689 9469 32723 9503
rect 34161 9469 34195 9503
rect 35909 9469 35943 9503
rect 3985 9401 4019 9435
rect 26433 9401 26467 9435
rect 2789 9333 2823 9367
rect 12909 9333 12943 9367
rect 16037 9333 16071 9367
rect 21373 9333 21407 9367
rect 21925 9333 21959 9367
rect 22293 9333 22327 9367
rect 23489 9333 23523 9367
rect 32137 9333 32171 9367
rect 33333 9333 33367 9367
rect 2237 9129 2271 9163
rect 2697 9129 2731 9163
rect 16405 9129 16439 9163
rect 19441 9129 19475 9163
rect 22293 9129 22327 9163
rect 24409 9129 24443 9163
rect 24685 9129 24719 9163
rect 25329 9129 25363 9163
rect 28917 9129 28951 9163
rect 32781 9129 32815 9163
rect 32965 9129 32999 9163
rect 34069 9129 34103 9163
rect 36737 9129 36771 9163
rect 14473 9061 14507 9095
rect 15945 9061 15979 9095
rect 30757 9061 30791 9095
rect 39865 9061 39899 9095
rect 3985 8993 4019 9027
rect 15301 8993 15335 9027
rect 15485 8993 15519 9027
rect 18153 8993 18187 9027
rect 20913 8993 20947 9027
rect 23765 8993 23799 9027
rect 24041 8993 24075 9027
rect 28365 8993 28399 9027
rect 32229 8993 32263 9027
rect 32505 8993 32539 9027
rect 33425 8993 33459 9027
rect 34345 8993 34379 9027
rect 34989 8993 35023 9027
rect 35173 8993 35207 9027
rect 49157 8993 49191 9027
rect 1593 8925 1627 8959
rect 3341 8925 3375 8959
rect 14289 8925 14323 8959
rect 15577 8925 15611 8959
rect 18705 8925 18739 8959
rect 21189 8925 21223 8959
rect 25605 8925 25639 8959
rect 33609 8925 33643 8959
rect 36553 8925 36587 8959
rect 37657 8925 37691 8959
rect 47961 8925 47995 8959
rect 3801 8857 3835 8891
rect 17877 8857 17911 8891
rect 28549 8857 28583 8891
rect 29745 8857 29779 8891
rect 39313 8857 39347 8891
rect 39497 8857 39531 8891
rect 14933 8789 14967 8823
rect 21833 8789 21867 8823
rect 24869 8789 24903 8823
rect 25789 8789 25823 8823
rect 27813 8789 27847 8823
rect 28457 8789 28491 8823
rect 30297 8789 30331 8823
rect 33701 8789 33735 8823
rect 35265 8789 35299 8823
rect 35633 8789 35667 8823
rect 37841 8789 37875 8823
rect 3065 8585 3099 8619
rect 18613 8585 18647 8619
rect 19073 8585 19107 8619
rect 19717 8585 19751 8619
rect 22017 8585 22051 8619
rect 31309 8585 31343 8619
rect 31769 8585 31803 8619
rect 34069 8585 34103 8619
rect 37657 8585 37691 8619
rect 13921 8517 13955 8551
rect 15761 8517 15795 8551
rect 16221 8517 16255 8551
rect 17141 8517 17175 8551
rect 21189 8517 21223 8551
rect 24133 8517 24167 8551
rect 29101 8517 29135 8551
rect 44189 8517 44223 8551
rect 44373 8517 44407 8551
rect 49157 8517 49191 8551
rect 2145 8449 2179 8483
rect 2973 8449 3007 8483
rect 13645 8449 13679 8483
rect 16865 8449 16899 8483
rect 23765 8449 23799 8483
rect 31401 8449 31435 8483
rect 32321 8449 32355 8483
rect 34805 8449 34839 8483
rect 37473 8449 37507 8483
rect 38945 8449 38979 8483
rect 40325 8449 40359 8483
rect 40785 8449 40819 8483
rect 45845 8449 45879 8483
rect 47961 8449 47995 8483
rect 2421 8381 2455 8415
rect 3433 8381 3467 8415
rect 15393 8381 15427 8415
rect 16405 8381 16439 8415
rect 21465 8381 21499 8415
rect 23489 8381 23523 8415
rect 28825 8381 28859 8415
rect 31217 8381 31251 8415
rect 32597 8381 32631 8415
rect 34345 8381 34379 8415
rect 34621 8381 34655 8415
rect 40509 8381 40543 8415
rect 46857 8381 46891 8415
rect 30573 8313 30607 8347
rect 39129 8313 39163 8347
rect 2237 8041 2271 8075
rect 18981 8041 19015 8075
rect 19441 8041 19475 8075
rect 22017 8041 22051 8075
rect 30389 8041 30423 8075
rect 31769 8041 31803 8075
rect 15761 7973 15795 8007
rect 37565 7973 37599 8007
rect 3249 7905 3283 7939
rect 16773 7905 16807 7939
rect 16957 7905 16991 7939
rect 18061 7905 18095 7939
rect 20913 7905 20947 7939
rect 22661 7905 22695 7939
rect 29929 7905 29963 7939
rect 31217 7905 31251 7939
rect 32505 7905 32539 7939
rect 33425 7905 33459 7939
rect 49157 7905 49191 7939
rect 1593 7837 1627 7871
rect 2697 7837 2731 7871
rect 15577 7837 15611 7871
rect 17049 7837 17083 7871
rect 21189 7837 21223 7871
rect 22385 7837 22419 7871
rect 31309 7837 31343 7871
rect 32689 7837 32723 7871
rect 38025 7837 38059 7871
rect 47961 7837 47995 7871
rect 18245 7769 18279 7803
rect 30757 7769 30791 7803
rect 38761 7769 38795 7803
rect 38945 7769 38979 7803
rect 2881 7701 2915 7735
rect 17417 7701 17451 7735
rect 18153 7701 18187 7735
rect 18613 7701 18647 7735
rect 21465 7701 21499 7735
rect 21649 7701 21683 7735
rect 22477 7701 22511 7735
rect 23121 7701 23155 7735
rect 30481 7701 30515 7735
rect 31401 7701 31435 7735
rect 32597 7701 32631 7735
rect 33057 7701 33091 7735
rect 38117 7701 38151 7735
rect 39221 7701 39255 7735
rect 2237 7497 2271 7531
rect 22477 7497 22511 7531
rect 23029 7497 23063 7531
rect 31125 7497 31159 7531
rect 32321 7497 32355 7531
rect 39037 7497 39071 7531
rect 3801 7429 3835 7463
rect 21373 7429 21407 7463
rect 31861 7429 31895 7463
rect 38577 7429 38611 7463
rect 49157 7429 49191 7463
rect 1593 7361 1627 7395
rect 3341 7361 3375 7395
rect 3617 7361 3651 7395
rect 18245 7361 18279 7395
rect 18705 7361 18739 7395
rect 18981 7361 19015 7395
rect 21281 7361 21315 7395
rect 22385 7361 22419 7395
rect 37841 7361 37875 7395
rect 44925 7361 44959 7395
rect 47961 7361 47995 7395
rect 21557 7293 21591 7327
rect 22569 7293 22603 7327
rect 22017 7225 22051 7259
rect 37381 7225 37415 7259
rect 38761 7225 38795 7259
rect 45109 7225 45143 7259
rect 2697 7157 2731 7191
rect 32873 7157 32907 7191
rect 37933 7157 37967 7191
rect 3249 6817 3283 6851
rect 49157 6817 49191 6851
rect 1593 6749 1627 6783
rect 2237 6749 2271 6783
rect 2697 6749 2731 6783
rect 3985 6749 4019 6783
rect 4445 6749 4479 6783
rect 17693 6749 17727 6783
rect 19625 6749 19659 6783
rect 46121 6749 46155 6783
rect 47961 6749 47995 6783
rect 47317 6681 47351 6715
rect 2881 6613 2915 6647
rect 4169 6613 4203 6647
rect 17877 6613 17911 6647
rect 19809 6613 19843 6647
rect 2789 6341 2823 6375
rect 2973 6341 3007 6375
rect 37565 6341 37599 6375
rect 38025 6341 38059 6375
rect 44005 6341 44039 6375
rect 49157 6341 49191 6375
rect 1593 6273 1627 6307
rect 2237 6273 2271 6307
rect 3433 6273 3467 6307
rect 47961 6273 47995 6307
rect 3985 6205 4019 6239
rect 18061 6205 18095 6239
rect 18245 6205 18279 6239
rect 3617 6137 3651 6171
rect 44189 6137 44223 6171
rect 18705 6069 18739 6103
rect 37657 6069 37691 6103
rect 49157 5729 49191 5763
rect 1593 5661 1627 5695
rect 2697 5661 2731 5695
rect 3341 5661 3375 5695
rect 3985 5661 4019 5695
rect 43729 5661 43763 5695
rect 47961 5661 47995 5695
rect 43913 5593 43947 5627
rect 2237 5525 2271 5559
rect 4169 5525 4203 5559
rect 3433 5321 3467 5355
rect 37381 5253 37415 5287
rect 37749 5253 37783 5287
rect 38485 5253 38519 5287
rect 38945 5253 38979 5287
rect 49157 5253 49191 5287
rect 2145 5185 2179 5219
rect 2881 5185 2915 5219
rect 18889 5185 18923 5219
rect 45845 5185 45879 5219
rect 47961 5185 47995 5219
rect 2421 5117 2455 5151
rect 3801 5117 3835 5151
rect 19073 5117 19107 5151
rect 46857 5117 46891 5151
rect 3065 5049 3099 5083
rect 38669 5049 38703 5083
rect 3617 4981 3651 5015
rect 19533 4981 19567 5015
rect 37841 4981 37875 5015
rect 2881 4777 2915 4811
rect 36829 4777 36863 4811
rect 22569 4709 22603 4743
rect 46489 4709 46523 4743
rect 47225 4709 47259 4743
rect 3249 4641 3283 4675
rect 20453 4641 20487 4675
rect 21925 4641 21959 4675
rect 49157 4641 49191 4675
rect 1593 4573 1627 4607
rect 2697 4573 2731 4607
rect 20637 4573 20671 4607
rect 22109 4573 22143 4607
rect 23096 4573 23130 4607
rect 37289 4573 37323 4607
rect 38025 4573 38059 4607
rect 38485 4573 38519 4607
rect 47961 4573 47995 4607
rect 2237 4505 2271 4539
rect 4077 4505 4111 4539
rect 25881 4505 25915 4539
rect 26801 4505 26835 4539
rect 26893 4505 26927 4539
rect 38209 4505 38243 4539
rect 46673 4505 46707 4539
rect 47409 4505 47443 4539
rect 4169 4437 4203 4471
rect 21097 4437 21131 4471
rect 23167 4437 23201 4471
rect 37381 4437 37415 4471
rect 46213 4437 46247 4471
rect 2237 4233 2271 4267
rect 17049 4165 17083 4199
rect 25881 4165 25915 4199
rect 28825 4165 28859 4199
rect 1593 4097 1627 4131
rect 3341 4097 3375 4131
rect 3801 4097 3835 4131
rect 15761 4097 15795 4131
rect 22360 4097 22394 4131
rect 22972 4097 23006 4131
rect 23075 4097 23109 4131
rect 23616 4097 23650 4131
rect 45845 4097 45879 4131
rect 47961 4097 47995 4131
rect 49157 4097 49191 4131
rect 3617 4029 3651 4063
rect 14565 4029 14599 4063
rect 24961 4029 24995 4063
rect 25973 4029 26007 4063
rect 27905 4029 27939 4063
rect 28917 4029 28951 4063
rect 46673 4029 46707 4063
rect 23719 3961 23753 3995
rect 2697 3893 2731 3927
rect 16957 3893 16991 3927
rect 22431 3893 22465 3927
rect 47685 3893 47719 3927
rect 23581 3689 23615 3723
rect 23949 3689 23983 3723
rect 36553 3689 36587 3723
rect 3157 3621 3191 3655
rect 2421 3553 2455 3587
rect 3433 3553 3467 3587
rect 16589 3553 16623 3587
rect 25329 3553 25363 3587
rect 45385 3553 45419 3587
rect 49157 3553 49191 3587
rect 2145 3485 2179 3519
rect 2973 3485 3007 3519
rect 9689 3485 9723 3519
rect 11161 3485 11195 3519
rect 11805 3485 11839 3519
rect 12357 3485 12391 3519
rect 15761 3485 15795 3519
rect 17601 3485 17635 3519
rect 21005 3485 21039 3519
rect 24041 3485 24075 3519
rect 36461 3485 36495 3519
rect 36921 3485 36955 3519
rect 46121 3485 46155 3519
rect 47961 3485 47995 3519
rect 14749 3417 14783 3451
rect 21281 3417 21315 3451
rect 26249 3417 26283 3451
rect 26341 3417 26375 3451
rect 45109 3417 45143 3451
rect 45569 3417 45603 3451
rect 47317 3417 47351 3451
rect 3801 3349 3835 3383
rect 10333 3349 10367 3383
rect 13001 3349 13035 3383
rect 22753 3349 22787 3383
rect 23121 3349 23155 3383
rect 29561 3349 29595 3383
rect 3617 3145 3651 3179
rect 10333 3145 10367 3179
rect 16313 3145 16347 3179
rect 19993 3145 20027 3179
rect 21465 3145 21499 3179
rect 25973 3145 26007 3179
rect 27537 3145 27571 3179
rect 31217 3145 31251 3179
rect 4169 3077 4203 3111
rect 14841 3077 14875 3111
rect 16681 3077 16715 3111
rect 17509 3077 17543 3111
rect 29193 3077 29227 3111
rect 31769 3077 31803 3111
rect 49157 3077 49191 3111
rect 1593 3009 1627 3043
rect 2789 3009 2823 3043
rect 3433 3009 3467 3043
rect 9689 3009 9723 3043
rect 13185 3009 13219 3043
rect 14565 3009 14599 3043
rect 19533 3009 19567 3043
rect 20177 3009 20211 3043
rect 20637 3009 20671 3043
rect 21281 3009 21315 3043
rect 22661 3009 22695 3043
rect 23765 3009 23799 3043
rect 26433 3009 26467 3043
rect 27997 3009 28031 3043
rect 28917 3009 28951 3043
rect 31401 3009 31435 3043
rect 33149 3009 33183 3043
rect 35265 3009 35299 3043
rect 38025 3009 38059 3043
rect 44005 3009 44039 3043
rect 45845 3009 45879 3043
rect 47961 3009 47995 3043
rect 2237 2941 2271 2975
rect 11989 2941 12023 2975
rect 17325 2941 17359 2975
rect 18337 2941 18371 2975
rect 24225 2941 24259 2975
rect 24501 2941 24535 2975
rect 38301 2941 38335 2975
rect 45201 2941 45235 2975
rect 46857 2941 46891 2975
rect 2973 2873 3007 2907
rect 20821 2873 20855 2907
rect 22201 2873 22235 2907
rect 32965 2873 32999 2907
rect 3985 2805 4019 2839
rect 9413 2805 9447 2839
rect 22385 2805 22419 2839
rect 23305 2805 23339 2839
rect 23489 2805 23523 2839
rect 26617 2805 26651 2839
rect 27905 2805 27939 2839
rect 30665 2805 30699 2839
rect 35081 2805 35115 2839
rect 2237 2601 2271 2635
rect 9597 2601 9631 2635
rect 26341 2601 26375 2635
rect 29009 2601 29043 2635
rect 31585 2601 31619 2635
rect 33701 2601 33735 2635
rect 35817 2601 35851 2635
rect 38117 2601 38151 2635
rect 4169 2533 4203 2567
rect 13277 2465 13311 2499
rect 15301 2465 15335 2499
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 25053 2465 25087 2499
rect 27629 2465 27663 2499
rect 41429 2465 41463 2499
rect 43821 2465 43855 2499
rect 49157 2465 49191 2499
rect 1593 2397 1627 2431
rect 2697 2397 2731 2431
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 9413 2397 9447 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 13737 2397 13771 2431
rect 16313 2397 16347 2431
rect 18245 2397 18279 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 22385 2397 22419 2431
rect 24593 2397 24627 2431
rect 27169 2397 27203 2431
rect 29193 2397 29227 2431
rect 29745 2397 29779 2431
rect 30941 2397 30975 2431
rect 31861 2397 31895 2431
rect 33057 2397 33091 2431
rect 35173 2397 35207 2431
rect 37473 2397 37507 2431
rect 40693 2397 40727 2431
rect 43545 2397 43579 2431
rect 45845 2397 45879 2431
rect 47961 2397 47995 2431
rect 17049 2329 17083 2363
rect 30389 2329 30423 2363
rect 47041 2329 47075 2363
rect 4905 2261 4939 2295
rect 18705 2261 18739 2295
rect 19625 2261 19659 2295
rect 32781 2261 32815 2295
rect 34897 2261 34931 2295
rect 37105 2261 37139 2295
rect 43269 2261 43303 2295
<< metal1 >>
rect 34054 26324 34060 26376
rect 34112 26364 34118 26376
rect 43346 26364 43352 26376
rect 34112 26336 43352 26364
rect 34112 26324 34118 26336
rect 43346 26324 43352 26336
rect 43404 26324 43410 26376
rect 4062 25168 4068 25220
rect 4120 25208 4126 25220
rect 9766 25208 9772 25220
rect 4120 25180 9772 25208
rect 4120 25168 4126 25180
rect 9766 25168 9772 25180
rect 9824 25168 9830 25220
rect 21542 24828 21548 24880
rect 21600 24868 21606 24880
rect 25958 24868 25964 24880
rect 21600 24840 25964 24868
rect 21600 24828 21606 24840
rect 25958 24828 25964 24840
rect 26016 24828 26022 24880
rect 16022 24760 16028 24812
rect 16080 24800 16086 24812
rect 24486 24800 24492 24812
rect 16080 24772 24492 24800
rect 16080 24760 16086 24772
rect 24486 24760 24492 24772
rect 24544 24760 24550 24812
rect 26326 24800 26332 24812
rect 24596 24772 26332 24800
rect 18874 24692 18880 24744
rect 18932 24732 18938 24744
rect 24596 24732 24624 24772
rect 26326 24760 26332 24772
rect 26384 24760 26390 24812
rect 26418 24760 26424 24812
rect 26476 24800 26482 24812
rect 35158 24800 35164 24812
rect 26476 24772 35164 24800
rect 26476 24760 26482 24772
rect 35158 24760 35164 24772
rect 35216 24760 35222 24812
rect 40586 24800 40592 24812
rect 35268 24772 40592 24800
rect 18932 24704 24624 24732
rect 18932 24692 18938 24704
rect 29546 24692 29552 24744
rect 29604 24732 29610 24744
rect 32858 24732 32864 24744
rect 29604 24704 32864 24732
rect 29604 24692 29610 24704
rect 32858 24692 32864 24704
rect 32916 24692 32922 24744
rect 34974 24692 34980 24744
rect 35032 24732 35038 24744
rect 35268 24732 35296 24772
rect 40586 24760 40592 24772
rect 40644 24760 40650 24812
rect 35032 24704 35296 24732
rect 35032 24692 35038 24704
rect 35526 24692 35532 24744
rect 35584 24732 35590 24744
rect 35584 24704 38976 24732
rect 35584 24692 35590 24704
rect 24762 24624 24768 24676
rect 24820 24664 24826 24676
rect 30374 24664 30380 24676
rect 24820 24636 30380 24664
rect 24820 24624 24826 24636
rect 30374 24624 30380 24636
rect 30432 24624 30438 24676
rect 30558 24624 30564 24676
rect 30616 24664 30622 24676
rect 38838 24664 38844 24676
rect 30616 24636 38844 24664
rect 30616 24624 30622 24636
rect 38838 24624 38844 24636
rect 38896 24624 38902 24676
rect 38948 24664 38976 24704
rect 39206 24692 39212 24744
rect 39264 24732 39270 24744
rect 43898 24732 43904 24744
rect 39264 24704 43904 24732
rect 39264 24692 39270 24704
rect 43898 24692 43904 24704
rect 43956 24692 43962 24744
rect 39390 24664 39396 24676
rect 38948 24636 39396 24664
rect 39390 24624 39396 24636
rect 39448 24624 39454 24676
rect 39574 24624 39580 24676
rect 39632 24664 39638 24676
rect 44358 24664 44364 24676
rect 39632 24636 44364 24664
rect 39632 24624 39638 24636
rect 44358 24624 44364 24636
rect 44416 24624 44422 24676
rect 45554 24624 45560 24676
rect 45612 24664 45618 24676
rect 46750 24664 46756 24676
rect 45612 24636 46756 24664
rect 45612 24624 45618 24636
rect 46750 24624 46756 24636
rect 46808 24624 46814 24676
rect 3602 24556 3608 24608
rect 3660 24596 3666 24608
rect 6546 24596 6552 24608
rect 3660 24568 6552 24596
rect 3660 24556 3666 24568
rect 6546 24556 6552 24568
rect 6604 24556 6610 24608
rect 20806 24556 20812 24608
rect 20864 24596 20870 24608
rect 29730 24596 29736 24608
rect 20864 24568 29736 24596
rect 20864 24556 20870 24568
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 31846 24556 31852 24608
rect 31904 24596 31910 24608
rect 39482 24596 39488 24608
rect 31904 24568 39488 24596
rect 31904 24556 31910 24568
rect 39482 24556 39488 24568
rect 39540 24556 39546 24608
rect 40402 24556 40408 24608
rect 40460 24596 40466 24608
rect 47118 24596 47124 24608
rect 40460 24568 47124 24596
rect 40460 24556 40466 24568
rect 47118 24556 47124 24568
rect 47176 24556 47182 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 19058 24352 19064 24404
rect 19116 24392 19122 24404
rect 19116 24364 25268 24392
rect 19116 24352 19122 24364
rect 9858 24324 9864 24336
rect 3988 24296 9864 24324
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 3510 24256 3516 24268
rect 3007 24228 3516 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 3421 24191 3479 24197
rect 3421 24157 3433 24191
rect 3467 24188 3479 24191
rect 3878 24188 3884 24200
rect 3467 24160 3884 24188
rect 3467 24157 3479 24160
rect 3421 24151 3479 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 3988 24197 4016 24296
rect 9858 24284 9864 24296
rect 9916 24284 9922 24336
rect 11882 24324 11888 24336
rect 10704 24296 11888 24324
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6730 24256 6736 24268
rect 5859 24228 6736 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6730 24216 6736 24228
rect 6788 24216 6794 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8662 24256 8668 24268
rect 8251 24228 8668 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 10704 24265 10732 24296
rect 11882 24284 11888 24296
rect 11940 24284 11946 24336
rect 19610 24324 19616 24336
rect 18432 24296 19616 24324
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24225 10747 24259
rect 12342 24256 12348 24268
rect 10689 24219 10747 24225
rect 11164 24228 12348 24256
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24157 6607 24191
rect 6549 24151 6607 24157
rect 2314 24080 2320 24132
rect 2372 24120 2378 24132
rect 4632 24120 4660 24151
rect 2372 24092 4660 24120
rect 6564 24120 6592 24151
rect 7098 24148 7104 24200
rect 7156 24188 7162 24200
rect 7377 24191 7435 24197
rect 7377 24188 7389 24191
rect 7156 24160 7389 24188
rect 7156 24148 7162 24160
rect 7377 24157 7389 24160
rect 7423 24188 7435 24191
rect 7466 24188 7472 24200
rect 7423 24160 7472 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 7466 24148 7472 24160
rect 7524 24148 7530 24200
rect 11164 24197 11192 24228
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 13265 24259 13323 24265
rect 13265 24225 13277 24259
rect 13311 24256 13323 24259
rect 13814 24256 13820 24268
rect 13311 24228 13820 24256
rect 13311 24225 13323 24228
rect 13265 24219 13323 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 15841 24259 15899 24265
rect 15841 24225 15853 24259
rect 15887 24256 15899 24259
rect 17678 24256 17684 24268
rect 15887 24228 17684 24256
rect 15887 24225 15899 24228
rect 15841 24219 15899 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 18432 24265 18460 24296
rect 19610 24284 19616 24296
rect 19668 24284 19674 24336
rect 20254 24284 20260 24336
rect 20312 24324 20318 24336
rect 20312 24296 22094 24324
rect 20312 24284 20318 24296
rect 18417 24259 18475 24265
rect 18417 24225 18429 24259
rect 18463 24225 18475 24259
rect 20622 24256 20628 24268
rect 18417 24219 18475 24225
rect 18524 24228 20628 24256
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 11149 24191 11207 24197
rect 9355 24160 10916 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9582 24120 9588 24132
rect 6564 24092 9588 24120
rect 2372 24080 2378 24092
rect 9582 24080 9588 24092
rect 9640 24080 9646 24132
rect 10888 24120 10916 24160
rect 11149 24157 11161 24191
rect 11195 24157 11207 24191
rect 11149 24151 11207 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 13630 24188 13636 24200
rect 11931 24160 13636 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 13722 24148 13728 24200
rect 13780 24148 13786 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24188 16359 24191
rect 18524 24188 18552 24228
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 22066 24256 22094 24296
rect 24486 24284 24492 24336
rect 24544 24324 24550 24336
rect 24581 24327 24639 24333
rect 24581 24324 24593 24327
rect 24544 24296 24593 24324
rect 24544 24284 24550 24296
rect 24581 24293 24593 24296
rect 24627 24293 24639 24327
rect 24581 24287 24639 24293
rect 25240 24265 25268 24364
rect 26418 24352 26424 24404
rect 26476 24352 26482 24404
rect 29730 24352 29736 24404
rect 29788 24352 29794 24404
rect 30190 24352 30196 24404
rect 30248 24392 30254 24404
rect 35894 24392 35900 24404
rect 30248 24364 35900 24392
rect 30248 24352 30254 24364
rect 35894 24352 35900 24364
rect 35952 24352 35958 24404
rect 37550 24352 37556 24404
rect 37608 24392 37614 24404
rect 39301 24395 39359 24401
rect 39301 24392 39313 24395
rect 37608 24364 39313 24392
rect 37608 24352 37614 24364
rect 39301 24361 39313 24364
rect 39347 24361 39359 24395
rect 39301 24355 39359 24361
rect 39390 24352 39396 24404
rect 39448 24392 39454 24404
rect 42613 24395 42671 24401
rect 42613 24392 42625 24395
rect 39448 24364 42625 24392
rect 39448 24352 39454 24364
rect 42613 24361 42625 24364
rect 42659 24361 42671 24395
rect 44266 24392 44272 24404
rect 42613 24355 42671 24361
rect 42996 24364 44272 24392
rect 25774 24284 25780 24336
rect 25832 24284 25838 24336
rect 26326 24284 26332 24336
rect 26384 24324 26390 24336
rect 27157 24327 27215 24333
rect 27157 24324 27169 24327
rect 26384 24296 27169 24324
rect 26384 24284 26390 24296
rect 27157 24293 27169 24296
rect 27203 24293 27215 24327
rect 27157 24287 27215 24293
rect 28626 24284 28632 24336
rect 28684 24324 28690 24336
rect 28684 24296 30512 24324
rect 28684 24284 28690 24296
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 22066 24228 22477 24256
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 25225 24259 25283 24265
rect 25225 24225 25237 24259
rect 25271 24225 25283 24259
rect 26602 24256 26608 24268
rect 25225 24219 25283 24225
rect 25516 24228 26608 24256
rect 16347 24160 18552 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 18874 24148 18880 24200
rect 18932 24148 18938 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 20806 24188 20812 24200
rect 19659 24160 20812 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 20806 24148 20812 24160
rect 20864 24148 20870 24200
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 15562 24120 15568 24132
rect 10888 24092 15568 24120
rect 15562 24080 15568 24092
rect 15620 24080 15626 24132
rect 17218 24080 17224 24132
rect 17276 24120 17282 24132
rect 21376 24120 21404 24151
rect 21450 24148 21456 24200
rect 21508 24188 21514 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21508 24160 22017 24188
rect 21508 24148 21514 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 23845 24191 23903 24197
rect 23845 24157 23857 24191
rect 23891 24188 23903 24191
rect 25406 24188 25412 24200
rect 23891 24160 25412 24188
rect 23891 24157 23903 24160
rect 23845 24151 23903 24157
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 22646 24120 22652 24132
rect 17276 24092 19564 24120
rect 21376 24092 22652 24120
rect 17276 24080 17282 24092
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24052 4215 24055
rect 6638 24052 6644 24064
rect 4203 24024 6644 24052
rect 4203 24021 4215 24024
rect 4157 24015 4215 24021
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 6733 24055 6791 24061
rect 6733 24021 6745 24055
rect 6779 24052 6791 24055
rect 7466 24052 7472 24064
rect 6779 24024 7472 24052
rect 6779 24021 6791 24024
rect 6733 24015 6791 24021
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 11146 24012 11152 24064
rect 11204 24052 11210 24064
rect 11701 24055 11759 24061
rect 11701 24052 11713 24055
rect 11204 24024 11713 24052
rect 11204 24012 11210 24024
rect 11701 24021 11713 24024
rect 11747 24021 11759 24055
rect 11701 24015 11759 24021
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 11848 24024 14289 24052
rect 11848 24012 11854 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 17037 24055 17095 24061
rect 17037 24021 17049 24055
rect 17083 24052 17095 24055
rect 18598 24052 18604 24064
rect 17083 24024 18604 24052
rect 17083 24021 17095 24024
rect 17037 24015 17095 24021
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 19536 24052 19564 24092
rect 22646 24080 22652 24092
rect 22704 24080 22710 24132
rect 24949 24123 25007 24129
rect 24949 24089 24961 24123
rect 24995 24120 25007 24123
rect 25314 24120 25320 24132
rect 24995 24092 25320 24120
rect 24995 24089 25007 24092
rect 24949 24083 25007 24089
rect 25314 24080 25320 24092
rect 25372 24080 25378 24132
rect 23934 24052 23940 24064
rect 19536 24024 23940 24052
rect 23934 24012 23940 24024
rect 23992 24012 23998 24064
rect 24029 24055 24087 24061
rect 24029 24021 24041 24055
rect 24075 24052 24087 24055
rect 24854 24052 24860 24064
rect 24075 24024 24860 24052
rect 24075 24021 24087 24024
rect 24029 24015 24087 24021
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25516 24052 25544 24228
rect 26602 24216 26608 24228
rect 26660 24216 26666 24268
rect 27338 24216 27344 24268
rect 27396 24256 27402 24268
rect 29181 24259 29239 24265
rect 29181 24256 29193 24259
rect 27396 24228 29193 24256
rect 27396 24216 27402 24228
rect 26050 24148 26056 24200
rect 26108 24188 26114 24200
rect 28552 24197 28580 24228
rect 29181 24225 29193 24228
rect 29227 24225 29239 24259
rect 29181 24219 29239 24225
rect 27893 24191 27951 24197
rect 27893 24188 27905 24191
rect 26108 24160 27905 24188
rect 26108 24148 26114 24160
rect 27893 24157 27905 24160
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24157 29975 24191
rect 29917 24151 29975 24157
rect 25961 24123 26019 24129
rect 25961 24089 25973 24123
rect 26007 24120 26019 24123
rect 26418 24120 26424 24132
rect 26007 24092 26424 24120
rect 26007 24089 26019 24092
rect 25961 24083 26019 24089
rect 26418 24080 26424 24092
rect 26476 24080 26482 24132
rect 26789 24123 26847 24129
rect 26789 24089 26801 24123
rect 26835 24120 26847 24123
rect 27246 24120 27252 24132
rect 26835 24092 27252 24120
rect 26835 24089 26847 24092
rect 26789 24083 26847 24089
rect 27246 24080 27252 24092
rect 27304 24080 27310 24132
rect 27338 24080 27344 24132
rect 27396 24080 27402 24132
rect 27908 24120 27936 24151
rect 28997 24123 29055 24129
rect 28997 24120 29009 24123
rect 27908 24092 29009 24120
rect 28997 24089 29009 24092
rect 29043 24089 29055 24123
rect 29932 24120 29960 24151
rect 30374 24148 30380 24200
rect 30432 24148 30438 24200
rect 30484 24188 30512 24296
rect 30558 24284 30564 24336
rect 30616 24324 30622 24336
rect 30616 24296 31156 24324
rect 30616 24284 30622 24296
rect 31128 24256 31156 24296
rect 31294 24284 31300 24336
rect 31352 24324 31358 24336
rect 32953 24327 33011 24333
rect 32953 24324 32965 24327
rect 31352 24296 32965 24324
rect 31352 24284 31358 24296
rect 32953 24293 32965 24296
rect 32999 24293 33011 24327
rect 32953 24287 33011 24293
rect 33042 24284 33048 24336
rect 33100 24324 33106 24336
rect 36446 24324 36452 24336
rect 33100 24296 36452 24324
rect 33100 24284 33106 24296
rect 36446 24284 36452 24296
rect 36504 24284 36510 24336
rect 38197 24327 38255 24333
rect 36556 24296 38148 24324
rect 31481 24259 31539 24265
rect 31481 24256 31493 24259
rect 31128 24228 31493 24256
rect 31481 24225 31493 24228
rect 31527 24225 31539 24259
rect 31481 24219 31539 24225
rect 31570 24216 31576 24268
rect 31628 24256 31634 24268
rect 31941 24259 31999 24265
rect 31941 24256 31953 24259
rect 31628 24228 31953 24256
rect 31628 24216 31634 24228
rect 31941 24225 31953 24228
rect 31987 24256 31999 24259
rect 32766 24256 32772 24268
rect 31987 24228 32772 24256
rect 31987 24225 31999 24228
rect 31941 24219 31999 24225
rect 32766 24216 32772 24228
rect 32824 24216 32830 24268
rect 34241 24259 34299 24265
rect 34241 24225 34253 24259
rect 34287 24256 34299 24259
rect 34330 24256 34336 24268
rect 34287 24228 34336 24256
rect 34287 24225 34299 24228
rect 34241 24219 34299 24225
rect 34330 24216 34336 24228
rect 34388 24216 34394 24268
rect 34974 24216 34980 24268
rect 35032 24216 35038 24268
rect 35158 24216 35164 24268
rect 35216 24216 35222 24268
rect 36556 24265 36584 24296
rect 36541 24259 36599 24265
rect 36541 24225 36553 24259
rect 36587 24225 36599 24259
rect 36541 24219 36599 24225
rect 36722 24216 36728 24268
rect 36780 24216 36786 24268
rect 37458 24216 37464 24268
rect 37516 24256 37522 24268
rect 37553 24259 37611 24265
rect 37553 24256 37565 24259
rect 37516 24228 37565 24256
rect 37516 24216 37522 24228
rect 37553 24225 37565 24228
rect 37599 24225 37611 24259
rect 38120 24256 38148 24296
rect 38197 24293 38209 24327
rect 38243 24324 38255 24327
rect 38654 24324 38660 24336
rect 38243 24296 38660 24324
rect 38243 24293 38255 24296
rect 38197 24287 38255 24293
rect 38654 24284 38660 24296
rect 38712 24284 38718 24336
rect 42886 24324 42892 24336
rect 41386 24296 42892 24324
rect 40126 24256 40132 24268
rect 37553 24219 37611 24225
rect 37752 24228 37964 24256
rect 38120 24228 40132 24256
rect 31021 24191 31079 24197
rect 31021 24188 31033 24191
rect 30484 24160 31033 24188
rect 31021 24157 31033 24160
rect 31067 24188 31079 24191
rect 31665 24191 31723 24197
rect 31665 24188 31677 24191
rect 31067 24160 31677 24188
rect 31067 24157 31079 24160
rect 31021 24151 31079 24157
rect 31665 24157 31677 24160
rect 31711 24157 31723 24191
rect 31665 24151 31723 24157
rect 32493 24191 32551 24197
rect 32493 24157 32505 24191
rect 32539 24188 32551 24191
rect 32858 24188 32864 24200
rect 32539 24160 32864 24188
rect 32539 24157 32551 24160
rect 32493 24151 32551 24157
rect 32858 24148 32864 24160
rect 32916 24148 32922 24200
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24188 33195 24191
rect 33318 24188 33324 24200
rect 33183 24160 33324 24188
rect 33183 24157 33195 24160
rect 33137 24151 33195 24157
rect 33318 24148 33324 24160
rect 33376 24148 33382 24200
rect 33870 24148 33876 24200
rect 33928 24188 33934 24200
rect 34992 24188 35020 24216
rect 33928 24160 35020 24188
rect 35176 24188 35204 24216
rect 37752 24197 37780 24228
rect 37737 24191 37795 24197
rect 37737 24188 37749 24191
rect 35176 24184 37596 24188
rect 37660 24184 37749 24188
rect 35176 24160 37749 24184
rect 33928 24148 33934 24160
rect 37568 24156 37688 24160
rect 37737 24157 37749 24160
rect 37783 24157 37795 24191
rect 37737 24151 37795 24157
rect 33965 24123 34023 24129
rect 29932 24092 33640 24120
rect 28997 24083 29055 24089
rect 25087 24024 25544 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 26970 24012 26976 24064
rect 27028 24052 27034 24064
rect 27798 24052 27804 24064
rect 27028 24024 27804 24052
rect 27028 24012 27034 24024
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 28077 24055 28135 24061
rect 28077 24021 28089 24055
rect 28123 24052 28135 24055
rect 28350 24052 28356 24064
rect 28123 24024 28356 24052
rect 28123 24021 28135 24024
rect 28077 24015 28135 24021
rect 28350 24012 28356 24024
rect 28408 24012 28414 24064
rect 28626 24012 28632 24064
rect 28684 24052 28690 24064
rect 28721 24055 28779 24061
rect 28721 24052 28733 24055
rect 28684 24024 28733 24052
rect 28684 24012 28690 24024
rect 28721 24021 28733 24024
rect 28767 24021 28779 24055
rect 28721 24015 28779 24021
rect 30558 24012 30564 24064
rect 30616 24012 30622 24064
rect 31110 24012 31116 24064
rect 31168 24052 31174 24064
rect 31205 24055 31263 24061
rect 31205 24052 31217 24055
rect 31168 24024 31217 24052
rect 31168 24012 31174 24024
rect 31205 24021 31217 24024
rect 31251 24021 31263 24055
rect 31205 24015 31263 24021
rect 32306 24012 32312 24064
rect 32364 24012 32370 24064
rect 33612 24061 33640 24092
rect 33965 24089 33977 24123
rect 34011 24120 34023 24123
rect 34422 24120 34428 24132
rect 34011 24092 34428 24120
rect 34011 24089 34023 24092
rect 33965 24083 34023 24089
rect 34422 24080 34428 24092
rect 34480 24080 34486 24132
rect 37936 24120 37964 24228
rect 40126 24216 40132 24228
rect 40184 24216 40190 24268
rect 40586 24216 40592 24268
rect 40644 24216 40650 24268
rect 38838 24148 38844 24200
rect 38896 24148 38902 24200
rect 39482 24148 39488 24200
rect 39540 24148 39546 24200
rect 40402 24148 40408 24200
rect 40460 24148 40466 24200
rect 41049 24123 41107 24129
rect 41049 24120 41061 24123
rect 37936 24092 41061 24120
rect 41049 24089 41061 24092
rect 41095 24120 41107 24123
rect 41386 24120 41414 24296
rect 42886 24284 42892 24296
rect 42944 24284 42950 24336
rect 42150 24256 42156 24268
rect 42076 24228 42156 24256
rect 42076 24197 42104 24228
rect 42150 24216 42156 24228
rect 42208 24256 42214 24268
rect 42996 24256 43024 24364
rect 44266 24352 44272 24364
rect 44324 24352 44330 24404
rect 46290 24352 46296 24404
rect 46348 24392 46354 24404
rect 47581 24395 47639 24401
rect 47581 24392 47593 24395
rect 46348 24364 47593 24392
rect 46348 24352 46354 24364
rect 47581 24361 47593 24364
rect 47627 24392 47639 24395
rect 47854 24392 47860 24404
rect 47627 24364 47860 24392
rect 47627 24361 47639 24364
rect 47581 24355 47639 24361
rect 47854 24352 47860 24364
rect 47912 24352 47918 24404
rect 43530 24284 43536 24336
rect 43588 24324 43594 24336
rect 43588 24296 45968 24324
rect 43588 24284 43594 24296
rect 45833 24259 45891 24265
rect 45833 24256 45845 24259
rect 42208 24228 43024 24256
rect 44376 24228 45845 24256
rect 42208 24216 42214 24228
rect 42061 24191 42119 24197
rect 42061 24157 42073 24191
rect 42107 24157 42119 24191
rect 42061 24151 42119 24157
rect 42797 24191 42855 24197
rect 42797 24157 42809 24191
rect 42843 24188 42855 24191
rect 43346 24188 43352 24200
rect 42843 24160 43352 24188
rect 42843 24157 42855 24160
rect 42797 24151 42855 24157
rect 43346 24148 43352 24160
rect 43404 24148 43410 24200
rect 43441 24191 43499 24197
rect 43441 24157 43453 24191
rect 43487 24188 43499 24191
rect 43530 24188 43536 24200
rect 43487 24160 43536 24188
rect 43487 24157 43499 24160
rect 43441 24151 43499 24157
rect 43530 24148 43536 24160
rect 43588 24148 43594 24200
rect 44376 24197 44404 24228
rect 45833 24225 45845 24228
rect 45879 24225 45891 24259
rect 45940 24256 45968 24296
rect 46750 24284 46756 24336
rect 46808 24324 46814 24336
rect 46808 24296 48360 24324
rect 46808 24284 46814 24296
rect 47213 24259 47271 24265
rect 47213 24256 47225 24259
rect 45940 24228 47225 24256
rect 45833 24219 45891 24225
rect 47213 24225 47225 24228
rect 47259 24225 47271 24259
rect 47213 24219 47271 24225
rect 44361 24191 44419 24197
rect 44361 24157 44373 24191
rect 44407 24157 44419 24191
rect 44361 24151 44419 24157
rect 44450 24148 44456 24200
rect 44508 24188 44514 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44508 24160 45201 24188
rect 44508 24148 44514 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 46937 24191 46995 24197
rect 46937 24157 46949 24191
rect 46983 24157 46995 24191
rect 46937 24151 46995 24157
rect 41095 24092 41414 24120
rect 41095 24089 41107 24092
rect 41049 24083 41107 24089
rect 42150 24080 42156 24132
rect 42208 24120 42214 24132
rect 43717 24123 43775 24129
rect 43717 24120 43729 24123
rect 42208 24092 43729 24120
rect 42208 24080 42214 24092
rect 43717 24089 43729 24092
rect 43763 24089 43775 24123
rect 43717 24083 43775 24089
rect 44726 24080 44732 24132
rect 44784 24120 44790 24132
rect 46952 24120 46980 24151
rect 47670 24148 47676 24200
rect 47728 24188 47734 24200
rect 48225 24191 48283 24197
rect 48225 24188 48237 24191
rect 47728 24160 48237 24188
rect 47728 24148 47734 24160
rect 48225 24157 48237 24160
rect 48271 24157 48283 24191
rect 48332 24188 48360 24296
rect 48961 24191 49019 24197
rect 48961 24188 48973 24191
rect 48332 24160 48973 24188
rect 48225 24151 48283 24157
rect 48961 24157 48973 24160
rect 49007 24188 49019 24191
rect 49421 24191 49479 24197
rect 49421 24188 49433 24191
rect 49007 24160 49433 24188
rect 49007 24157 49019 24160
rect 48961 24151 49019 24157
rect 49421 24157 49433 24160
rect 49467 24157 49479 24191
rect 49421 24151 49479 24157
rect 49237 24123 49295 24129
rect 49237 24120 49249 24123
rect 44784 24092 49249 24120
rect 44784 24080 44790 24092
rect 49237 24089 49249 24092
rect 49283 24089 49295 24123
rect 49237 24083 49295 24089
rect 33597 24055 33655 24061
rect 33597 24021 33609 24055
rect 33643 24021 33655 24055
rect 33597 24015 33655 24021
rect 34054 24012 34060 24064
rect 34112 24012 34118 24064
rect 35250 24012 35256 24064
rect 35308 24012 35314 24064
rect 35618 24012 35624 24064
rect 35676 24012 35682 24064
rect 36078 24012 36084 24064
rect 36136 24012 36142 24064
rect 36449 24055 36507 24061
rect 36449 24021 36461 24055
rect 36495 24052 36507 24055
rect 36814 24052 36820 24064
rect 36495 24024 36820 24052
rect 36495 24021 36507 24024
rect 36449 24015 36507 24021
rect 36814 24012 36820 24024
rect 36872 24012 36878 24064
rect 37826 24012 37832 24064
rect 37884 24012 37890 24064
rect 38378 24012 38384 24064
rect 38436 24052 38442 24064
rect 38657 24055 38715 24061
rect 38657 24052 38669 24055
rect 38436 24024 38669 24052
rect 38436 24012 38442 24024
rect 38657 24021 38669 24024
rect 38703 24021 38715 24055
rect 38657 24015 38715 24021
rect 40034 24012 40040 24064
rect 40092 24012 40098 24064
rect 40497 24055 40555 24061
rect 40497 24021 40509 24055
rect 40543 24052 40555 24055
rect 40954 24052 40960 24064
rect 40543 24024 40960 24052
rect 40543 24021 40555 24024
rect 40497 24015 40555 24021
rect 40954 24012 40960 24024
rect 41012 24012 41018 24064
rect 41417 24055 41475 24061
rect 41417 24021 41429 24055
rect 41463 24052 41475 24055
rect 42610 24052 42616 24064
rect 41463 24024 42616 24052
rect 41463 24021 41475 24024
rect 41417 24015 41475 24021
rect 42610 24012 42616 24024
rect 42668 24012 42674 24064
rect 42794 24012 42800 24064
rect 42852 24052 42858 24064
rect 43257 24055 43315 24061
rect 43257 24052 43269 24055
rect 42852 24024 43269 24052
rect 42852 24012 42858 24024
rect 43257 24021 43269 24024
rect 43303 24021 43315 24055
rect 43257 24015 43315 24021
rect 44174 24012 44180 24064
rect 44232 24012 44238 24064
rect 44634 24012 44640 24064
rect 44692 24012 44698 24064
rect 45370 24012 45376 24064
rect 45428 24052 45434 24064
rect 46293 24055 46351 24061
rect 46293 24052 46305 24055
rect 45428 24024 46305 24052
rect 45428 24012 45434 24024
rect 46293 24021 46305 24024
rect 46339 24021 46351 24055
rect 46293 24015 46351 24021
rect 48038 24012 48044 24064
rect 48096 24012 48102 24064
rect 48774 24012 48780 24064
rect 48832 24012 48838 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 2314 23808 2320 23860
rect 2372 23808 2378 23860
rect 7469 23851 7527 23857
rect 7469 23817 7481 23851
rect 7515 23848 7527 23851
rect 19610 23848 19616 23860
rect 7515 23820 12434 23848
rect 7515 23817 7527 23820
rect 7469 23811 7527 23817
rect 11790 23780 11796 23792
rect 2148 23752 6592 23780
rect 2148 23721 2176 23752
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 4062 23672 4068 23724
rect 4120 23672 4126 23724
rect 4706 23672 4712 23724
rect 4764 23672 4770 23724
rect 3697 23647 3755 23653
rect 3697 23613 3709 23647
rect 3743 23644 3755 23647
rect 4154 23644 4160 23656
rect 3743 23616 4160 23644
rect 3743 23613 3755 23616
rect 3697 23607 3755 23613
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 3970 23536 3976 23588
rect 4028 23576 4034 23588
rect 5810 23576 5816 23588
rect 4028 23548 5816 23576
rect 4028 23536 4034 23548
rect 5810 23536 5816 23548
rect 5868 23536 5874 23588
rect 6564 23576 6592 23752
rect 9324 23752 11796 23780
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 7285 23715 7343 23721
rect 7285 23681 7297 23715
rect 7331 23712 7343 23715
rect 8570 23712 8576 23724
rect 7331 23684 8576 23712
rect 7331 23681 7343 23684
rect 7285 23675 7343 23681
rect 6840 23644 6868 23675
rect 8570 23672 8576 23684
rect 8628 23672 8634 23724
rect 9324 23721 9352 23752
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23712 11207 23715
rect 12158 23712 12164 23724
rect 11195 23684 12164 23712
rect 11195 23681 11207 23684
rect 11149 23675 11207 23681
rect 12158 23672 12164 23684
rect 12216 23672 12222 23724
rect 12406 23712 12434 23820
rect 16316 23820 19616 23848
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 14366 23780 14372 23792
rect 14323 23752 14372 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 14366 23740 14372 23752
rect 14424 23740 14430 23792
rect 16316 23721 16344 23820
rect 19610 23808 19616 23820
rect 19668 23808 19674 23860
rect 21450 23808 21456 23860
rect 21508 23808 21514 23860
rect 28445 23851 28503 23857
rect 28445 23848 28457 23851
rect 22066 23820 28457 23848
rect 19242 23740 19248 23792
rect 19300 23740 19306 23792
rect 20257 23783 20315 23789
rect 20257 23749 20269 23783
rect 20303 23780 20315 23783
rect 20346 23780 20352 23792
rect 20303 23752 20352 23780
rect 20303 23749 20315 23752
rect 20257 23743 20315 23749
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 22066 23780 22094 23820
rect 28445 23817 28457 23820
rect 28491 23817 28503 23851
rect 32309 23851 32367 23857
rect 32309 23848 32321 23851
rect 28445 23811 28503 23817
rect 28644 23820 32321 23848
rect 23474 23780 23480 23792
rect 21468 23752 22094 23780
rect 22848 23752 23480 23780
rect 13081 23715 13139 23721
rect 13081 23712 13093 23715
rect 12406 23684 13093 23712
rect 13081 23681 13093 23684
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23681 16359 23715
rect 16301 23675 16359 23681
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 21269 23715 21327 23721
rect 18279 23684 19104 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 8386 23644 8392 23656
rect 6840 23616 8392 23644
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 8849 23647 8907 23653
rect 8849 23613 8861 23647
rect 8895 23644 8907 23647
rect 9214 23644 9220 23656
rect 8895 23616 9220 23644
rect 8895 23613 8907 23616
rect 8849 23607 8907 23613
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 10594 23604 10600 23656
rect 10652 23604 10658 23656
rect 12345 23647 12403 23653
rect 12345 23613 12357 23647
rect 12391 23613 12403 23647
rect 12345 23607 12403 23613
rect 10318 23576 10324 23588
rect 6564 23548 10324 23576
rect 10318 23536 10324 23548
rect 10376 23536 10382 23588
rect 12360 23576 12388 23607
rect 12618 23604 12624 23656
rect 12676 23604 12682 23656
rect 15841 23647 15899 23653
rect 15841 23613 15853 23647
rect 15887 23644 15899 23647
rect 16390 23644 16396 23656
rect 15887 23616 16396 23644
rect 15887 23613 15899 23616
rect 15841 23607 15899 23613
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18322 23644 18328 23656
rect 17911 23616 18328 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 17218 23576 17224 23588
rect 12360 23548 17224 23576
rect 17218 23536 17224 23548
rect 17276 23536 17282 23588
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 5718 23508 5724 23520
rect 2832 23480 5724 23508
rect 2832 23468 2838 23480
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 5994 23468 6000 23520
rect 6052 23508 6058 23520
rect 6641 23511 6699 23517
rect 6641 23508 6653 23511
rect 6052 23480 6653 23508
rect 6052 23468 6058 23480
rect 6641 23477 6653 23480
rect 6687 23477 6699 23511
rect 6641 23471 6699 23477
rect 18782 23468 18788 23520
rect 18840 23468 18846 23520
rect 19076 23508 19104 23684
rect 21269 23681 21281 23715
rect 21315 23712 21327 23715
rect 21468 23712 21496 23752
rect 22848 23721 22876 23752
rect 23474 23740 23480 23752
rect 23532 23780 23538 23792
rect 24489 23783 24547 23789
rect 24489 23780 24501 23783
rect 23532 23752 24501 23780
rect 23532 23740 23538 23752
rect 24489 23749 24501 23752
rect 24535 23749 24547 23783
rect 24489 23743 24547 23749
rect 25866 23740 25872 23792
rect 25924 23740 25930 23792
rect 26329 23783 26387 23789
rect 26329 23749 26341 23783
rect 26375 23780 26387 23783
rect 27706 23780 27712 23792
rect 26375 23752 27712 23780
rect 26375 23749 26387 23752
rect 26329 23743 26387 23749
rect 27706 23740 27712 23752
rect 27764 23740 27770 23792
rect 21315 23684 21496 23712
rect 22833 23715 22891 23721
rect 21315 23681 21327 23684
rect 21269 23675 21327 23681
rect 22833 23681 22845 23715
rect 22879 23681 22891 23715
rect 22833 23675 22891 23681
rect 23566 23672 23572 23724
rect 23624 23712 23630 23724
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23624 23684 23673 23712
rect 23624 23672 23630 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23712 24455 23715
rect 24946 23712 24952 23724
rect 24443 23684 24952 23712
rect 24443 23681 24455 23684
rect 24397 23675 24455 23681
rect 24946 23672 24952 23684
rect 25004 23672 25010 23724
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 20533 23647 20591 23653
rect 20533 23613 20545 23647
rect 20579 23644 20591 23647
rect 21726 23644 21732 23656
rect 20579 23616 21732 23644
rect 20579 23613 20591 23616
rect 20533 23607 20591 23613
rect 21726 23604 21732 23616
rect 21784 23604 21790 23656
rect 22554 23604 22560 23656
rect 22612 23604 22618 23656
rect 23750 23604 23756 23656
rect 23808 23604 23814 23656
rect 23845 23647 23903 23653
rect 23845 23613 23857 23647
rect 23891 23613 23903 23647
rect 23845 23607 23903 23613
rect 22738 23576 22744 23588
rect 20456 23548 22744 23576
rect 20456 23508 20484 23548
rect 22738 23536 22744 23548
rect 22796 23536 22802 23588
rect 23658 23536 23664 23588
rect 23716 23576 23722 23588
rect 23860 23576 23888 23607
rect 24854 23604 24860 23656
rect 24912 23644 24918 23656
rect 25590 23644 25596 23656
rect 24912 23616 25596 23644
rect 24912 23604 24918 23616
rect 25590 23604 25596 23616
rect 25648 23604 25654 23656
rect 26602 23604 26608 23656
rect 26660 23604 26666 23656
rect 27356 23576 27384 23675
rect 27798 23672 27804 23724
rect 27856 23712 27862 23724
rect 28534 23712 28540 23724
rect 27856 23684 28540 23712
rect 27856 23672 27862 23684
rect 28534 23672 28540 23684
rect 28592 23672 28598 23724
rect 28644 23721 28672 23820
rect 32309 23817 32321 23820
rect 32355 23817 32367 23851
rect 32309 23811 32367 23817
rect 32769 23851 32827 23857
rect 32769 23817 32781 23851
rect 32815 23848 32827 23851
rect 37461 23851 37519 23857
rect 37461 23848 37473 23851
rect 32815 23820 37473 23848
rect 32815 23817 32827 23820
rect 32769 23811 32827 23817
rect 37461 23817 37473 23820
rect 37507 23817 37519 23851
rect 37461 23811 37519 23817
rect 37829 23851 37887 23857
rect 37829 23817 37841 23851
rect 37875 23848 37887 23851
rect 40034 23848 40040 23860
rect 37875 23820 40040 23848
rect 37875 23817 37887 23820
rect 37829 23811 37887 23817
rect 40034 23808 40040 23820
rect 40092 23808 40098 23860
rect 41690 23848 41696 23860
rect 41386 23820 41696 23848
rect 31018 23740 31024 23792
rect 31076 23780 31082 23792
rect 31386 23780 31392 23792
rect 31076 23752 31392 23780
rect 31076 23740 31082 23752
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 31481 23783 31539 23789
rect 31481 23749 31493 23783
rect 31527 23780 31539 23783
rect 32490 23780 32496 23792
rect 31527 23752 32496 23780
rect 31527 23749 31539 23752
rect 31481 23743 31539 23749
rect 32490 23740 32496 23752
rect 32548 23780 32554 23792
rect 33042 23780 33048 23792
rect 32548 23752 33048 23780
rect 32548 23740 32554 23752
rect 33042 23740 33048 23752
rect 33100 23740 33106 23792
rect 35618 23740 35624 23792
rect 35676 23780 35682 23792
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 35676 23752 37933 23780
rect 35676 23740 35682 23752
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 39206 23740 39212 23792
rect 39264 23740 39270 23792
rect 39301 23783 39359 23789
rect 39301 23749 39313 23783
rect 39347 23780 39359 23783
rect 41386 23780 41414 23820
rect 41690 23808 41696 23820
rect 41748 23848 41754 23860
rect 42518 23848 42524 23860
rect 41748 23820 42524 23848
rect 41748 23808 41754 23820
rect 42518 23808 42524 23820
rect 42576 23808 42582 23860
rect 44637 23851 44695 23857
rect 44637 23848 44649 23851
rect 42904 23820 44649 23848
rect 42429 23783 42487 23789
rect 42429 23780 42441 23783
rect 39347 23752 41414 23780
rect 41892 23752 42441 23780
rect 39347 23749 39359 23752
rect 39301 23743 39359 23749
rect 28629 23715 28687 23721
rect 28629 23681 28641 23715
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 29089 23715 29147 23721
rect 29089 23681 29101 23715
rect 29135 23712 29147 23715
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 29135 23684 29561 23712
rect 29135 23681 29147 23684
rect 29089 23675 29147 23681
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 28442 23604 28448 23656
rect 28500 23644 28506 23656
rect 29104 23644 29132 23675
rect 32674 23672 32680 23724
rect 32732 23672 32738 23724
rect 32766 23672 32772 23724
rect 32824 23712 32830 23724
rect 36265 23715 36323 23721
rect 32824 23684 33994 23712
rect 32824 23672 32830 23684
rect 36265 23681 36277 23715
rect 36311 23712 36323 23715
rect 36311 23684 38148 23712
rect 36311 23681 36323 23684
rect 36265 23675 36323 23681
rect 28500 23616 29132 23644
rect 28500 23604 28506 23616
rect 29178 23604 29184 23656
rect 29236 23644 29242 23656
rect 31018 23644 31024 23656
rect 29236 23616 31024 23644
rect 29236 23604 29242 23616
rect 31018 23604 31024 23616
rect 31076 23604 31082 23656
rect 31754 23604 31760 23656
rect 31812 23604 31818 23656
rect 32953 23647 33011 23653
rect 32953 23613 32965 23647
rect 32999 23644 33011 23647
rect 32999 23616 33640 23644
rect 32999 23613 33011 23616
rect 32953 23607 33011 23613
rect 29730 23576 29736 23588
rect 23716 23548 23888 23576
rect 23952 23548 24992 23576
rect 27356 23548 29736 23576
rect 23716 23536 23722 23548
rect 19076 23480 20484 23508
rect 20806 23468 20812 23520
rect 20864 23508 20870 23520
rect 20901 23511 20959 23517
rect 20901 23508 20913 23511
rect 20864 23480 20913 23508
rect 20864 23468 20870 23480
rect 20901 23477 20913 23480
rect 20947 23477 20959 23511
rect 20901 23471 20959 23477
rect 20990 23468 20996 23520
rect 21048 23508 21054 23520
rect 23293 23511 23351 23517
rect 23293 23508 23305 23511
rect 21048 23480 23305 23508
rect 21048 23468 21054 23480
rect 23293 23477 23305 23480
rect 23339 23477 23351 23511
rect 23293 23471 23351 23477
rect 23842 23468 23848 23520
rect 23900 23508 23906 23520
rect 23952 23508 23980 23548
rect 23900 23480 23980 23508
rect 23900 23468 23906 23480
rect 24854 23468 24860 23520
rect 24912 23468 24918 23520
rect 24964 23508 24992 23548
rect 29730 23536 29736 23548
rect 29788 23536 29794 23588
rect 29822 23536 29828 23588
rect 29880 23576 29886 23588
rect 29880 23548 30420 23576
rect 29880 23536 29886 23548
rect 27157 23511 27215 23517
rect 27157 23508 27169 23511
rect 24964 23480 27169 23508
rect 27157 23477 27169 23480
rect 27203 23477 27215 23511
rect 27157 23471 27215 23477
rect 27798 23468 27804 23520
rect 27856 23508 27862 23520
rect 27985 23511 28043 23517
rect 27985 23508 27997 23511
rect 27856 23480 27997 23508
rect 27856 23468 27862 23480
rect 27985 23477 27997 23480
rect 28031 23477 28043 23511
rect 27985 23471 28043 23477
rect 29270 23468 29276 23520
rect 29328 23468 29334 23520
rect 30009 23511 30067 23517
rect 30009 23477 30021 23511
rect 30055 23508 30067 23511
rect 30282 23508 30288 23520
rect 30055 23480 30288 23508
rect 30055 23477 30067 23480
rect 30009 23471 30067 23477
rect 30282 23468 30288 23480
rect 30340 23468 30346 23520
rect 30392 23508 30420 23548
rect 32306 23508 32312 23520
rect 30392 23480 32312 23508
rect 32306 23468 32312 23480
rect 32364 23468 32370 23520
rect 33612 23517 33640 23616
rect 34974 23604 34980 23656
rect 35032 23644 35038 23656
rect 35345 23647 35403 23653
rect 35345 23644 35357 23647
rect 35032 23616 35357 23644
rect 35032 23604 35038 23616
rect 35345 23613 35357 23616
rect 35391 23644 35403 23647
rect 35391 23616 36124 23644
rect 35391 23613 35403 23616
rect 35345 23607 35403 23613
rect 35894 23536 35900 23588
rect 35952 23536 35958 23588
rect 36096 23576 36124 23616
rect 36170 23604 36176 23656
rect 36228 23644 36234 23656
rect 36357 23647 36415 23653
rect 36357 23644 36369 23647
rect 36228 23616 36369 23644
rect 36228 23604 36234 23616
rect 36357 23613 36369 23616
rect 36403 23613 36415 23647
rect 36357 23607 36415 23613
rect 36446 23604 36452 23656
rect 36504 23604 36510 23656
rect 36538 23604 36544 23656
rect 36596 23644 36602 23656
rect 38013 23647 38071 23653
rect 38013 23644 38025 23647
rect 36596 23616 38025 23644
rect 36596 23604 36602 23616
rect 38013 23613 38025 23616
rect 38059 23613 38071 23647
rect 38120 23644 38148 23684
rect 38838 23672 38844 23724
rect 38896 23712 38902 23724
rect 41892 23712 41920 23752
rect 42429 23749 42441 23752
rect 42475 23749 42487 23783
rect 42904 23780 42932 23820
rect 44637 23817 44649 23820
rect 44683 23817 44695 23851
rect 44637 23811 44695 23817
rect 47302 23808 47308 23860
rect 47360 23848 47366 23860
rect 47581 23851 47639 23857
rect 47581 23848 47593 23851
rect 47360 23820 47593 23848
rect 47360 23808 47366 23820
rect 47581 23817 47593 23820
rect 47627 23817 47639 23851
rect 47581 23811 47639 23817
rect 49142 23808 49148 23860
rect 49200 23808 49206 23860
rect 49510 23808 49516 23860
rect 49568 23808 49574 23860
rect 42429 23743 42487 23749
rect 42628 23752 42932 23780
rect 38896 23684 41920 23712
rect 42061 23715 42119 23721
rect 38896 23672 38902 23684
rect 42061 23681 42073 23715
rect 42107 23712 42119 23715
rect 42628 23712 42656 23752
rect 42978 23740 42984 23792
rect 43036 23780 43042 23792
rect 43349 23783 43407 23789
rect 43349 23780 43361 23783
rect 43036 23752 43361 23780
rect 43036 23740 43042 23752
rect 43349 23749 43361 23752
rect 43395 23749 43407 23783
rect 43349 23743 43407 23749
rect 44192 23752 46888 23780
rect 44192 23721 44220 23752
rect 46860 23724 46888 23752
rect 42107 23684 42656 23712
rect 44177 23715 44235 23721
rect 42107 23681 42119 23684
rect 42061 23675 42119 23681
rect 44177 23681 44189 23715
rect 44223 23681 44235 23715
rect 44177 23675 44235 23681
rect 44818 23672 44824 23724
rect 44876 23672 44882 23724
rect 45925 23715 45983 23721
rect 45925 23681 45937 23715
rect 45971 23681 45983 23715
rect 45925 23675 45983 23681
rect 39393 23647 39451 23653
rect 38120 23616 38884 23644
rect 38013 23607 38071 23613
rect 38856 23585 38884 23616
rect 39393 23613 39405 23647
rect 39439 23613 39451 23647
rect 39393 23607 39451 23613
rect 36909 23579 36967 23585
rect 36909 23576 36921 23579
rect 36096 23548 36921 23576
rect 36909 23545 36921 23548
rect 36955 23545 36967 23579
rect 36909 23539 36967 23545
rect 38841 23579 38899 23585
rect 38841 23545 38853 23579
rect 38887 23545 38899 23579
rect 38841 23539 38899 23545
rect 33597 23511 33655 23517
rect 33597 23477 33609 23511
rect 33643 23508 33655 23511
rect 34514 23508 34520 23520
rect 33643 23480 34520 23508
rect 33643 23477 33655 23480
rect 33597 23471 33655 23477
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 35087 23511 35145 23517
rect 35087 23477 35099 23511
rect 35133 23508 35145 23511
rect 35434 23508 35440 23520
rect 35133 23480 35440 23508
rect 35133 23477 35145 23480
rect 35087 23471 35145 23477
rect 35434 23468 35440 23480
rect 35492 23508 35498 23520
rect 36538 23508 36544 23520
rect 35492 23480 36544 23508
rect 35492 23468 35498 23480
rect 36538 23468 36544 23480
rect 36596 23468 36602 23520
rect 36924 23508 36952 23539
rect 39408 23520 39436 23607
rect 39758 23604 39764 23656
rect 39816 23644 39822 23656
rect 39945 23647 40003 23653
rect 39945 23644 39957 23647
rect 39816 23616 39957 23644
rect 39816 23604 39822 23616
rect 39945 23613 39957 23616
rect 39991 23644 40003 23647
rect 40313 23647 40371 23653
rect 40313 23644 40325 23647
rect 39991 23616 40325 23644
rect 39991 23613 40003 23616
rect 39945 23607 40003 23613
rect 40313 23613 40325 23616
rect 40359 23644 40371 23647
rect 41046 23644 41052 23656
rect 40359 23616 41052 23644
rect 40359 23613 40371 23616
rect 40313 23607 40371 23613
rect 41046 23604 41052 23616
rect 41104 23604 41110 23656
rect 43165 23647 43223 23653
rect 43165 23644 43177 23647
rect 41156 23616 43177 23644
rect 39482 23536 39488 23588
rect 39540 23576 39546 23588
rect 41156 23576 41184 23616
rect 43165 23613 43177 23616
rect 43211 23613 43223 23647
rect 45940 23644 45968 23675
rect 46382 23672 46388 23724
rect 46440 23672 46446 23724
rect 46842 23672 46848 23724
rect 46900 23712 46906 23724
rect 47305 23715 47363 23721
rect 47305 23712 47317 23715
rect 46900 23684 47317 23712
rect 46900 23672 46906 23684
rect 47305 23681 47317 23684
rect 47351 23681 47363 23715
rect 47305 23675 47363 23681
rect 48222 23672 48228 23724
rect 48280 23712 48286 23724
rect 48777 23715 48835 23721
rect 48777 23712 48789 23715
rect 48280 23684 48789 23712
rect 48280 23672 48286 23684
rect 48777 23681 48789 23684
rect 48823 23681 48835 23715
rect 48777 23675 48835 23681
rect 47029 23647 47087 23653
rect 47029 23644 47041 23647
rect 45940 23616 47041 23644
rect 43165 23607 43223 23613
rect 47029 23613 47041 23616
rect 47075 23613 47087 23647
rect 47029 23607 47087 23613
rect 41506 23576 41512 23588
rect 39540 23548 41184 23576
rect 41386 23548 41512 23576
rect 39540 23536 39546 23548
rect 38562 23508 38568 23520
rect 36924 23480 38568 23508
rect 38562 23468 38568 23480
rect 38620 23468 38626 23520
rect 39390 23468 39396 23520
rect 39448 23508 39454 23520
rect 41386 23508 41414 23548
rect 41506 23536 41512 23548
rect 41564 23576 41570 23588
rect 42981 23579 43039 23585
rect 42981 23576 42993 23579
rect 41564 23548 42993 23576
rect 41564 23536 41570 23548
rect 42981 23545 42993 23548
rect 43027 23545 43039 23579
rect 42981 23539 43039 23545
rect 43530 23536 43536 23588
rect 43588 23536 43594 23588
rect 43990 23536 43996 23588
rect 44048 23536 44054 23588
rect 46014 23536 46020 23588
rect 46072 23576 46078 23588
rect 48133 23579 48191 23585
rect 48133 23576 48145 23579
rect 46072 23548 48145 23576
rect 46072 23536 46078 23548
rect 48133 23545 48145 23548
rect 48179 23545 48191 23579
rect 48133 23539 48191 23545
rect 39448 23480 41414 23508
rect 39448 23468 39454 23480
rect 42426 23468 42432 23520
rect 42484 23508 42490 23520
rect 42613 23511 42671 23517
rect 42613 23508 42625 23511
rect 42484 23480 42625 23508
rect 42484 23468 42490 23480
rect 42613 23477 42625 23480
rect 42659 23477 42671 23511
rect 42613 23471 42671 23477
rect 42886 23468 42892 23520
rect 42944 23508 42950 23520
rect 43622 23508 43628 23520
rect 42944 23480 43628 23508
rect 42944 23468 42950 23480
rect 43622 23468 43628 23480
rect 43680 23468 43686 23520
rect 44726 23468 44732 23520
rect 44784 23508 44790 23520
rect 45281 23511 45339 23517
rect 45281 23508 45293 23511
rect 44784 23480 45293 23508
rect 44784 23468 44790 23480
rect 45281 23477 45293 23480
rect 45327 23477 45339 23511
rect 45281 23471 45339 23477
rect 47857 23511 47915 23517
rect 47857 23477 47869 23511
rect 47903 23508 47915 23511
rect 48038 23508 48044 23520
rect 47903 23480 48044 23508
rect 47903 23477 47915 23480
rect 47857 23471 47915 23477
rect 48038 23468 48044 23480
rect 48096 23468 48102 23520
rect 49326 23468 49332 23520
rect 49384 23468 49390 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 4706 23264 4712 23316
rect 4764 23264 4770 23316
rect 23658 23304 23664 23316
rect 20364 23276 23664 23304
rect 20364 23248 20392 23276
rect 23658 23264 23664 23276
rect 23716 23264 23722 23316
rect 23750 23264 23756 23316
rect 23808 23304 23814 23316
rect 27893 23307 27951 23313
rect 27893 23304 27905 23307
rect 23808 23276 27905 23304
rect 23808 23264 23814 23276
rect 27893 23273 27905 23276
rect 27939 23273 27951 23307
rect 27893 23267 27951 23273
rect 28534 23264 28540 23316
rect 28592 23304 28598 23316
rect 28997 23307 29055 23313
rect 28997 23304 29009 23307
rect 28592 23276 29009 23304
rect 28592 23264 28598 23276
rect 28997 23273 29009 23276
rect 29043 23273 29055 23307
rect 28997 23267 29055 23273
rect 29178 23264 29184 23316
rect 29236 23264 29242 23316
rect 29730 23264 29736 23316
rect 29788 23264 29794 23316
rect 29914 23264 29920 23316
rect 29972 23304 29978 23316
rect 33318 23304 33324 23316
rect 29972 23276 33324 23304
rect 29972 23264 29978 23276
rect 33318 23264 33324 23276
rect 33376 23304 33382 23316
rect 34149 23307 34207 23313
rect 34149 23304 34161 23307
rect 33376 23276 34161 23304
rect 33376 23264 33382 23276
rect 34149 23273 34161 23276
rect 34195 23273 34207 23307
rect 34149 23267 34207 23273
rect 35066 23264 35072 23316
rect 35124 23304 35130 23316
rect 36630 23304 36636 23316
rect 35124 23276 36636 23304
rect 35124 23264 35130 23276
rect 36630 23264 36636 23276
rect 36688 23264 36694 23316
rect 39022 23304 39028 23316
rect 37292 23276 39028 23304
rect 5626 23236 5632 23248
rect 4172 23208 5632 23236
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23100 3019 23103
rect 4172 23100 4200 23208
rect 5626 23196 5632 23208
rect 5684 23196 5690 23248
rect 15838 23236 15844 23248
rect 10060 23208 15844 23236
rect 4908 23140 6040 23168
rect 3007 23072 4200 23100
rect 4249 23103 4307 23109
rect 3007 23069 3019 23072
rect 2961 23063 3019 23069
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4430 23100 4436 23112
rect 4295 23072 4436 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4430 23060 4436 23072
rect 4488 23060 4494 23112
rect 4908 23109 4936 23140
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 1762 22992 1768 23044
rect 1820 22992 1826 23044
rect 3602 22992 3608 23044
rect 3660 23032 3666 23044
rect 5368 23032 5396 23063
rect 3660 23004 5396 23032
rect 6012 23032 6040 23140
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 10060 23177 10088 23208
rect 15838 23196 15844 23208
rect 15896 23196 15902 23248
rect 19610 23196 19616 23248
rect 19668 23196 19674 23248
rect 20346 23196 20352 23248
rect 20404 23196 20410 23248
rect 22738 23196 22744 23248
rect 22796 23236 22802 23248
rect 24581 23239 24639 23245
rect 24581 23236 24593 23239
rect 22796 23208 24593 23236
rect 22796 23196 22802 23208
rect 24581 23205 24593 23208
rect 24627 23205 24639 23239
rect 24581 23199 24639 23205
rect 25225 23239 25283 23245
rect 25225 23205 25237 23239
rect 25271 23236 25283 23239
rect 25406 23236 25412 23248
rect 25271 23208 25412 23236
rect 25271 23205 25283 23208
rect 25225 23199 25283 23205
rect 25406 23196 25412 23208
rect 25464 23196 25470 23248
rect 31294 23236 31300 23248
rect 30116 23208 31300 23236
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23137 10103 23171
rect 10045 23131 10103 23137
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13354 23168 13360 23180
rect 13311 23140 13360 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 15746 23128 15752 23180
rect 15804 23128 15810 23180
rect 17586 23168 17592 23180
rect 16224 23140 17592 23168
rect 6638 23060 6644 23112
rect 6696 23100 6702 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 6696 23072 7205 23100
rect 6696 23060 6702 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 9122 23060 9128 23112
rect 9180 23100 9186 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 9180 23072 9321 23100
rect 9180 23060 9186 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 11882 23060 11888 23112
rect 11940 23060 11946 23112
rect 13725 23103 13783 23109
rect 13725 23069 13737 23103
rect 13771 23100 13783 23103
rect 13906 23100 13912 23112
rect 13771 23072 13912 23100
rect 13771 23069 13783 23072
rect 13725 23063 13783 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23100 14887 23103
rect 16224 23100 16252 23140
rect 17586 23128 17592 23140
rect 17644 23128 17650 23180
rect 18230 23128 18236 23180
rect 18288 23168 18294 23180
rect 18601 23171 18659 23177
rect 18601 23168 18613 23171
rect 18288 23140 18613 23168
rect 18288 23128 18294 23140
rect 18601 23137 18613 23140
rect 18647 23168 18659 23171
rect 19058 23168 19064 23180
rect 18647 23140 19064 23168
rect 18647 23137 18659 23140
rect 18601 23131 18659 23137
rect 19058 23128 19064 23140
rect 19116 23128 19122 23180
rect 19242 23128 19248 23180
rect 19300 23168 19306 23180
rect 19337 23171 19395 23177
rect 19337 23168 19349 23171
rect 19300 23140 19349 23168
rect 19300 23128 19306 23140
rect 19337 23137 19349 23140
rect 19383 23168 19395 23171
rect 20806 23168 20812 23180
rect 19383 23140 20812 23168
rect 19383 23137 19395 23140
rect 19337 23131 19395 23137
rect 20806 23128 20812 23140
rect 20864 23128 20870 23180
rect 21726 23128 21732 23180
rect 21784 23168 21790 23180
rect 22097 23171 22155 23177
rect 22097 23168 22109 23171
rect 21784 23140 22109 23168
rect 21784 23128 21790 23140
rect 22097 23137 22109 23140
rect 22143 23137 22155 23171
rect 22097 23131 22155 23137
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 24854 23168 24860 23180
rect 23983 23140 24860 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 24854 23128 24860 23140
rect 24912 23168 24918 23180
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 24912 23140 25973 23168
rect 24912 23128 24918 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 25961 23131 26019 23137
rect 26326 23128 26332 23180
rect 26384 23168 26390 23180
rect 28445 23171 28503 23177
rect 28445 23168 28457 23171
rect 26384 23140 28457 23168
rect 26384 23128 26390 23140
rect 28445 23137 28457 23140
rect 28491 23137 28503 23171
rect 28445 23131 28503 23137
rect 14875 23072 16252 23100
rect 16669 23103 16727 23109
rect 14875 23069 14887 23072
rect 14829 23063 14887 23069
rect 16669 23069 16681 23103
rect 16715 23100 16727 23103
rect 16715 23072 17356 23100
rect 16715 23069 16727 23072
rect 16669 23063 16727 23069
rect 7834 23032 7840 23044
rect 6012 23004 7840 23032
rect 3660 22992 3666 23004
rect 7834 22992 7840 23004
rect 7892 22992 7898 23044
rect 4065 22967 4123 22973
rect 4065 22933 4077 22967
rect 4111 22964 4123 22967
rect 4614 22964 4620 22976
rect 4111 22936 4620 22964
rect 4111 22933 4123 22936
rect 4065 22927 4123 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 5442 22924 5448 22976
rect 5500 22964 5506 22976
rect 9217 22967 9275 22973
rect 9217 22964 9229 22967
rect 5500 22936 9229 22964
rect 5500 22924 5506 22936
rect 9217 22933 9229 22936
rect 9263 22933 9275 22967
rect 9217 22927 9275 22933
rect 14182 22924 14188 22976
rect 14240 22924 14246 22976
rect 14366 22924 14372 22976
rect 14424 22924 14430 22976
rect 14642 22924 14648 22976
rect 14700 22924 14706 22976
rect 17129 22967 17187 22973
rect 17129 22933 17141 22967
rect 17175 22964 17187 22967
rect 17218 22964 17224 22976
rect 17175 22936 17224 22964
rect 17175 22933 17187 22936
rect 17129 22927 17187 22933
rect 17218 22924 17224 22936
rect 17276 22924 17282 22976
rect 17328 22964 17356 23072
rect 18874 23060 18880 23112
rect 18932 23060 18938 23112
rect 23753 23103 23811 23109
rect 23753 23069 23765 23103
rect 23799 23100 23811 23103
rect 23799 23072 25636 23100
rect 23799 23069 23811 23072
rect 23753 23063 23811 23069
rect 18506 23032 18512 23044
rect 18170 23004 18512 23032
rect 18506 22992 18512 23004
rect 18564 22992 18570 23044
rect 19518 23032 19524 23044
rect 18708 23004 19524 23032
rect 18708 22964 18736 23004
rect 19518 22992 19524 23004
rect 19576 22992 19582 23044
rect 19794 22992 19800 23044
rect 19852 22992 19858 23044
rect 21542 23032 21548 23044
rect 21390 23004 21548 23032
rect 21542 22992 21548 23004
rect 21600 22992 21606 23044
rect 21818 22992 21824 23044
rect 21876 22992 21882 23044
rect 21910 22992 21916 23044
rect 21968 23032 21974 23044
rect 22557 23035 22615 23041
rect 22557 23032 22569 23035
rect 21968 23004 22569 23032
rect 21968 22992 21974 23004
rect 22557 23001 22569 23004
rect 22603 23001 22615 23035
rect 22557 22995 22615 23001
rect 22741 23035 22799 23041
rect 22741 23001 22753 23035
rect 22787 23032 22799 23035
rect 24670 23032 24676 23044
rect 22787 23004 24676 23032
rect 22787 23001 22799 23004
rect 22741 22995 22799 23001
rect 24670 22992 24676 23004
rect 24728 22992 24734 23044
rect 24762 22992 24768 23044
rect 24820 22992 24826 23044
rect 17328 22936 18736 22964
rect 18782 22924 18788 22976
rect 18840 22964 18846 22976
rect 22002 22964 22008 22976
rect 18840 22936 22008 22964
rect 18840 22924 18846 22936
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 23290 22924 23296 22976
rect 23348 22924 23354 22976
rect 23658 22924 23664 22976
rect 23716 22924 23722 22976
rect 25314 22924 25320 22976
rect 25372 22924 25378 22976
rect 25608 22964 25636 23072
rect 25682 23060 25688 23112
rect 25740 23060 25746 23112
rect 28261 23103 28319 23109
rect 28261 23069 28273 23103
rect 28307 23100 28319 23103
rect 30116 23100 30144 23208
rect 31294 23196 31300 23208
rect 31352 23196 31358 23248
rect 32858 23196 32864 23248
rect 32916 23236 32922 23248
rect 34333 23239 34391 23245
rect 34333 23236 34345 23239
rect 32916 23208 34345 23236
rect 32916 23196 32922 23208
rect 34333 23205 34345 23208
rect 34379 23205 34391 23239
rect 34333 23199 34391 23205
rect 30190 23128 30196 23180
rect 30248 23128 30254 23180
rect 30282 23128 30288 23180
rect 30340 23128 30346 23180
rect 30837 23171 30895 23177
rect 30837 23137 30849 23171
rect 30883 23168 30895 23171
rect 31018 23168 31024 23180
rect 30883 23140 31024 23168
rect 30883 23137 30895 23140
rect 30837 23131 30895 23137
rect 31018 23128 31024 23140
rect 31076 23128 31082 23180
rect 31389 23171 31447 23177
rect 31389 23137 31401 23171
rect 31435 23168 31447 23171
rect 31662 23168 31668 23180
rect 31435 23140 31668 23168
rect 31435 23137 31447 23140
rect 31389 23131 31447 23137
rect 31662 23128 31668 23140
rect 31720 23168 31726 23180
rect 31754 23168 31760 23180
rect 31720 23140 31760 23168
rect 31720 23128 31726 23140
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 33137 23171 33195 23177
rect 33137 23137 33149 23171
rect 33183 23168 33195 23171
rect 33318 23168 33324 23180
rect 33183 23140 33324 23168
rect 33183 23137 33195 23140
rect 33137 23131 33195 23137
rect 33318 23128 33324 23140
rect 33376 23168 33382 23180
rect 33778 23168 33784 23180
rect 33376 23140 33784 23168
rect 33376 23128 33382 23140
rect 33778 23128 33784 23140
rect 33836 23128 33842 23180
rect 34514 23128 34520 23180
rect 34572 23168 34578 23180
rect 35345 23171 35403 23177
rect 35345 23168 35357 23171
rect 34572 23140 35357 23168
rect 34572 23128 34578 23140
rect 35345 23137 35357 23140
rect 35391 23137 35403 23171
rect 35345 23131 35403 23137
rect 35710 23128 35716 23180
rect 35768 23168 35774 23180
rect 37292 23177 37320 23276
rect 39022 23264 39028 23276
rect 39080 23264 39086 23316
rect 39298 23264 39304 23316
rect 39356 23304 39362 23316
rect 39356 23276 41552 23304
rect 39356 23264 39362 23276
rect 41524 23236 41552 23276
rect 41598 23264 41604 23316
rect 41656 23304 41662 23316
rect 43530 23304 43536 23316
rect 41656 23276 43536 23304
rect 41656 23264 41662 23276
rect 43530 23264 43536 23276
rect 43588 23264 43594 23316
rect 43622 23264 43628 23316
rect 43680 23304 43686 23316
rect 44542 23304 44548 23316
rect 43680 23276 44548 23304
rect 43680 23264 43686 23276
rect 44542 23264 44548 23276
rect 44600 23264 44606 23316
rect 44637 23307 44695 23313
rect 44637 23273 44649 23307
rect 44683 23304 44695 23307
rect 44818 23304 44824 23316
rect 44683 23276 44824 23304
rect 44683 23273 44695 23276
rect 44637 23267 44695 23273
rect 44818 23264 44824 23276
rect 44876 23264 44882 23316
rect 48222 23264 48228 23316
rect 48280 23264 48286 23316
rect 42242 23236 42248 23248
rect 39500 23208 41414 23236
rect 41524 23208 42248 23236
rect 37277 23171 37335 23177
rect 37277 23168 37289 23171
rect 35768 23140 37289 23168
rect 35768 23128 35774 23140
rect 37277 23137 37289 23140
rect 37323 23137 37335 23171
rect 37277 23131 37335 23137
rect 38654 23128 38660 23180
rect 38712 23168 38718 23180
rect 39025 23171 39083 23177
rect 39025 23168 39037 23171
rect 38712 23140 39037 23168
rect 38712 23128 38718 23140
rect 39025 23137 39037 23140
rect 39071 23168 39083 23171
rect 39206 23168 39212 23180
rect 39071 23140 39212 23168
rect 39071 23137 39083 23140
rect 39025 23131 39083 23137
rect 39206 23128 39212 23140
rect 39264 23168 39270 23180
rect 39500 23177 39528 23208
rect 39485 23171 39543 23177
rect 39485 23168 39497 23171
rect 39264 23140 39497 23168
rect 39264 23128 39270 23140
rect 39485 23137 39497 23140
rect 39531 23137 39543 23171
rect 39485 23131 39543 23137
rect 40589 23171 40647 23177
rect 40589 23137 40601 23171
rect 40635 23137 40647 23171
rect 40589 23131 40647 23137
rect 28307 23072 30144 23100
rect 28307 23069 28319 23072
rect 28261 23063 28319 23069
rect 27246 23032 27252 23044
rect 27186 23004 27252 23032
rect 27246 22992 27252 23004
rect 27304 22992 27310 23044
rect 27614 23032 27620 23044
rect 27356 23004 27620 23032
rect 27356 22964 27384 23004
rect 27614 22992 27620 23004
rect 27672 22992 27678 23044
rect 28353 23035 28411 23041
rect 28353 23001 28365 23035
rect 28399 23032 28411 23035
rect 30300 23032 30328 23128
rect 32766 23060 32772 23112
rect 32824 23060 32830 23112
rect 33873 23103 33931 23109
rect 33873 23100 33885 23103
rect 33060 23072 33885 23100
rect 31665 23035 31723 23041
rect 31665 23032 31677 23035
rect 28399 23004 29408 23032
rect 30300 23004 31677 23032
rect 28399 23001 28411 23004
rect 28353 22995 28411 23001
rect 29380 22976 29408 23004
rect 31665 23001 31677 23004
rect 31711 23001 31723 23035
rect 31665 22995 31723 23001
rect 25608 22936 27384 22964
rect 27430 22924 27436 22976
rect 27488 22924 27494 22976
rect 29362 22924 29368 22976
rect 29420 22924 29426 22976
rect 30098 22924 30104 22976
rect 30156 22924 30162 22976
rect 30742 22924 30748 22976
rect 30800 22964 30806 22976
rect 31021 22967 31079 22973
rect 31021 22964 31033 22967
rect 30800 22936 31033 22964
rect 30800 22924 30806 22936
rect 31021 22933 31033 22936
rect 31067 22933 31079 22967
rect 31021 22927 31079 22933
rect 31202 22924 31208 22976
rect 31260 22964 31266 22976
rect 33060 22964 33088 23072
rect 33873 23069 33885 23072
rect 33919 23100 33931 23103
rect 34238 23100 34244 23112
rect 33919 23072 34244 23100
rect 33919 23069 33931 23072
rect 33873 23063 33931 23069
rect 34238 23060 34244 23072
rect 34296 23060 34302 23112
rect 34974 23060 34980 23112
rect 35032 23100 35038 23112
rect 35069 23103 35127 23109
rect 35069 23100 35081 23103
rect 35032 23072 35081 23100
rect 35032 23060 35038 23072
rect 35069 23069 35081 23072
rect 35115 23069 35127 23103
rect 37366 23100 37372 23112
rect 35069 23063 35127 23069
rect 36648 23072 37372 23100
rect 33226 22992 33232 23044
rect 33284 23032 33290 23044
rect 33284 23004 33916 23032
rect 33284 22992 33290 23004
rect 31260 22936 33088 22964
rect 33689 22967 33747 22973
rect 31260 22924 31266 22936
rect 33689 22933 33701 22967
rect 33735 22964 33747 22967
rect 33778 22964 33784 22976
rect 33735 22936 33784 22964
rect 33735 22933 33747 22936
rect 33689 22927 33747 22933
rect 33778 22924 33784 22936
rect 33836 22924 33842 22976
rect 33888 22964 33916 23004
rect 34330 22992 34336 23044
rect 34388 23032 34394 23044
rect 35618 23032 35624 23044
rect 34388 23004 35624 23032
rect 34388 22992 34394 23004
rect 35618 22992 35624 23004
rect 35676 22992 35682 23044
rect 35986 22992 35992 23044
rect 36044 22992 36050 23044
rect 34514 22964 34520 22976
rect 33888 22936 34520 22964
rect 34514 22924 34520 22936
rect 34572 22924 34578 22976
rect 34606 22924 34612 22976
rect 34664 22964 34670 22976
rect 34701 22967 34759 22973
rect 34701 22964 34713 22967
rect 34664 22936 34713 22964
rect 34664 22924 34670 22936
rect 34701 22933 34713 22936
rect 34747 22933 34759 22967
rect 34701 22927 34759 22933
rect 34790 22924 34796 22976
rect 34848 22964 34854 22976
rect 36648 22964 36676 23072
rect 37366 23060 37372 23072
rect 37424 23060 37430 23112
rect 40604 23100 40632 23131
rect 41046 23128 41052 23180
rect 41104 23128 41110 23180
rect 41386 23168 41414 23208
rect 42242 23196 42248 23208
rect 42300 23196 42306 23248
rect 44266 23196 44272 23248
rect 44324 23236 44330 23248
rect 45925 23239 45983 23245
rect 45925 23236 45937 23239
rect 44324 23208 45937 23236
rect 44324 23196 44330 23208
rect 45925 23205 45937 23208
rect 45971 23205 45983 23239
rect 45925 23199 45983 23205
rect 47026 23196 47032 23248
rect 47084 23236 47090 23248
rect 48590 23236 48596 23248
rect 47084 23208 48596 23236
rect 47084 23196 47090 23208
rect 48590 23196 48596 23208
rect 48648 23196 48654 23248
rect 43533 23171 43591 23177
rect 43533 23168 43545 23171
rect 41386 23140 43545 23168
rect 43533 23137 43545 23140
rect 43579 23168 43591 23171
rect 45741 23171 45799 23177
rect 45741 23168 45753 23171
rect 43579 23140 45753 23168
rect 43579 23137 43591 23140
rect 43533 23131 43591 23137
rect 45741 23137 45753 23140
rect 45787 23137 45799 23171
rect 48038 23168 48044 23180
rect 45741 23131 45799 23137
rect 47136 23140 48044 23168
rect 39040 23072 40632 23100
rect 36998 22992 37004 23044
rect 37056 23032 37062 23044
rect 37056 23004 37582 23032
rect 37056 22992 37062 23004
rect 34848 22936 36676 22964
rect 36817 22967 36875 22973
rect 34848 22924 34854 22936
rect 36817 22933 36829 22967
rect 36863 22964 36875 22967
rect 36906 22964 36912 22976
rect 36863 22936 36912 22964
rect 36863 22933 36875 22936
rect 36817 22927 36875 22933
rect 36906 22924 36912 22936
rect 36964 22924 36970 22976
rect 37476 22964 37504 23004
rect 38654 22992 38660 23044
rect 38712 23032 38718 23044
rect 38749 23035 38807 23041
rect 38749 23032 38761 23035
rect 38712 23004 38761 23032
rect 38712 22992 38718 23004
rect 38749 23001 38761 23004
rect 38795 23032 38807 23035
rect 39040 23032 39068 23072
rect 41506 23060 41512 23112
rect 41564 23060 41570 23112
rect 42150 23060 42156 23112
rect 42208 23060 42214 23112
rect 43993 23103 44051 23109
rect 43993 23069 44005 23103
rect 44039 23100 44051 23103
rect 44174 23100 44180 23112
rect 44039 23072 44180 23100
rect 44039 23069 44051 23072
rect 43993 23063 44051 23069
rect 44174 23060 44180 23072
rect 44232 23060 44238 23112
rect 44542 23060 44548 23112
rect 44600 23100 44606 23112
rect 45189 23103 45247 23109
rect 45189 23100 45201 23103
rect 44600 23072 45201 23100
rect 44600 23060 44606 23072
rect 45189 23069 45201 23072
rect 45235 23069 45247 23103
rect 45189 23063 45247 23069
rect 45370 23060 45376 23112
rect 45428 23060 45434 23112
rect 47136 23109 47164 23140
rect 48038 23128 48044 23140
rect 48096 23128 48102 23180
rect 47121 23103 47179 23109
rect 47121 23069 47133 23103
rect 47167 23069 47179 23103
rect 47121 23063 47179 23069
rect 47578 23060 47584 23112
rect 47636 23060 47642 23112
rect 49326 23060 49332 23112
rect 49384 23060 49390 23112
rect 38795 23004 39068 23032
rect 40405 23035 40463 23041
rect 38795 23001 38807 23004
rect 38749 22995 38807 23001
rect 40405 23001 40417 23035
rect 40451 23032 40463 23035
rect 41230 23032 41236 23044
rect 40451 23004 41236 23032
rect 40451 23001 40463 23004
rect 40405 22995 40463 23001
rect 41230 22992 41236 23004
rect 41288 22992 41294 23044
rect 39758 22964 39764 22976
rect 37476 22936 39764 22964
rect 39758 22924 39764 22936
rect 39816 22924 39822 22976
rect 39942 22924 39948 22976
rect 40000 22964 40006 22976
rect 40037 22967 40095 22973
rect 40037 22964 40049 22967
rect 40000 22936 40049 22964
rect 40000 22924 40006 22936
rect 40037 22933 40049 22936
rect 40083 22933 40095 22967
rect 40037 22927 40095 22933
rect 40494 22924 40500 22976
rect 40552 22924 40558 22976
rect 41046 22924 41052 22976
rect 41104 22964 41110 22976
rect 42168 22964 42196 23060
rect 43257 23035 43315 23041
rect 43257 23001 43269 23035
rect 43303 23032 43315 23035
rect 44726 23032 44732 23044
rect 43303 23004 44732 23032
rect 43303 23001 43315 23004
rect 43257 22995 43315 23001
rect 44726 22992 44732 23004
rect 44784 22992 44790 23044
rect 46109 23035 46167 23041
rect 46109 23032 46121 23035
rect 44836 23004 46121 23032
rect 41104 22936 42196 22964
rect 41104 22924 41110 22936
rect 43346 22924 43352 22976
rect 43404 22964 43410 22976
rect 44836 22964 44864 23004
rect 46109 23001 46121 23004
rect 46155 23001 46167 23035
rect 46109 22995 46167 23001
rect 43404 22936 44864 22964
rect 46477 22967 46535 22973
rect 43404 22924 43410 22936
rect 46477 22933 46489 22967
rect 46523 22964 46535 22967
rect 46750 22964 46756 22976
rect 46523 22936 46756 22964
rect 46523 22933 46535 22936
rect 46477 22927 46535 22933
rect 46750 22924 46756 22936
rect 46808 22924 46814 22976
rect 48314 22924 48320 22976
rect 48372 22964 48378 22976
rect 48685 22967 48743 22973
rect 48685 22964 48697 22967
rect 48372 22936 48697 22964
rect 48372 22924 48378 22936
rect 48685 22933 48697 22936
rect 48731 22933 48743 22967
rect 48685 22927 48743 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 3418 22760 3424 22772
rect 1636 22732 3424 22760
rect 1636 22720 1642 22732
rect 3418 22720 3424 22732
rect 3476 22720 3482 22772
rect 9493 22763 9551 22769
rect 3896 22732 8064 22760
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3896 22624 3924 22732
rect 4798 22652 4804 22704
rect 4856 22652 4862 22704
rect 7558 22692 7564 22704
rect 5920 22664 7564 22692
rect 3007 22596 3924 22624
rect 3973 22627 4031 22633
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 3973 22593 3985 22627
rect 4019 22624 4031 22627
rect 5920 22624 5948 22664
rect 7558 22652 7564 22664
rect 7616 22652 7622 22704
rect 4019 22596 5948 22624
rect 4019 22593 4031 22596
rect 3973 22587 4031 22593
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 7190 22624 7196 22636
rect 6687 22596 7196 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 7466 22584 7472 22636
rect 7524 22584 7530 22636
rect 2501 22559 2559 22565
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 2547 22528 2774 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 2746 22500 2774 22528
rect 7098 22516 7104 22568
rect 7156 22516 7162 22568
rect 7374 22516 7380 22568
rect 7432 22556 7438 22568
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7432 22528 7941 22556
rect 7432 22516 7438 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 8036 22556 8064 22732
rect 9493 22729 9505 22763
rect 9539 22760 9551 22763
rect 12618 22760 12624 22772
rect 9539 22732 12624 22760
rect 9539 22729 9551 22732
rect 9493 22723 9551 22729
rect 12618 22720 12624 22732
rect 12676 22760 12682 22772
rect 13538 22760 13544 22772
rect 12676 22732 13544 22760
rect 12676 22720 12682 22732
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 14182 22720 14188 22772
rect 14240 22760 14246 22772
rect 14550 22760 14556 22772
rect 14240 22732 14556 22760
rect 14240 22720 14246 22732
rect 14550 22720 14556 22732
rect 14608 22720 14614 22772
rect 18874 22760 18880 22772
rect 16868 22732 18880 22760
rect 9950 22652 9956 22704
rect 10008 22652 10014 22704
rect 12802 22652 12808 22704
rect 12860 22652 12866 22704
rect 15102 22652 15108 22704
rect 15160 22652 15166 22704
rect 11146 22584 11152 22636
rect 11204 22584 11210 22636
rect 11422 22584 11428 22636
rect 11480 22624 11486 22636
rect 11885 22627 11943 22633
rect 11885 22624 11897 22627
rect 11480 22596 11897 22624
rect 11480 22584 11486 22596
rect 11885 22593 11897 22596
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22624 14059 22627
rect 14642 22624 14648 22636
rect 14047 22596 14648 22624
rect 14047 22593 14059 22596
rect 14001 22587 14059 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 16868 22633 16896 22732
rect 18874 22720 18880 22732
rect 18932 22760 18938 22772
rect 19061 22763 19119 22769
rect 19061 22760 19073 22763
rect 18932 22732 19073 22760
rect 18932 22720 18938 22732
rect 19061 22729 19073 22732
rect 19107 22760 19119 22763
rect 19334 22760 19340 22772
rect 19107 22732 19340 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 21174 22720 21180 22772
rect 21232 22760 21238 22772
rect 21818 22760 21824 22772
rect 21232 22732 21824 22760
rect 21232 22720 21238 22732
rect 21818 22720 21824 22732
rect 21876 22720 21882 22772
rect 22002 22720 22008 22772
rect 22060 22760 22066 22772
rect 27246 22760 27252 22772
rect 22060 22720 22094 22760
rect 18506 22692 18512 22704
rect 18354 22664 18512 22692
rect 18506 22652 18512 22664
rect 18564 22692 18570 22704
rect 18969 22695 19027 22701
rect 18969 22692 18981 22695
rect 18564 22664 18981 22692
rect 18564 22652 18570 22664
rect 18969 22661 18981 22664
rect 19015 22692 19027 22695
rect 19242 22692 19248 22704
rect 19015 22664 19248 22692
rect 19015 22661 19027 22664
rect 18969 22655 19027 22661
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 22066 22692 22094 22720
rect 25240 22732 26004 22760
rect 22281 22695 22339 22701
rect 22281 22692 22293 22695
rect 22066 22664 22293 22692
rect 22281 22661 22293 22664
rect 22327 22661 22339 22695
rect 22281 22655 22339 22661
rect 23934 22652 23940 22704
rect 23992 22692 23998 22704
rect 24121 22695 24179 22701
rect 24121 22692 24133 22695
rect 23992 22664 24133 22692
rect 23992 22652 23998 22664
rect 24121 22661 24133 22664
rect 24167 22661 24179 22695
rect 24121 22655 24179 22661
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16853 22627 16911 22633
rect 16347 22596 16712 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 8036 22528 12434 22556
rect 7929 22519 7987 22525
rect 2746 22460 2780 22500
rect 2774 22448 2780 22460
rect 2832 22448 2838 22500
rect 4157 22491 4215 22497
rect 4157 22457 4169 22491
rect 4203 22488 4215 22491
rect 6454 22488 6460 22500
rect 4203 22460 6460 22488
rect 4203 22457 4215 22460
rect 4157 22451 4215 22457
rect 6454 22448 6460 22460
rect 6512 22448 6518 22500
rect 6825 22491 6883 22497
rect 6825 22457 6837 22491
rect 6871 22488 6883 22491
rect 9122 22488 9128 22500
rect 6871 22460 9128 22488
rect 6871 22457 6883 22460
rect 6825 22451 6883 22457
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 11701 22491 11759 22497
rect 11701 22488 11713 22491
rect 9232 22460 11713 22488
rect 3786 22380 3792 22432
rect 3844 22420 3850 22432
rect 5994 22420 6000 22432
rect 3844 22392 6000 22420
rect 3844 22380 3850 22392
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 7742 22380 7748 22432
rect 7800 22420 7806 22432
rect 9232 22420 9260 22460
rect 11701 22457 11713 22460
rect 11747 22457 11759 22491
rect 12406 22488 12434 22528
rect 15378 22488 15384 22500
rect 12406 22460 15384 22488
rect 11701 22451 11759 22457
rect 15378 22448 15384 22460
rect 15436 22448 15442 22500
rect 7800 22392 9260 22420
rect 9309 22423 9367 22429
rect 7800 22380 7806 22392
rect 9309 22389 9321 22423
rect 9355 22420 9367 22423
rect 11974 22420 11980 22432
rect 9355 22392 11980 22420
rect 9355 22389 9367 22392
rect 9309 22383 9367 22389
rect 11974 22380 11980 22392
rect 12032 22380 12038 22432
rect 12250 22380 12256 22432
rect 12308 22380 12314 22432
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 14461 22423 14519 22429
rect 14461 22420 14473 22423
rect 14424 22392 14473 22420
rect 14424 22380 14430 22392
rect 14461 22389 14473 22392
rect 14507 22420 14519 22423
rect 16206 22420 16212 22432
rect 14507 22392 16212 22420
rect 14507 22389 14519 22392
rect 14461 22383 14519 22389
rect 16206 22380 16212 22392
rect 16264 22380 16270 22432
rect 16684 22420 16712 22596
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 19429 22627 19487 22633
rect 19429 22624 19441 22627
rect 19392 22596 19441 22624
rect 19392 22584 19398 22596
rect 19429 22593 19441 22596
rect 19475 22593 19487 22627
rect 19429 22587 19487 22593
rect 20806 22584 20812 22636
rect 20864 22624 20870 22636
rect 21542 22624 21548 22636
rect 20864 22596 21548 22624
rect 20864 22584 20870 22596
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 22002 22624 22008 22636
rect 21784 22596 22008 22624
rect 21784 22584 21790 22596
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 23750 22624 23756 22636
rect 23414 22596 23756 22624
rect 23750 22584 23756 22596
rect 23808 22624 23814 22636
rect 24397 22627 24455 22633
rect 24397 22624 24409 22627
rect 23808 22596 24409 22624
rect 23808 22584 23814 22596
rect 24397 22593 24409 22596
rect 24443 22624 24455 22627
rect 24946 22624 24952 22636
rect 24443 22596 24952 22624
rect 24443 22593 24455 22596
rect 24397 22587 24455 22593
rect 24946 22584 24952 22596
rect 25004 22624 25010 22636
rect 25240 22624 25268 22732
rect 25866 22652 25872 22704
rect 25924 22692 25930 22704
rect 25976 22692 26004 22732
rect 26252 22732 27252 22760
rect 26252 22692 26280 22732
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 27338 22720 27344 22772
rect 27396 22720 27402 22772
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 27488 22732 30512 22760
rect 27488 22720 27494 22732
rect 25924 22664 26280 22692
rect 26329 22695 26387 22701
rect 25924 22652 25930 22664
rect 26329 22661 26341 22695
rect 26375 22692 26387 22695
rect 27448 22692 27476 22720
rect 26375 22664 27476 22692
rect 26375 22661 26387 22664
rect 26329 22655 26387 22661
rect 29454 22652 29460 22704
rect 29512 22692 29518 22704
rect 29549 22695 29607 22701
rect 29549 22692 29561 22695
rect 29512 22664 29561 22692
rect 29512 22652 29518 22664
rect 29549 22661 29561 22664
rect 29595 22692 29607 22695
rect 30006 22692 30012 22704
rect 29595 22664 30012 22692
rect 29595 22661 29607 22664
rect 29549 22655 29607 22661
rect 30006 22652 30012 22664
rect 30064 22652 30070 22704
rect 25004 22610 25268 22624
rect 25004 22596 25254 22610
rect 25004 22584 25010 22596
rect 27154 22584 27160 22636
rect 27212 22584 27218 22636
rect 27246 22584 27252 22636
rect 27304 22624 27310 22636
rect 27709 22627 27767 22633
rect 27709 22624 27721 22627
rect 27304 22596 27721 22624
rect 27304 22584 27310 22596
rect 27709 22593 27721 22596
rect 27755 22624 27767 22627
rect 28258 22624 28264 22636
rect 27755 22596 28264 22624
rect 27755 22593 27767 22596
rect 27709 22587 27767 22593
rect 28258 22584 28264 22596
rect 28316 22624 28322 22636
rect 28316 22610 28474 22624
rect 28316 22596 28488 22610
rect 28316 22584 28322 22596
rect 17126 22516 17132 22568
rect 17184 22516 17190 22568
rect 18414 22516 18420 22568
rect 18472 22556 18478 22568
rect 19705 22559 19763 22565
rect 19705 22556 19717 22559
rect 18472 22528 19717 22556
rect 18472 22516 18478 22528
rect 19705 22525 19717 22528
rect 19751 22525 19763 22559
rect 23290 22556 23296 22568
rect 19705 22519 19763 22525
rect 20732 22528 23296 22556
rect 18156 22460 18736 22488
rect 18156 22420 18184 22460
rect 16684 22392 18184 22420
rect 18322 22380 18328 22432
rect 18380 22420 18386 22432
rect 18601 22423 18659 22429
rect 18601 22420 18613 22423
rect 18380 22392 18613 22420
rect 18380 22380 18386 22392
rect 18601 22389 18613 22392
rect 18647 22389 18659 22423
rect 18708 22420 18736 22460
rect 20732 22420 20760 22528
rect 23290 22516 23296 22528
rect 23348 22516 23354 22568
rect 23658 22516 23664 22568
rect 23716 22556 23722 22568
rect 23716 22528 26556 22556
rect 23716 22516 23722 22528
rect 21818 22448 21824 22500
rect 21876 22488 21882 22500
rect 21876 22460 22094 22488
rect 21876 22448 21882 22460
rect 18708 22392 20760 22420
rect 18601 22383 18659 22389
rect 21634 22380 21640 22432
rect 21692 22380 21698 22432
rect 22066 22420 22094 22460
rect 23382 22448 23388 22500
rect 23440 22488 23446 22500
rect 24854 22488 24860 22500
rect 23440 22460 24860 22488
rect 23440 22448 23446 22460
rect 24854 22448 24860 22460
rect 24912 22448 24918 22500
rect 26528 22488 26556 22528
rect 26602 22516 26608 22568
rect 26660 22556 26666 22568
rect 28460 22556 28488 22596
rect 28902 22556 28908 22568
rect 26660 22528 28396 22556
rect 28460 22528 28908 22556
rect 26660 22516 26666 22528
rect 27522 22488 27528 22500
rect 26528 22460 27528 22488
rect 27522 22448 27528 22460
rect 27580 22448 27586 22500
rect 27706 22448 27712 22500
rect 27764 22488 27770 22500
rect 28074 22488 28080 22500
rect 27764 22460 28080 22488
rect 27764 22448 27770 22460
rect 28074 22448 28080 22460
rect 28132 22448 28138 22500
rect 23474 22420 23480 22432
rect 22066 22392 23480 22420
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 23753 22423 23811 22429
rect 23753 22389 23765 22423
rect 23799 22420 23811 22423
rect 24026 22420 24032 22432
rect 23799 22392 24032 22420
rect 23799 22389 23811 22392
rect 23753 22383 23811 22389
rect 24026 22380 24032 22392
rect 24084 22380 24090 22432
rect 24578 22380 24584 22432
rect 24636 22380 24642 22432
rect 25130 22380 25136 22432
rect 25188 22420 25194 22432
rect 26326 22420 26332 22432
rect 25188 22392 26332 22420
rect 25188 22380 25194 22392
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 28368 22420 28396 22528
rect 28902 22516 28908 22528
rect 28960 22516 28966 22568
rect 29825 22559 29883 22565
rect 29825 22525 29837 22559
rect 29871 22556 29883 22559
rect 30374 22556 30380 22568
rect 29871 22528 30380 22556
rect 29871 22525 29883 22528
rect 29825 22519 29883 22525
rect 29932 22420 29960 22528
rect 30374 22516 30380 22528
rect 30432 22516 30438 22568
rect 30484 22556 30512 22732
rect 30834 22720 30840 22772
rect 30892 22760 30898 22772
rect 32309 22763 32367 22769
rect 32309 22760 32321 22763
rect 30892 22732 32321 22760
rect 30892 22720 30898 22732
rect 32309 22729 32321 22732
rect 32355 22729 32367 22763
rect 32309 22723 32367 22729
rect 32677 22763 32735 22769
rect 32677 22729 32689 22763
rect 32723 22760 32735 22763
rect 33226 22760 33232 22772
rect 32723 22732 33232 22760
rect 32723 22729 32735 22732
rect 32677 22723 32735 22729
rect 33226 22720 33232 22732
rect 33284 22720 33290 22772
rect 34974 22760 34980 22772
rect 33704 22732 34980 22760
rect 33594 22692 33600 22704
rect 31680 22664 33600 22692
rect 30650 22584 30656 22636
rect 30708 22584 30714 22636
rect 30742 22584 30748 22636
rect 30800 22584 30806 22636
rect 31680 22633 31708 22664
rect 33594 22652 33600 22664
rect 33652 22652 33658 22704
rect 33704 22633 33732 22732
rect 34974 22720 34980 22732
rect 35032 22720 35038 22772
rect 35434 22720 35440 22772
rect 35492 22720 35498 22772
rect 35805 22763 35863 22769
rect 35805 22729 35817 22763
rect 35851 22760 35863 22763
rect 35894 22760 35900 22772
rect 35851 22732 35900 22760
rect 35851 22729 35863 22732
rect 35805 22723 35863 22729
rect 35894 22720 35900 22732
rect 35952 22720 35958 22772
rect 37461 22763 37519 22769
rect 37461 22729 37473 22763
rect 37507 22760 37519 22763
rect 38654 22760 38660 22772
rect 37507 22732 38660 22760
rect 37507 22729 37519 22732
rect 37461 22723 37519 22729
rect 33870 22652 33876 22704
rect 33928 22692 33934 22704
rect 33965 22695 34023 22701
rect 33965 22692 33977 22695
rect 33928 22664 33977 22692
rect 33928 22652 33934 22664
rect 33965 22661 33977 22664
rect 34011 22661 34023 22695
rect 33965 22655 34023 22661
rect 34606 22652 34612 22704
rect 34664 22652 34670 22704
rect 36354 22652 36360 22704
rect 36412 22692 36418 22704
rect 37274 22692 37280 22704
rect 36412 22664 37280 22692
rect 36412 22652 36418 22664
rect 37274 22652 37280 22664
rect 37332 22652 37338 22704
rect 31665 22627 31723 22633
rect 31665 22593 31677 22627
rect 31711 22593 31723 22627
rect 31665 22587 31723 22593
rect 32769 22627 32827 22633
rect 32769 22593 32781 22627
rect 32815 22624 32827 22627
rect 33689 22627 33747 22633
rect 32815 22596 32996 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 30837 22559 30895 22565
rect 30837 22556 30849 22559
rect 30484 22528 30849 22556
rect 30837 22525 30849 22528
rect 30883 22525 30895 22559
rect 32861 22559 32919 22565
rect 32861 22556 32873 22559
rect 30837 22519 30895 22525
rect 30944 22528 32873 22556
rect 30006 22448 30012 22500
rect 30064 22488 30070 22500
rect 30944 22488 30972 22528
rect 32861 22525 32873 22528
rect 32907 22525 32919 22559
rect 32861 22519 32919 22525
rect 30064 22460 30972 22488
rect 30064 22448 30070 22460
rect 31202 22448 31208 22500
rect 31260 22488 31266 22500
rect 32968 22488 32996 22596
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 35526 22584 35532 22636
rect 35584 22624 35590 22636
rect 36449 22627 36507 22633
rect 36449 22624 36461 22627
rect 35584 22596 36461 22624
rect 35584 22584 35590 22596
rect 36449 22593 36461 22596
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 34422 22516 34428 22568
rect 34480 22556 34486 22568
rect 36541 22559 36599 22565
rect 36541 22556 36553 22559
rect 34480 22528 36124 22556
rect 34480 22516 34486 22528
rect 33686 22488 33692 22500
rect 31260 22460 31616 22488
rect 32968 22460 33692 22488
rect 31260 22448 31266 22460
rect 28368 22392 29960 22420
rect 30190 22380 30196 22432
rect 30248 22420 30254 22432
rect 30285 22423 30343 22429
rect 30285 22420 30297 22423
rect 30248 22392 30297 22420
rect 30248 22380 30254 22392
rect 30285 22389 30297 22392
rect 30331 22389 30343 22423
rect 30285 22383 30343 22389
rect 30466 22380 30472 22432
rect 30524 22420 30530 22432
rect 30834 22420 30840 22432
rect 30524 22392 30840 22420
rect 30524 22380 30530 22392
rect 30834 22380 30840 22392
rect 30892 22380 30898 22432
rect 31478 22380 31484 22432
rect 31536 22380 31542 22432
rect 31588 22420 31616 22460
rect 33686 22448 33692 22460
rect 33744 22448 33750 22500
rect 36096 22497 36124 22528
rect 36464 22528 36553 22556
rect 36464 22500 36492 22528
rect 36541 22525 36553 22528
rect 36587 22525 36599 22559
rect 36541 22519 36599 22525
rect 36725 22559 36783 22565
rect 36725 22525 36737 22559
rect 36771 22556 36783 22559
rect 37476 22556 37504 22723
rect 38654 22720 38660 22732
rect 38712 22720 38718 22772
rect 38930 22720 38936 22772
rect 38988 22760 38994 22772
rect 43257 22763 43315 22769
rect 38988 22732 42104 22760
rect 38988 22720 38994 22732
rect 38838 22652 38844 22704
rect 38896 22692 38902 22704
rect 42076 22692 42104 22732
rect 43257 22729 43269 22763
rect 43303 22760 43315 22763
rect 44450 22760 44456 22772
rect 43303 22732 44456 22760
rect 43303 22729 43315 22732
rect 43257 22723 43315 22729
rect 44450 22720 44456 22732
rect 44508 22720 44514 22772
rect 46569 22763 46627 22769
rect 46569 22729 46581 22763
rect 46615 22760 46627 22763
rect 47578 22760 47584 22772
rect 46615 22732 47584 22760
rect 46615 22729 46627 22732
rect 46569 22723 46627 22729
rect 47578 22720 47584 22732
rect 47636 22720 47642 22772
rect 38896 22664 41460 22692
rect 38896 22652 38902 22664
rect 37826 22584 37832 22636
rect 37884 22584 37890 22636
rect 39206 22584 39212 22636
rect 39264 22624 39270 22636
rect 39485 22627 39543 22633
rect 39485 22624 39497 22627
rect 39264 22596 39497 22624
rect 39264 22584 39270 22596
rect 39485 22593 39497 22596
rect 39531 22593 39543 22627
rect 39485 22587 39543 22593
rect 39758 22584 39764 22636
rect 39816 22584 39822 22636
rect 40402 22584 40408 22636
rect 40460 22584 40466 22636
rect 40497 22627 40555 22633
rect 40497 22593 40509 22627
rect 40543 22624 40555 22627
rect 41138 22624 41144 22636
rect 40543 22596 41144 22624
rect 40543 22593 40555 22596
rect 40497 22587 40555 22593
rect 41138 22584 41144 22596
rect 41196 22584 41202 22636
rect 41432 22633 41460 22664
rect 42076 22664 42748 22692
rect 41417 22627 41475 22633
rect 41417 22593 41429 22627
rect 41463 22624 41475 22627
rect 41598 22624 41604 22636
rect 41463 22596 41604 22624
rect 41463 22593 41475 22596
rect 41417 22587 41475 22593
rect 41598 22584 41604 22596
rect 41656 22584 41662 22636
rect 42076 22633 42104 22664
rect 42061 22627 42119 22633
rect 42061 22593 42073 22627
rect 42107 22593 42119 22627
rect 42061 22587 42119 22593
rect 42610 22584 42616 22636
rect 42668 22584 42674 22636
rect 42720 22624 42748 22664
rect 44082 22652 44088 22704
rect 44140 22692 44146 22704
rect 44726 22692 44732 22704
rect 44140 22664 44732 22692
rect 44140 22652 44146 22664
rect 44726 22652 44732 22664
rect 44784 22692 44790 22704
rect 45189 22695 45247 22701
rect 45189 22692 45201 22695
rect 44784 22664 45201 22692
rect 44784 22652 44790 22664
rect 45189 22661 45201 22664
rect 45235 22661 45247 22695
rect 45189 22655 45247 22661
rect 45738 22652 45744 22704
rect 45796 22652 45802 22704
rect 45925 22695 45983 22701
rect 45925 22661 45937 22695
rect 45971 22692 45983 22695
rect 47302 22692 47308 22704
rect 45971 22664 47308 22692
rect 45971 22661 45983 22664
rect 45925 22655 45983 22661
rect 47302 22652 47308 22664
rect 47360 22652 47366 22704
rect 47854 22652 47860 22704
rect 47912 22692 47918 22704
rect 47949 22695 48007 22701
rect 47949 22692 47961 22695
rect 47912 22664 47961 22692
rect 47912 22652 47918 22664
rect 47949 22661 47961 22664
rect 47995 22661 48007 22695
rect 47949 22655 48007 22661
rect 44174 22624 44180 22636
rect 42720 22596 44180 22624
rect 44174 22584 44180 22596
rect 44232 22584 44238 22636
rect 47213 22627 47271 22633
rect 47213 22593 47225 22627
rect 47259 22624 47271 22627
rect 49142 22624 49148 22636
rect 47259 22596 49148 22624
rect 47259 22593 47271 22596
rect 47213 22587 47271 22593
rect 49142 22584 49148 22596
rect 49200 22584 49206 22636
rect 49234 22584 49240 22636
rect 49292 22624 49298 22636
rect 49329 22627 49387 22633
rect 49329 22624 49341 22627
rect 49292 22596 49341 22624
rect 49292 22584 49298 22596
rect 49329 22593 49341 22596
rect 49375 22593 49387 22627
rect 49329 22587 49387 22593
rect 36771 22528 37504 22556
rect 36771 22525 36783 22528
rect 36725 22519 36783 22525
rect 37642 22516 37648 22568
rect 37700 22556 37706 22568
rect 38838 22556 38844 22568
rect 37700 22528 38844 22556
rect 37700 22516 37706 22528
rect 38838 22516 38844 22528
rect 38896 22516 38902 22568
rect 38933 22559 38991 22565
rect 38933 22525 38945 22559
rect 38979 22556 38991 22559
rect 40589 22559 40647 22565
rect 40589 22556 40601 22559
rect 38979 22528 39160 22556
rect 38979 22525 38991 22528
rect 38933 22519 38991 22525
rect 36081 22491 36139 22497
rect 34992 22460 35848 22488
rect 33413 22423 33471 22429
rect 33413 22420 33425 22423
rect 31588 22392 33425 22420
rect 33413 22389 33425 22392
rect 33459 22420 33471 22423
rect 33962 22420 33968 22432
rect 33459 22392 33968 22420
rect 33459 22389 33471 22392
rect 33413 22383 33471 22389
rect 33962 22380 33968 22392
rect 34020 22380 34026 22432
rect 34514 22380 34520 22432
rect 34572 22420 34578 22432
rect 34992 22420 35020 22460
rect 35820 22432 35848 22460
rect 36081 22457 36093 22491
rect 36127 22457 36139 22491
rect 36081 22451 36139 22457
rect 36446 22448 36452 22500
rect 36504 22448 36510 22500
rect 37550 22488 37556 22500
rect 36556 22460 37556 22488
rect 34572 22392 35020 22420
rect 34572 22380 34578 22392
rect 35802 22380 35808 22432
rect 35860 22420 35866 22432
rect 36556 22420 36584 22460
rect 37550 22448 37556 22460
rect 37608 22448 37614 22500
rect 39132 22488 39160 22528
rect 39408 22528 40601 22556
rect 39298 22488 39304 22500
rect 39132 22460 39304 22488
rect 39298 22448 39304 22460
rect 39356 22448 39362 22500
rect 35860 22392 36584 22420
rect 35860 22380 35866 22392
rect 36906 22380 36912 22432
rect 36964 22420 36970 22432
rect 39408 22420 39436 22528
rect 40589 22525 40601 22528
rect 40635 22525 40647 22559
rect 40589 22519 40647 22525
rect 40678 22516 40684 22568
rect 40736 22556 40742 22568
rect 43717 22559 43775 22565
rect 43717 22556 43729 22559
rect 40736 22528 43729 22556
rect 40736 22516 40742 22528
rect 43717 22525 43729 22528
rect 43763 22525 43775 22559
rect 43717 22519 43775 22525
rect 39482 22448 39488 22500
rect 39540 22488 39546 22500
rect 41233 22491 41291 22497
rect 41233 22488 41245 22491
rect 39540 22460 41245 22488
rect 39540 22448 39546 22460
rect 41233 22457 41245 22460
rect 41279 22457 41291 22491
rect 43732 22488 43760 22519
rect 43990 22516 43996 22568
rect 44048 22516 44054 22568
rect 46658 22516 46664 22568
rect 46716 22556 46722 22568
rect 47578 22556 47584 22568
rect 46716 22528 47584 22556
rect 46716 22516 46722 22528
rect 47578 22516 47584 22528
rect 47636 22516 47642 22568
rect 47854 22516 47860 22568
rect 47912 22556 47918 22568
rect 48685 22559 48743 22565
rect 48685 22556 48697 22559
rect 47912 22528 48697 22556
rect 47912 22516 47918 22528
rect 48685 22525 48697 22528
rect 48731 22525 48743 22559
rect 48685 22519 48743 22525
rect 44542 22488 44548 22500
rect 43732 22460 44548 22488
rect 41233 22451 41291 22457
rect 44542 22448 44548 22460
rect 44600 22448 44606 22500
rect 45002 22448 45008 22500
rect 45060 22448 45066 22500
rect 47596 22488 47624 22516
rect 48317 22491 48375 22497
rect 48317 22488 48329 22491
rect 47596 22460 48329 22488
rect 48317 22457 48329 22460
rect 48363 22457 48375 22491
rect 48317 22451 48375 22457
rect 36964 22392 39436 22420
rect 36964 22380 36970 22392
rect 40034 22380 40040 22432
rect 40092 22380 40098 22432
rect 40310 22380 40316 22432
rect 40368 22420 40374 22432
rect 41877 22423 41935 22429
rect 41877 22420 41889 22423
rect 40368 22392 41889 22420
rect 40368 22380 40374 22392
rect 41877 22389 41889 22392
rect 41923 22389 41935 22423
rect 41877 22383 41935 22389
rect 45278 22380 45284 22432
rect 45336 22420 45342 22432
rect 47857 22423 47915 22429
rect 47857 22420 47869 22423
rect 45336 22392 47869 22420
rect 45336 22380 45342 22392
rect 47857 22389 47869 22392
rect 47903 22389 47915 22423
rect 47857 22383 47915 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 4246 22216 4252 22228
rect 2280 22188 4252 22216
rect 2280 22176 2286 22188
rect 4246 22176 4252 22188
rect 4304 22176 4310 22228
rect 11882 22176 11888 22228
rect 11940 22216 11946 22228
rect 12345 22219 12403 22225
rect 12345 22216 12357 22219
rect 11940 22188 12357 22216
rect 11940 22176 11946 22188
rect 12345 22185 12357 22188
rect 12391 22185 12403 22219
rect 15197 22219 15255 22225
rect 15197 22216 15209 22219
rect 12345 22179 12403 22185
rect 14108 22188 15209 22216
rect 3970 22108 3976 22160
rect 4028 22148 4034 22160
rect 4028 22120 6040 22148
rect 4028 22108 4034 22120
rect 3510 22040 3516 22092
rect 3568 22080 3574 22092
rect 3786 22080 3792 22092
rect 3568 22052 3792 22080
rect 3568 22040 3574 22052
rect 3786 22040 3792 22052
rect 3844 22040 3850 22092
rect 6012 22089 6040 22120
rect 5997 22083 6055 22089
rect 5997 22049 6009 22083
rect 6043 22049 6055 22083
rect 9674 22080 9680 22092
rect 5997 22043 6055 22049
rect 7852 22052 9680 22080
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 21981 3019 22015
rect 2961 21975 3019 21981
rect 1026 21904 1032 21956
rect 1084 21944 1090 21956
rect 1765 21947 1823 21953
rect 1765 21944 1777 21947
rect 1084 21916 1777 21944
rect 1084 21904 1090 21916
rect 1765 21913 1777 21916
rect 1811 21913 1823 21947
rect 1765 21907 1823 21913
rect 2976 21876 3004 21975
rect 5350 21972 5356 22024
rect 5408 21972 5414 22024
rect 7852 22021 7880 22052
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 11885 22083 11943 22089
rect 11885 22049 11897 22083
rect 11931 22080 11943 22083
rect 11974 22080 11980 22092
rect 11931 22052 11980 22080
rect 11931 22049 11943 22052
rect 11885 22043 11943 22049
rect 11974 22040 11980 22052
rect 12032 22040 12038 22092
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22080 13691 22083
rect 14108 22080 14136 22188
rect 15197 22185 15209 22188
rect 15243 22216 15255 22219
rect 17126 22216 17132 22228
rect 15243 22188 17132 22216
rect 15243 22185 15255 22188
rect 15197 22179 15255 22185
rect 17126 22176 17132 22188
rect 17184 22176 17190 22228
rect 19794 22176 19800 22228
rect 19852 22216 19858 22228
rect 27062 22216 27068 22228
rect 19852 22188 27068 22216
rect 19852 22176 19858 22188
rect 27062 22176 27068 22188
rect 27120 22176 27126 22228
rect 27614 22176 27620 22228
rect 27672 22216 27678 22228
rect 28353 22219 28411 22225
rect 28353 22216 28365 22219
rect 27672 22188 28365 22216
rect 27672 22176 27678 22188
rect 28353 22185 28365 22188
rect 28399 22185 28411 22219
rect 30650 22216 30656 22228
rect 28353 22179 28411 22185
rect 29656 22188 30656 22216
rect 14185 22151 14243 22157
rect 14185 22117 14197 22151
rect 14231 22148 14243 22151
rect 14366 22148 14372 22160
rect 14231 22120 14372 22148
rect 14231 22117 14243 22120
rect 14185 22111 14243 22117
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 17034 22108 17040 22160
rect 17092 22148 17098 22160
rect 17092 22120 17632 22148
rect 17092 22108 17098 22120
rect 17604 22089 17632 22120
rect 19702 22108 19708 22160
rect 19760 22148 19766 22160
rect 19760 22120 22048 22148
rect 19760 22108 19766 22120
rect 13679 22052 14136 22080
rect 17589 22083 17647 22089
rect 13679 22049 13691 22052
rect 13633 22043 13691 22049
rect 17589 22049 17601 22083
rect 17635 22049 17647 22083
rect 17589 22043 17647 22049
rect 18966 22040 18972 22092
rect 19024 22080 19030 22092
rect 22020 22089 22048 22120
rect 23474 22108 23480 22160
rect 23532 22148 23538 22160
rect 23532 22120 24532 22148
rect 23532 22108 23538 22120
rect 19889 22083 19947 22089
rect 19889 22080 19901 22083
rect 19024 22052 19901 22080
rect 19024 22040 19030 22052
rect 19889 22049 19901 22052
rect 19935 22049 19947 22083
rect 19889 22043 19947 22049
rect 22005 22083 22063 22089
rect 22005 22049 22017 22083
rect 22051 22049 22063 22083
rect 22005 22043 22063 22049
rect 22646 22040 22652 22092
rect 22704 22080 22710 22092
rect 23201 22083 23259 22089
rect 23201 22080 23213 22083
rect 22704 22052 23213 22080
rect 22704 22040 22710 22052
rect 23201 22049 23213 22052
rect 23247 22080 23259 22083
rect 23382 22080 23388 22092
rect 23247 22052 23388 22080
rect 23247 22049 23259 22052
rect 23201 22043 23259 22049
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 24504 22080 24532 22120
rect 24854 22108 24860 22160
rect 24912 22148 24918 22160
rect 24912 22120 26556 22148
rect 24912 22108 24918 22120
rect 25130 22080 25136 22092
rect 24504 22052 25136 22080
rect 25130 22040 25136 22052
rect 25188 22040 25194 22092
rect 26528 22089 26556 22120
rect 26602 22108 26608 22160
rect 26660 22148 26666 22160
rect 26660 22120 27108 22148
rect 26660 22108 26666 22120
rect 26513 22083 26571 22089
rect 26513 22049 26525 22083
rect 26559 22080 26571 22083
rect 27080 22080 27108 22120
rect 27154 22108 27160 22160
rect 27212 22148 27218 22160
rect 29656 22148 29684 22188
rect 30650 22176 30656 22188
rect 30708 22176 30714 22228
rect 31478 22176 31484 22228
rect 31536 22216 31542 22228
rect 31662 22216 31668 22228
rect 31536 22188 31668 22216
rect 31536 22176 31542 22188
rect 31662 22176 31668 22188
rect 31720 22176 31726 22228
rect 34238 22176 34244 22228
rect 34296 22176 34302 22228
rect 39114 22216 39120 22228
rect 36280 22188 39120 22216
rect 27212 22120 29684 22148
rect 27212 22108 27218 22120
rect 29730 22108 29736 22160
rect 29788 22108 29794 22160
rect 35434 22148 35440 22160
rect 33704 22120 35440 22148
rect 27709 22083 27767 22089
rect 27709 22080 27721 22083
rect 26559 22052 26593 22080
rect 27080 22052 27721 22080
rect 26559 22049 26571 22052
rect 26513 22043 26571 22049
rect 27709 22049 27721 22052
rect 27755 22049 27767 22083
rect 27709 22043 27767 22049
rect 28074 22040 28080 22092
rect 28132 22080 28138 22092
rect 28902 22080 28908 22092
rect 28132 22052 28908 22080
rect 28132 22040 28138 22052
rect 28902 22040 28908 22052
rect 28960 22040 28966 22092
rect 30190 22080 30196 22092
rect 29012 22052 30196 22080
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22012 7251 22015
rect 7837 22015 7895 22021
rect 7239 21984 7788 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 3510 21904 3516 21956
rect 3568 21944 3574 21956
rect 4157 21947 4215 21953
rect 4157 21944 4169 21947
rect 3568 21916 4169 21944
rect 3568 21904 3574 21916
rect 4157 21913 4169 21916
rect 4203 21913 4215 21947
rect 4157 21907 4215 21913
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 5684 21916 7665 21944
rect 5684 21904 5690 21916
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 7760 21944 7788 21984
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 8478 21944 8484 21956
rect 7760 21916 8484 21944
rect 7653 21907 7711 21913
rect 8478 21904 8484 21916
rect 8536 21904 8542 21956
rect 8294 21876 8300 21888
rect 2976 21848 8300 21876
rect 8294 21836 8300 21848
rect 8352 21836 8358 21888
rect 8386 21836 8392 21888
rect 8444 21836 8450 21888
rect 8588 21876 8616 21975
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 11606 21972 11612 22024
rect 11664 21972 11670 22024
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 14461 22015 14519 22021
rect 14461 22012 14473 22015
rect 13780 21984 14473 22012
rect 13780 21972 13786 21984
rect 14461 21981 14473 21984
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 16942 21972 16948 22024
rect 17000 21972 17006 22024
rect 18506 22012 18512 22024
rect 17052 21984 18512 22012
rect 11422 21904 11428 21956
rect 11480 21944 11486 21956
rect 12710 21944 12716 21956
rect 11480 21916 12716 21944
rect 11480 21904 11486 21916
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 14642 21904 14648 21956
rect 14700 21904 14706 21956
rect 16206 21904 16212 21956
rect 16264 21944 16270 21956
rect 16264 21916 16344 21944
rect 16264 21904 16270 21916
rect 12989 21879 13047 21885
rect 12989 21876 13001 21879
rect 8588 21848 13001 21876
rect 12989 21845 13001 21848
rect 13035 21845 13047 21879
rect 12989 21839 13047 21845
rect 13354 21836 13360 21888
rect 13412 21836 13418 21888
rect 13449 21879 13507 21885
rect 13449 21845 13461 21879
rect 13495 21876 13507 21879
rect 15286 21876 15292 21888
rect 13495 21848 15292 21876
rect 13495 21845 13507 21848
rect 13449 21839 13507 21845
rect 15286 21836 15292 21848
rect 15344 21836 15350 21888
rect 16316 21876 16344 21916
rect 16666 21904 16672 21956
rect 16724 21904 16730 21956
rect 17052 21876 17080 21984
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 18785 22015 18843 22021
rect 18785 21981 18797 22015
rect 18831 21981 18843 22015
rect 18785 21975 18843 21981
rect 17218 21904 17224 21956
rect 17276 21944 17282 21956
rect 18800 21944 18828 21975
rect 19426 21972 19432 22024
rect 19484 21972 19490 22024
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 22012 21235 22015
rect 21836 22012 21956 22028
rect 22278 22012 22284 22024
rect 21223 22000 22284 22012
rect 21223 21984 21864 22000
rect 21928 21984 22284 22000
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 22278 21972 22284 21984
rect 22336 22012 22342 22024
rect 22922 22012 22928 22024
rect 22336 21984 22928 22012
rect 22336 21972 22342 21984
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 22012 23075 22015
rect 23934 22012 23940 22024
rect 23063 21984 23940 22012
rect 23063 21981 23075 21984
rect 23017 21975 23075 21981
rect 23934 21972 23940 21984
rect 23992 21972 23998 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 24854 22012 24860 22024
rect 24075 21984 24860 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 24854 21972 24860 21984
rect 24912 21972 24918 22024
rect 25590 21972 25596 22024
rect 25648 22012 25654 22024
rect 25685 22015 25743 22021
rect 25685 22012 25697 22015
rect 25648 21984 25697 22012
rect 25648 21972 25654 21984
rect 25685 21981 25697 21984
rect 25731 22012 25743 22015
rect 26421 22015 26479 22021
rect 25731 21984 26372 22012
rect 25731 21981 25743 21984
rect 25685 21975 25743 21981
rect 21726 21944 21732 21956
rect 17276 21916 17816 21944
rect 18800 21916 21732 21944
rect 17276 21904 17282 21916
rect 16316 21848 17080 21876
rect 17788 21876 17816 21916
rect 21726 21904 21732 21916
rect 21784 21904 21790 21956
rect 21821 21947 21879 21953
rect 21821 21913 21833 21947
rect 21867 21913 21879 21947
rect 21821 21907 21879 21913
rect 21913 21947 21971 21953
rect 21913 21913 21925 21947
rect 21959 21944 21971 21947
rect 23474 21944 23480 21956
rect 21959 21916 23480 21944
rect 21959 21913 21971 21916
rect 21913 21907 21971 21913
rect 18966 21876 18972 21888
rect 17788 21848 18972 21876
rect 18966 21836 18972 21848
rect 19024 21836 19030 21888
rect 21450 21836 21456 21888
rect 21508 21836 21514 21888
rect 21836 21876 21864 21907
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 23566 21904 23572 21956
rect 23624 21944 23630 21956
rect 24949 21947 25007 21953
rect 23624 21916 24624 21944
rect 23624 21904 23630 21916
rect 22462 21876 22468 21888
rect 21836 21848 22468 21876
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 22612 21848 22661 21876
rect 22612 21836 22618 21848
rect 22649 21845 22661 21848
rect 22695 21845 22707 21879
rect 22649 21839 22707 21845
rect 22922 21836 22928 21888
rect 22980 21876 22986 21888
rect 23109 21879 23167 21885
rect 23109 21876 23121 21879
rect 22980 21848 23121 21876
rect 22980 21836 22986 21848
rect 23109 21845 23121 21848
rect 23155 21845 23167 21879
rect 23109 21839 23167 21845
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 24596 21885 24624 21916
rect 24949 21913 24961 21947
rect 24995 21944 25007 21947
rect 26050 21944 26056 21956
rect 24995 21916 26056 21944
rect 24995 21913 25007 21916
rect 24949 21907 25007 21913
rect 26050 21904 26056 21916
rect 26108 21904 26114 21956
rect 26344 21953 26372 21984
rect 26421 21981 26433 22015
rect 26467 22012 26479 22015
rect 29012 22012 29040 22052
rect 30190 22040 30196 22052
rect 30248 22040 30254 22092
rect 31570 22080 31576 22092
rect 30852 22052 31576 22080
rect 30852 22024 30880 22052
rect 31570 22040 31576 22052
rect 31628 22040 31634 22092
rect 32766 22040 32772 22092
rect 32824 22080 32830 22092
rect 33336 22089 33548 22094
rect 33704 22089 33732 22120
rect 35434 22108 35440 22120
rect 35492 22108 35498 22160
rect 33336 22083 33563 22089
rect 33336 22080 33517 22083
rect 32824 22066 33517 22080
rect 32824 22052 33364 22066
rect 32824 22040 32830 22052
rect 33505 22049 33517 22066
rect 33551 22080 33563 22083
rect 33689 22083 33747 22089
rect 33551 22052 33585 22080
rect 33551 22049 33563 22052
rect 33505 22043 33563 22049
rect 33689 22049 33701 22083
rect 33735 22049 33747 22083
rect 33689 22043 33747 22049
rect 33962 22040 33968 22092
rect 34020 22080 34026 22092
rect 35069 22083 35127 22089
rect 35069 22080 35081 22083
rect 34020 22052 35081 22080
rect 34020 22040 34026 22052
rect 35069 22049 35081 22052
rect 35115 22080 35127 22083
rect 35894 22080 35900 22092
rect 35115 22052 35900 22080
rect 35115 22049 35127 22052
rect 35069 22043 35127 22049
rect 35894 22040 35900 22052
rect 35952 22040 35958 22092
rect 36280 22089 36308 22188
rect 39114 22176 39120 22188
rect 39172 22176 39178 22228
rect 39206 22176 39212 22228
rect 39264 22216 39270 22228
rect 39393 22219 39451 22225
rect 39393 22216 39405 22219
rect 39264 22188 39405 22216
rect 39264 22176 39270 22188
rect 39393 22185 39405 22188
rect 39439 22216 39451 22219
rect 39574 22216 39580 22228
rect 39439 22188 39580 22216
rect 39439 22185 39451 22188
rect 39393 22179 39451 22185
rect 36814 22108 36820 22160
rect 36872 22108 36878 22160
rect 36265 22083 36323 22089
rect 36265 22049 36277 22083
rect 36311 22049 36323 22083
rect 37090 22080 37096 22092
rect 36265 22043 36323 22049
rect 36464 22052 37096 22080
rect 26467 21984 29040 22012
rect 26467 21981 26479 21984
rect 26421 21975 26479 21981
rect 29914 21972 29920 22024
rect 29972 21972 29978 22024
rect 30374 21972 30380 22024
rect 30432 22012 30438 22024
rect 30834 22012 30840 22024
rect 30432 21984 30840 22012
rect 30432 21972 30438 21984
rect 30834 21972 30840 21984
rect 30892 21972 30898 22024
rect 32214 21972 32220 22024
rect 32272 22012 32278 22024
rect 36464 22021 36492 22052
rect 37090 22040 37096 22052
rect 37148 22040 37154 22092
rect 37642 22040 37648 22092
rect 37700 22080 37706 22092
rect 37826 22080 37832 22092
rect 37700 22052 37832 22080
rect 37700 22040 37706 22052
rect 36449 22015 36507 22021
rect 32272 21984 33916 22012
rect 32272 21972 32278 21984
rect 26329 21947 26387 21953
rect 26329 21913 26341 21947
rect 26375 21944 26387 21947
rect 26878 21944 26884 21956
rect 26375 21916 26884 21944
rect 26375 21913 26387 21916
rect 26329 21907 26387 21913
rect 26878 21904 26884 21916
rect 26936 21904 26942 21956
rect 27525 21947 27583 21953
rect 27525 21913 27537 21947
rect 27571 21944 27583 21947
rect 27798 21944 27804 21956
rect 27571 21916 27804 21944
rect 27571 21913 27583 21916
rect 27525 21907 27583 21913
rect 27798 21904 27804 21916
rect 27856 21944 27862 21956
rect 28534 21944 28540 21956
rect 27856 21916 28540 21944
rect 27856 21904 27862 21916
rect 28534 21904 28540 21916
rect 28592 21904 28598 21956
rect 28718 21904 28724 21956
rect 28776 21904 28782 21956
rect 28813 21947 28871 21953
rect 28813 21913 28825 21947
rect 28859 21944 28871 21947
rect 30466 21944 30472 21956
rect 28859 21916 30472 21944
rect 28859 21913 28871 21916
rect 28813 21907 28871 21913
rect 30466 21904 30472 21916
rect 30524 21904 30530 21956
rect 31113 21947 31171 21953
rect 31113 21913 31125 21947
rect 31159 21944 31171 21947
rect 31202 21944 31208 21956
rect 31159 21916 31208 21944
rect 31159 21913 31171 21916
rect 31113 21907 31171 21913
rect 31202 21904 31208 21916
rect 31260 21904 31266 21956
rect 33686 21944 33692 21956
rect 32416 21916 33692 21944
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 23716 21848 23857 21876
rect 23716 21836 23722 21848
rect 23845 21845 23857 21848
rect 23891 21845 23903 21879
rect 23845 21839 23903 21845
rect 24581 21879 24639 21885
rect 24581 21845 24593 21879
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 24762 21836 24768 21888
rect 24820 21876 24826 21888
rect 25041 21879 25099 21885
rect 25041 21876 25053 21879
rect 24820 21848 25053 21876
rect 24820 21836 24826 21848
rect 25041 21845 25053 21848
rect 25087 21876 25099 21879
rect 25314 21876 25320 21888
rect 25087 21848 25320 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 25774 21836 25780 21888
rect 25832 21876 25838 21888
rect 25961 21879 26019 21885
rect 25961 21876 25973 21879
rect 25832 21848 25973 21876
rect 25832 21836 25838 21848
rect 25961 21845 25973 21848
rect 26007 21845 26019 21879
rect 25961 21839 26019 21845
rect 26694 21836 26700 21888
rect 26752 21876 26758 21888
rect 27157 21879 27215 21885
rect 27157 21876 27169 21879
rect 26752 21848 27169 21876
rect 26752 21836 26758 21848
rect 27157 21845 27169 21848
rect 27203 21845 27215 21879
rect 27157 21839 27215 21845
rect 27617 21879 27675 21885
rect 27617 21845 27629 21879
rect 27663 21876 27675 21879
rect 29638 21876 29644 21888
rect 27663 21848 29644 21876
rect 27663 21845 27675 21848
rect 27617 21839 27675 21845
rect 29638 21836 29644 21848
rect 29696 21876 29702 21888
rect 30193 21879 30251 21885
rect 30193 21876 30205 21879
rect 29696 21848 30205 21876
rect 29696 21836 29702 21848
rect 30193 21845 30205 21848
rect 30239 21845 30251 21879
rect 30193 21839 30251 21845
rect 30374 21836 30380 21888
rect 30432 21836 30438 21888
rect 30742 21836 30748 21888
rect 30800 21876 30806 21888
rect 32416 21876 32444 21916
rect 33686 21904 33692 21916
rect 33744 21904 33750 21956
rect 33888 21944 33916 21984
rect 36449 21981 36461 22015
rect 36495 21981 36507 22015
rect 37752 21998 37780 22052
rect 37826 22040 37832 22052
rect 37884 22040 37890 22092
rect 39117 22083 39175 22089
rect 39117 22049 39129 22083
rect 39163 22080 39175 22083
rect 39500 22080 39528 22188
rect 39574 22176 39580 22188
rect 39632 22176 39638 22228
rect 40221 22219 40279 22225
rect 40221 22185 40233 22219
rect 40267 22216 40279 22219
rect 40494 22216 40500 22228
rect 40267 22188 40500 22216
rect 40267 22185 40279 22188
rect 40221 22179 40279 22185
rect 40494 22176 40500 22188
rect 40552 22176 40558 22228
rect 44726 22176 44732 22228
rect 44784 22176 44790 22228
rect 47026 22176 47032 22228
rect 47084 22216 47090 22228
rect 47213 22219 47271 22225
rect 47213 22216 47225 22219
rect 47084 22188 47225 22216
rect 47084 22176 47090 22188
rect 47213 22185 47225 22188
rect 47259 22185 47271 22219
rect 47213 22179 47271 22185
rect 39850 22108 39856 22160
rect 39908 22108 39914 22160
rect 45278 22148 45284 22160
rect 39960 22120 42104 22148
rect 39163 22052 39528 22080
rect 39163 22049 39175 22052
rect 39117 22043 39175 22049
rect 36449 21975 36507 21981
rect 34057 21947 34115 21953
rect 34057 21944 34069 21947
rect 33888 21916 34069 21944
rect 34057 21913 34069 21916
rect 34103 21944 34115 21947
rect 34425 21947 34483 21953
rect 34425 21944 34437 21947
rect 34103 21916 34437 21944
rect 34103 21913 34115 21916
rect 34057 21907 34115 21913
rect 34425 21913 34437 21916
rect 34471 21944 34483 21947
rect 34606 21944 34612 21956
rect 34471 21916 34612 21944
rect 34471 21913 34483 21916
rect 34425 21907 34483 21913
rect 34606 21904 34612 21916
rect 34664 21904 34670 21956
rect 36538 21904 36544 21956
rect 36596 21944 36602 21956
rect 36596 21916 37504 21944
rect 36596 21904 36602 21916
rect 30800 21848 32444 21876
rect 30800 21836 30806 21848
rect 32490 21836 32496 21888
rect 32548 21876 32554 21888
rect 32585 21879 32643 21885
rect 32585 21876 32597 21879
rect 32548 21848 32597 21876
rect 32548 21836 32554 21848
rect 32585 21845 32597 21848
rect 32631 21845 32643 21879
rect 32585 21839 32643 21845
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32732 21848 33057 21876
rect 32732 21836 32738 21848
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 33410 21836 33416 21888
rect 33468 21836 33474 21888
rect 35158 21836 35164 21888
rect 35216 21836 35222 21888
rect 35250 21836 35256 21888
rect 35308 21836 35314 21888
rect 35621 21879 35679 21885
rect 35621 21845 35633 21879
rect 35667 21876 35679 21879
rect 36170 21876 36176 21888
rect 35667 21848 36176 21876
rect 35667 21845 35679 21848
rect 35621 21839 35679 21845
rect 36170 21836 36176 21848
rect 36228 21836 36234 21888
rect 36354 21836 36360 21888
rect 36412 21836 36418 21888
rect 37366 21836 37372 21888
rect 37424 21836 37430 21888
rect 37476 21876 37504 21916
rect 38838 21904 38844 21956
rect 38896 21904 38902 21956
rect 39298 21876 39304 21888
rect 37476 21848 39304 21876
rect 39298 21836 39304 21848
rect 39356 21876 39362 21888
rect 39960 21876 39988 22120
rect 40310 22040 40316 22092
rect 40368 22080 40374 22092
rect 40678 22080 40684 22092
rect 40368 22052 40684 22080
rect 40368 22040 40374 22052
rect 40678 22040 40684 22052
rect 40736 22040 40742 22092
rect 40880 22089 40908 22120
rect 40865 22083 40923 22089
rect 40865 22049 40877 22083
rect 40911 22049 40923 22083
rect 41966 22080 41972 22092
rect 40865 22043 40923 22049
rect 40972 22052 41972 22080
rect 40972 22012 41000 22052
rect 41966 22040 41972 22052
rect 42024 22040 42030 22092
rect 42076 22089 42104 22120
rect 42720 22120 45284 22148
rect 42061 22083 42119 22089
rect 42061 22049 42073 22083
rect 42107 22049 42119 22083
rect 42061 22043 42119 22049
rect 42150 22040 42156 22092
rect 42208 22080 42214 22092
rect 42521 22083 42579 22089
rect 42521 22080 42533 22083
rect 42208 22052 42533 22080
rect 42208 22040 42214 22052
rect 42521 22049 42533 22052
rect 42567 22080 42579 22083
rect 42720 22080 42748 22120
rect 45278 22108 45284 22120
rect 45336 22108 45342 22160
rect 42567 22052 42748 22080
rect 42567 22049 42579 22052
rect 42521 22043 42579 22049
rect 42794 22040 42800 22092
rect 42852 22080 42858 22092
rect 43073 22083 43131 22089
rect 43073 22080 43085 22083
rect 42852 22052 43085 22080
rect 42852 22040 42858 22052
rect 43073 22049 43085 22052
rect 43119 22080 43131 22083
rect 44361 22083 44419 22089
rect 44361 22080 44373 22083
rect 43119 22052 44373 22080
rect 43119 22049 43131 22052
rect 43073 22043 43131 22049
rect 44361 22049 44373 22052
rect 44407 22049 44419 22083
rect 44361 22043 44419 22049
rect 44542 22040 44548 22092
rect 44600 22040 44606 22092
rect 45186 22040 45192 22092
rect 45244 22040 45250 22092
rect 46842 22040 46848 22092
rect 46900 22080 46906 22092
rect 47029 22083 47087 22089
rect 47029 22080 47041 22083
rect 46900 22052 47041 22080
rect 46900 22040 46906 22052
rect 47029 22049 47041 22052
rect 47075 22049 47087 22083
rect 47029 22043 47087 22049
rect 47581 22083 47639 22089
rect 47581 22049 47593 22083
rect 47627 22080 47639 22083
rect 47670 22080 47676 22092
rect 47627 22052 47676 22080
rect 47627 22049 47639 22052
rect 47581 22043 47639 22049
rect 47670 22040 47676 22052
rect 47728 22040 47734 22092
rect 49510 22080 49516 22092
rect 48240 22052 49516 22080
rect 43349 22015 43407 22021
rect 40604 21984 41000 22012
rect 41386 21984 42748 22012
rect 40604 21888 40632 21984
rect 40678 21904 40684 21956
rect 40736 21944 40742 21956
rect 41386 21944 41414 21984
rect 40736 21916 41414 21944
rect 41785 21947 41843 21953
rect 40736 21904 40742 21916
rect 41785 21913 41797 21947
rect 41831 21944 41843 21947
rect 42610 21944 42616 21956
rect 41831 21916 42616 21944
rect 41831 21913 41843 21916
rect 41785 21907 41843 21913
rect 42610 21904 42616 21916
rect 42668 21904 42674 21956
rect 39356 21848 39988 21876
rect 39356 21836 39362 21848
rect 40586 21836 40592 21888
rect 40644 21836 40650 21888
rect 41230 21836 41236 21888
rect 41288 21876 41294 21888
rect 41417 21879 41475 21885
rect 41417 21876 41429 21879
rect 41288 21848 41429 21876
rect 41288 21836 41294 21848
rect 41417 21845 41429 21848
rect 41463 21845 41475 21879
rect 41417 21839 41475 21845
rect 41690 21836 41696 21888
rect 41748 21876 41754 21888
rect 42720 21885 42748 21984
rect 43349 21981 43361 22015
rect 43395 22012 43407 22015
rect 43438 22012 43444 22024
rect 43395 21984 43444 22012
rect 43395 21981 43407 21984
rect 43349 21975 43407 21981
rect 43438 21972 43444 21984
rect 43496 21972 43502 22024
rect 44174 21972 44180 22024
rect 44232 21972 44238 22024
rect 45462 21972 45468 22024
rect 45520 21972 45526 22024
rect 46750 21972 46756 22024
rect 46808 21972 46814 22024
rect 48240 22021 48268 22052
rect 49510 22040 49516 22052
rect 49568 22040 49574 22092
rect 48225 22015 48283 22021
rect 48225 21981 48237 22015
rect 48271 21981 48283 22015
rect 49326 22012 49332 22024
rect 48225 21975 48283 21981
rect 48792 21984 49332 22012
rect 42794 21904 42800 21956
rect 42852 21944 42858 21956
rect 45830 21944 45836 21956
rect 42852 21916 45836 21944
rect 42852 21904 42858 21916
rect 45830 21904 45836 21916
rect 45888 21904 45894 21956
rect 47486 21904 47492 21956
rect 47544 21944 47550 21956
rect 48792 21944 48820 21984
rect 49326 21972 49332 21984
rect 49384 21972 49390 22024
rect 47544 21916 48820 21944
rect 47544 21904 47550 21916
rect 41877 21879 41935 21885
rect 41877 21876 41889 21879
rect 41748 21848 41889 21876
rect 41748 21836 41754 21848
rect 41877 21845 41889 21848
rect 41923 21845 41935 21879
rect 41877 21839 41935 21845
rect 42705 21879 42763 21885
rect 42705 21845 42717 21879
rect 42751 21876 42763 21879
rect 45002 21876 45008 21888
rect 42751 21848 45008 21876
rect 42751 21845 42763 21848
rect 42705 21839 42763 21845
rect 45002 21836 45008 21848
rect 45060 21836 45066 21888
rect 46566 21836 46572 21888
rect 46624 21836 46630 21888
rect 48682 21836 48688 21888
rect 48740 21836 48746 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 5408 21644 9536 21672
rect 5408 21632 5414 21644
rect 3326 21564 3332 21616
rect 3384 21604 3390 21616
rect 3605 21607 3663 21613
rect 3605 21604 3617 21607
rect 3384 21576 3617 21604
rect 3384 21564 3390 21576
rect 3605 21573 3617 21576
rect 3651 21573 3663 21607
rect 3605 21567 3663 21573
rect 3694 21564 3700 21616
rect 3752 21604 3758 21616
rect 9508 21604 9536 21644
rect 9582 21632 9588 21684
rect 9640 21672 9646 21684
rect 10505 21675 10563 21681
rect 10505 21672 10517 21675
rect 9640 21644 10517 21672
rect 9640 21632 9646 21644
rect 10505 21641 10517 21644
rect 10551 21641 10563 21675
rect 11514 21672 11520 21684
rect 10505 21635 10563 21641
rect 10612 21644 11520 21672
rect 10612 21604 10640 21644
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 11701 21675 11759 21681
rect 11701 21641 11713 21675
rect 11747 21672 11759 21675
rect 11747 21644 12572 21672
rect 11747 21641 11759 21644
rect 11701 21635 11759 21641
rect 12544 21604 12572 21644
rect 12618 21632 12624 21684
rect 12676 21672 12682 21684
rect 13173 21675 13231 21681
rect 13173 21672 13185 21675
rect 12676 21644 13185 21672
rect 12676 21632 12682 21644
rect 13173 21641 13185 21644
rect 13219 21641 13231 21675
rect 13173 21635 13231 21641
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 13998 21632 14004 21684
rect 14056 21672 14062 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 14056 21644 17417 21672
rect 14056 21632 14062 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17405 21635 17463 21641
rect 17865 21675 17923 21681
rect 17865 21641 17877 21675
rect 17911 21672 17923 21675
rect 20990 21672 20996 21684
rect 17911 21644 20996 21672
rect 17911 21641 17923 21644
rect 17865 21635 17923 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 22830 21672 22836 21684
rect 21376 21644 22836 21672
rect 12802 21604 12808 21616
rect 3752 21576 8892 21604
rect 9508 21576 10640 21604
rect 10704 21576 12480 21604
rect 12544 21576 12808 21604
rect 3752 21564 3758 21576
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 1762 21428 1768 21480
rect 1820 21428 1826 21480
rect 2976 21332 3004 21499
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21536 5779 21539
rect 6362 21536 6368 21548
rect 5767 21508 6368 21536
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 6362 21496 6368 21508
rect 6420 21496 6426 21548
rect 6546 21496 6552 21548
rect 6604 21496 6610 21548
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21505 8447 21539
rect 8389 21499 8447 21505
rect 5810 21428 5816 21480
rect 5868 21468 5874 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 5868 21440 7021 21468
rect 5868 21428 5874 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 5905 21403 5963 21409
rect 5905 21369 5917 21403
rect 5951 21400 5963 21403
rect 8404 21400 8432 21499
rect 8864 21477 8892 21576
rect 10704 21545 10732 21576
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 12250 21496 12256 21548
rect 12308 21536 12314 21548
rect 12343 21539 12401 21545
rect 12343 21536 12355 21539
rect 12308 21508 12355 21536
rect 12308 21496 12314 21508
rect 12343 21505 12355 21508
rect 12389 21505 12401 21539
rect 12452 21536 12480 21576
rect 12802 21564 12808 21576
rect 12860 21564 12866 21616
rect 12912 21576 14228 21604
rect 12618 21536 12624 21548
rect 12452 21508 12624 21536
rect 12343 21499 12401 21505
rect 12618 21496 12624 21508
rect 12676 21496 12682 21548
rect 12912 21536 12940 21576
rect 12728 21508 12940 21536
rect 13265 21539 13323 21545
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21437 8907 21471
rect 8849 21431 8907 21437
rect 10229 21471 10287 21477
rect 10229 21437 10241 21471
rect 10275 21468 10287 21471
rect 11422 21468 11428 21480
rect 10275 21440 11428 21468
rect 10275 21437 10287 21440
rect 10229 21431 10287 21437
rect 11422 21428 11428 21440
rect 11480 21428 11486 21480
rect 12161 21471 12219 21477
rect 12161 21437 12173 21471
rect 12207 21468 12219 21471
rect 12434 21468 12440 21480
rect 12207 21440 12440 21468
rect 12207 21437 12219 21440
rect 12161 21431 12219 21437
rect 12434 21428 12440 21440
rect 12492 21428 12498 21480
rect 12728 21468 12756 21508
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 13906 21536 13912 21548
rect 13311 21508 13912 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 13906 21496 13912 21508
rect 13964 21496 13970 21548
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21505 14151 21539
rect 14200 21536 14228 21576
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 14829 21607 14887 21613
rect 14829 21604 14841 21607
rect 14332 21576 14841 21604
rect 14332 21564 14338 21576
rect 14829 21573 14841 21576
rect 14875 21573 14887 21607
rect 16206 21604 16212 21616
rect 16054 21576 16212 21604
rect 14829 21567 14887 21573
rect 16206 21564 16212 21576
rect 16264 21564 16270 21616
rect 16761 21607 16819 21613
rect 16761 21573 16773 21607
rect 16807 21604 16819 21607
rect 17218 21604 17224 21616
rect 16807 21576 17224 21604
rect 16807 21573 16819 21576
rect 16761 21567 16819 21573
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 18782 21604 18788 21616
rect 18432 21576 18788 21604
rect 17773 21539 17831 21545
rect 14200 21508 14596 21536
rect 14093 21499 14151 21505
rect 12636 21440 12756 21468
rect 5951 21372 8432 21400
rect 11149 21403 11207 21409
rect 5951 21369 5963 21372
rect 5905 21363 5963 21369
rect 11149 21369 11161 21403
rect 11195 21400 11207 21403
rect 11790 21400 11796 21412
rect 11195 21372 11796 21400
rect 11195 21369 11207 21372
rect 11149 21363 11207 21369
rect 11790 21360 11796 21372
rect 11848 21360 11854 21412
rect 11885 21403 11943 21409
rect 11885 21369 11897 21403
rect 11931 21400 11943 21403
rect 12342 21400 12348 21412
rect 11931 21372 12348 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 12342 21360 12348 21372
rect 12400 21400 12406 21412
rect 12636 21400 12664 21440
rect 13998 21400 14004 21412
rect 12400 21372 12664 21400
rect 12728 21372 14004 21400
rect 12400 21360 12406 21372
rect 7650 21332 7656 21344
rect 2976 21304 7656 21332
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11698 21332 11704 21344
rect 11379 21304 11704 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 11974 21292 11980 21344
rect 12032 21332 12038 21344
rect 12728 21332 12756 21372
rect 13998 21360 14004 21372
rect 14056 21360 14062 21412
rect 12032 21304 12756 21332
rect 12805 21335 12863 21341
rect 12032 21292 12038 21304
rect 12805 21301 12817 21335
rect 12851 21332 12863 21335
rect 13722 21332 13728 21344
rect 12851 21304 13728 21332
rect 12851 21301 12863 21304
rect 12805 21295 12863 21301
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 14108 21332 14136 21499
rect 14568 21480 14596 21508
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 18322 21536 18328 21548
rect 17819 21508 18328 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 14550 21428 14556 21480
rect 14608 21428 14614 21480
rect 15286 21428 15292 21480
rect 15344 21468 15350 21480
rect 16758 21468 16764 21480
rect 15344 21440 16764 21468
rect 15344 21428 15350 21440
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21468 18107 21471
rect 18432 21468 18460 21576
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 19426 21564 19432 21616
rect 19484 21564 19490 21616
rect 20622 21564 20628 21616
rect 20680 21604 20686 21616
rect 21376 21613 21404 21644
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 25406 21672 25412 21684
rect 23124 21644 25412 21672
rect 21177 21607 21235 21613
rect 21177 21604 21189 21607
rect 20680 21576 21189 21604
rect 20680 21564 20686 21576
rect 21177 21573 21189 21576
rect 21223 21573 21235 21607
rect 21177 21567 21235 21573
rect 21361 21607 21419 21613
rect 21361 21573 21373 21607
rect 21407 21573 21419 21607
rect 21361 21567 21419 21573
rect 21542 21564 21548 21616
rect 21600 21604 21606 21616
rect 23124 21604 23152 21644
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 26421 21675 26479 21681
rect 26421 21641 26433 21675
rect 26467 21641 26479 21675
rect 26421 21635 26479 21641
rect 24118 21604 24124 21616
rect 21600 21576 23152 21604
rect 23966 21576 24124 21604
rect 21600 21564 21606 21576
rect 24118 21564 24124 21576
rect 24176 21564 24182 21616
rect 26436 21604 26464 21635
rect 27614 21632 27620 21684
rect 27672 21672 27678 21684
rect 28353 21675 28411 21681
rect 28353 21672 28365 21675
rect 27672 21644 28365 21672
rect 27672 21632 27678 21644
rect 28353 21641 28365 21644
rect 28399 21641 28411 21675
rect 28353 21635 28411 21641
rect 28718 21632 28724 21684
rect 28776 21672 28782 21684
rect 30558 21672 30564 21684
rect 28776 21644 30564 21672
rect 28776 21632 28782 21644
rect 30558 21632 30564 21644
rect 30616 21672 30622 21684
rect 31113 21675 31171 21681
rect 30616 21644 30972 21672
rect 30616 21632 30622 21644
rect 27525 21607 27583 21613
rect 24228 21576 26464 21604
rect 26528 21576 27476 21604
rect 18095 21440 18460 21468
rect 18601 21471 18659 21477
rect 18095 21437 18107 21440
rect 18049 21431 18107 21437
rect 18601 21437 18613 21471
rect 18647 21437 18659 21471
rect 18601 21431 18659 21437
rect 17034 21360 17040 21412
rect 17092 21400 17098 21412
rect 17129 21403 17187 21409
rect 17129 21400 17141 21403
rect 17092 21372 17141 21400
rect 17092 21360 17098 21372
rect 17129 21369 17141 21372
rect 17175 21400 17187 21403
rect 18616 21400 18644 21431
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 19024 21440 22094 21468
rect 19024 21428 19030 21440
rect 17175 21372 18644 21400
rect 17175 21369 17187 21372
rect 17129 21363 17187 21369
rect 15930 21332 15936 21344
rect 14108 21304 15936 21332
rect 15930 21292 15936 21304
rect 15988 21292 15994 21344
rect 16301 21335 16359 21341
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 16574 21332 16580 21344
rect 16347 21304 16580 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 16945 21335 17003 21341
rect 16945 21301 16957 21335
rect 16991 21332 17003 21335
rect 17494 21332 17500 21344
rect 16991 21304 17500 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 18616 21332 18644 21372
rect 20349 21403 20407 21409
rect 20349 21369 20361 21403
rect 20395 21400 20407 21403
rect 21358 21400 21364 21412
rect 20395 21372 21364 21400
rect 20395 21369 20407 21372
rect 20349 21363 20407 21369
rect 21358 21360 21364 21372
rect 21416 21360 21422 21412
rect 22066 21400 22094 21440
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22244 21440 22477 21468
rect 22244 21428 22250 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22465 21431 22523 21437
rect 22572 21440 22753 21468
rect 22572 21400 22600 21440
rect 22741 21437 22753 21440
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 22830 21428 22836 21480
rect 22888 21468 22894 21480
rect 24228 21468 24256 21576
rect 25130 21496 25136 21548
rect 25188 21496 25194 21548
rect 26528 21536 26556 21576
rect 25332 21508 26556 21536
rect 26605 21539 26663 21545
rect 22888 21440 24256 21468
rect 22888 21428 22894 21440
rect 24578 21428 24584 21480
rect 24636 21468 24642 21480
rect 25222 21468 25228 21480
rect 24636 21440 25228 21468
rect 24636 21428 24642 21440
rect 25222 21428 25228 21440
rect 25280 21428 25286 21480
rect 24765 21403 24823 21409
rect 24765 21400 24777 21403
rect 22066 21372 22600 21400
rect 23768 21372 24777 21400
rect 19334 21332 19340 21344
rect 18616 21304 19340 21332
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 20625 21335 20683 21341
rect 20625 21332 20637 21335
rect 19484 21304 20637 21332
rect 19484 21292 19490 21304
rect 20625 21301 20637 21304
rect 20671 21332 20683 21335
rect 20809 21335 20867 21341
rect 20809 21332 20821 21335
rect 20671 21304 20821 21332
rect 20671 21301 20683 21304
rect 20625 21295 20683 21301
rect 20809 21301 20821 21304
rect 20855 21332 20867 21335
rect 21634 21332 21640 21344
rect 20855 21304 21640 21332
rect 20855 21301 20867 21304
rect 20809 21295 20867 21301
rect 21634 21292 21640 21304
rect 21692 21332 21698 21344
rect 21913 21335 21971 21341
rect 21913 21332 21925 21335
rect 21692 21304 21925 21332
rect 21692 21292 21698 21304
rect 21913 21301 21925 21304
rect 21959 21332 21971 21335
rect 22186 21332 22192 21344
rect 21959 21304 22192 21332
rect 21959 21301 21971 21304
rect 21913 21295 21971 21301
rect 22186 21292 22192 21304
rect 22244 21292 22250 21344
rect 22462 21292 22468 21344
rect 22520 21332 22526 21344
rect 23768 21332 23796 21372
rect 24765 21369 24777 21372
rect 24811 21369 24823 21403
rect 25332 21400 25360 21508
rect 26605 21505 26617 21539
rect 26651 21536 26663 21539
rect 26970 21536 26976 21548
rect 26651 21508 26976 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 26970 21496 26976 21508
rect 27028 21496 27034 21548
rect 27448 21536 27476 21576
rect 27525 21573 27537 21607
rect 27571 21604 27583 21607
rect 29822 21604 29828 21616
rect 27571 21576 29828 21604
rect 27571 21573 27583 21576
rect 27525 21567 27583 21573
rect 29822 21564 29828 21576
rect 29880 21564 29886 21616
rect 30944 21604 30972 21644
rect 31113 21641 31125 21675
rect 31159 21672 31171 21675
rect 31202 21672 31208 21684
rect 31159 21644 31208 21672
rect 31159 21641 31171 21644
rect 31113 21635 31171 21641
rect 31202 21632 31208 21644
rect 31260 21632 31266 21684
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21672 32827 21675
rect 33410 21672 33416 21684
rect 32815 21644 33416 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 33410 21632 33416 21644
rect 33468 21632 33474 21684
rect 33594 21632 33600 21684
rect 33652 21632 33658 21684
rect 34790 21632 34796 21684
rect 34848 21632 34854 21684
rect 35066 21632 35072 21684
rect 35124 21672 35130 21684
rect 36081 21675 36139 21681
rect 35124 21644 36032 21672
rect 35124 21632 35130 21644
rect 32582 21604 32588 21616
rect 30944 21576 32588 21604
rect 32582 21564 32588 21576
rect 32640 21564 32646 21616
rect 33612 21604 33640 21632
rect 35618 21604 35624 21616
rect 33612 21576 35624 21604
rect 35618 21564 35624 21576
rect 35676 21564 35682 21616
rect 36004 21604 36032 21644
rect 36081 21641 36093 21675
rect 36127 21672 36139 21675
rect 40034 21672 40040 21684
rect 36127 21644 40040 21672
rect 36127 21641 36139 21644
rect 36081 21635 36139 21641
rect 40034 21632 40040 21644
rect 40092 21632 40098 21684
rect 40954 21632 40960 21684
rect 41012 21672 41018 21684
rect 41322 21672 41328 21684
rect 41012 21644 41328 21672
rect 41012 21632 41018 21644
rect 41322 21632 41328 21644
rect 41380 21672 41386 21684
rect 41380 21644 42564 21672
rect 41380 21632 41386 21644
rect 36004 21576 37228 21604
rect 27448 21508 27844 21536
rect 25406 21428 25412 21480
rect 25464 21428 25470 21480
rect 26050 21428 26056 21480
rect 26108 21428 26114 21480
rect 27338 21428 27344 21480
rect 27396 21468 27402 21480
rect 27617 21471 27675 21477
rect 27617 21468 27629 21471
rect 27396 21440 27629 21468
rect 27396 21428 27402 21440
rect 27617 21437 27629 21440
rect 27663 21437 27675 21471
rect 27617 21431 27675 21437
rect 27709 21471 27767 21477
rect 27709 21437 27721 21471
rect 27755 21437 27767 21471
rect 27709 21431 27767 21437
rect 24765 21363 24823 21369
rect 25056 21372 25360 21400
rect 25424 21400 25452 21428
rect 27724 21400 27752 21431
rect 25424 21372 27752 21400
rect 27816 21400 27844 21508
rect 27890 21496 27896 21548
rect 27948 21536 27954 21548
rect 28721 21539 28779 21545
rect 28721 21536 28733 21539
rect 27948 21508 28733 21536
rect 27948 21496 27954 21508
rect 28721 21505 28733 21508
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 29917 21539 29975 21545
rect 29917 21505 29929 21539
rect 29963 21505 29975 21539
rect 29917 21499 29975 21505
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 30926 21536 30932 21548
rect 30055 21508 30932 21536
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 28810 21428 28816 21480
rect 28868 21428 28874 21480
rect 28902 21428 28908 21480
rect 28960 21428 28966 21480
rect 29454 21400 29460 21412
rect 27816 21372 29460 21400
rect 22520 21304 23796 21332
rect 24213 21335 24271 21341
rect 22520 21292 22526 21304
rect 24213 21301 24225 21335
rect 24259 21332 24271 21335
rect 25056 21332 25084 21372
rect 29454 21360 29460 21372
rect 29512 21360 29518 21412
rect 29932 21400 29960 21499
rect 30926 21496 30932 21508
rect 30984 21496 30990 21548
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 33502 21536 33508 21548
rect 31251 21508 33508 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 33502 21496 33508 21508
rect 33560 21496 33566 21548
rect 33686 21496 33692 21548
rect 33744 21536 33750 21548
rect 34701 21539 34759 21545
rect 34701 21536 34713 21539
rect 33744 21508 34713 21536
rect 33744 21496 33750 21508
rect 34701 21505 34713 21508
rect 34747 21536 34759 21539
rect 37200 21536 37228 21576
rect 37274 21564 37280 21616
rect 37332 21604 37338 21616
rect 37826 21604 37832 21616
rect 37332 21576 37832 21604
rect 37332 21564 37338 21576
rect 37826 21564 37832 21576
rect 37884 21604 37890 21616
rect 38562 21604 38568 21616
rect 37884 21576 38568 21604
rect 37884 21564 37890 21576
rect 38562 21564 38568 21576
rect 38620 21564 38626 21616
rect 39758 21604 39764 21616
rect 39514 21576 39764 21604
rect 39758 21564 39764 21576
rect 39816 21604 39822 21616
rect 40313 21607 40371 21613
rect 40313 21604 40325 21607
rect 39816 21576 40325 21604
rect 39816 21564 39822 21576
rect 40313 21573 40325 21576
rect 40359 21604 40371 21607
rect 40405 21607 40463 21613
rect 40405 21604 40417 21607
rect 40359 21576 40417 21604
rect 40359 21573 40371 21576
rect 40313 21567 40371 21573
rect 40405 21573 40417 21576
rect 40451 21604 40463 21607
rect 40589 21607 40647 21613
rect 40589 21604 40601 21607
rect 40451 21576 40601 21604
rect 40451 21573 40463 21576
rect 40405 21567 40463 21573
rect 40589 21573 40601 21576
rect 40635 21573 40647 21607
rect 42536 21604 42564 21644
rect 42610 21632 42616 21684
rect 42668 21632 42674 21684
rect 44450 21632 44456 21684
rect 44508 21672 44514 21684
rect 49234 21672 49240 21684
rect 44508 21644 49240 21672
rect 44508 21632 44514 21644
rect 49234 21632 49240 21644
rect 49292 21632 49298 21684
rect 44634 21604 44640 21616
rect 42536 21576 44640 21604
rect 40589 21567 40647 21573
rect 44634 21564 44640 21576
rect 44692 21604 44698 21616
rect 45281 21607 45339 21613
rect 45281 21604 45293 21607
rect 44692 21576 45293 21604
rect 44692 21564 44698 21576
rect 45281 21573 45293 21576
rect 45327 21573 45339 21607
rect 45281 21567 45339 21573
rect 45465 21607 45523 21613
rect 45465 21573 45477 21607
rect 45511 21604 45523 21607
rect 47026 21604 47032 21616
rect 45511 21576 47032 21604
rect 45511 21573 45523 21576
rect 45465 21567 45523 21573
rect 47026 21564 47032 21576
rect 47084 21564 47090 21616
rect 47121 21607 47179 21613
rect 47121 21573 47133 21607
rect 47167 21604 47179 21607
rect 48682 21604 48688 21616
rect 47167 21576 48688 21604
rect 47167 21573 47179 21576
rect 47121 21567 47179 21573
rect 48682 21564 48688 21576
rect 48740 21564 48746 21616
rect 37550 21536 37556 21548
rect 34747 21508 37044 21536
rect 37200 21508 37556 21536
rect 34747 21505 34759 21508
rect 34701 21499 34759 21505
rect 30193 21471 30251 21477
rect 30193 21437 30205 21471
rect 30239 21468 30251 21471
rect 30282 21468 30288 21480
rect 30239 21440 30288 21468
rect 30239 21437 30251 21440
rect 30193 21431 30251 21437
rect 30282 21428 30288 21440
rect 30340 21428 30346 21480
rect 30742 21428 30748 21480
rect 30800 21468 30806 21480
rect 31389 21471 31447 21477
rect 31389 21468 31401 21471
rect 30800 21440 31401 21468
rect 30800 21428 30806 21440
rect 31389 21437 31401 21440
rect 31435 21468 31447 21471
rect 31757 21471 31815 21477
rect 31757 21468 31769 21471
rect 31435 21440 31769 21468
rect 31435 21437 31447 21440
rect 31389 21431 31447 21437
rect 31757 21437 31769 21440
rect 31803 21437 31815 21471
rect 31757 21431 31815 21437
rect 33321 21471 33379 21477
rect 33321 21437 33333 21471
rect 33367 21437 33379 21471
rect 33321 21431 33379 21437
rect 34609 21471 34667 21477
rect 34609 21437 34621 21471
rect 34655 21468 34667 21471
rect 35986 21468 35992 21480
rect 34655 21440 35992 21468
rect 34655 21437 34667 21440
rect 34609 21431 34667 21437
rect 30558 21400 30564 21412
rect 29932 21372 30564 21400
rect 30558 21360 30564 21372
rect 30616 21360 30622 21412
rect 24259 21304 25084 21332
rect 24259 21301 24271 21304
rect 24213 21295 24271 21301
rect 25130 21292 25136 21344
rect 25188 21332 25194 21344
rect 25866 21332 25872 21344
rect 25188 21304 25872 21332
rect 25188 21292 25194 21304
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 26050 21292 26056 21344
rect 26108 21332 26114 21344
rect 27157 21335 27215 21341
rect 27157 21332 27169 21335
rect 26108 21304 27169 21332
rect 26108 21292 26114 21304
rect 27157 21301 27169 21304
rect 27203 21301 27215 21335
rect 27157 21295 27215 21301
rect 27246 21292 27252 21344
rect 27304 21332 27310 21344
rect 29549 21335 29607 21341
rect 29549 21332 29561 21335
rect 27304 21304 29561 21332
rect 27304 21292 27310 21304
rect 29549 21301 29561 21304
rect 29595 21301 29607 21335
rect 29549 21295 29607 21301
rect 30190 21292 30196 21344
rect 30248 21332 30254 21344
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 30248 21304 30757 21332
rect 30248 21292 30254 21304
rect 30745 21301 30757 21304
rect 30791 21301 30803 21335
rect 33336 21332 33364 21431
rect 35986 21428 35992 21440
rect 36044 21428 36050 21480
rect 36170 21428 36176 21480
rect 36228 21428 36234 21480
rect 36262 21428 36268 21480
rect 36320 21428 36326 21480
rect 37016 21477 37044 21508
rect 37550 21496 37556 21508
rect 37608 21496 37614 21548
rect 40218 21496 40224 21548
rect 40276 21536 40282 21548
rect 42426 21536 42432 21548
rect 40276 21508 42432 21536
rect 40276 21496 40282 21508
rect 42426 21496 42432 21508
rect 42484 21536 42490 21548
rect 42797 21539 42855 21545
rect 42797 21536 42809 21539
rect 42484 21508 42809 21536
rect 42484 21496 42490 21508
rect 42797 21505 42809 21508
rect 42843 21505 42855 21539
rect 42797 21499 42855 21505
rect 43346 21496 43352 21548
rect 43404 21536 43410 21548
rect 43441 21539 43499 21545
rect 43441 21536 43453 21539
rect 43404 21508 43453 21536
rect 43404 21496 43410 21508
rect 43441 21505 43453 21508
rect 43487 21505 43499 21539
rect 43441 21499 43499 21505
rect 43806 21496 43812 21548
rect 43864 21536 43870 21548
rect 43901 21539 43959 21545
rect 43901 21536 43913 21539
rect 43864 21508 43913 21536
rect 43864 21496 43870 21508
rect 43901 21505 43913 21508
rect 43947 21505 43959 21539
rect 43901 21499 43959 21505
rect 45186 21496 45192 21548
rect 45244 21536 45250 21548
rect 45833 21539 45891 21545
rect 45833 21536 45845 21539
rect 45244 21508 45845 21536
rect 45244 21496 45250 21508
rect 45833 21505 45845 21508
rect 45879 21505 45891 21539
rect 45833 21499 45891 21505
rect 46385 21539 46443 21545
rect 46385 21505 46397 21539
rect 46431 21536 46443 21539
rect 47394 21536 47400 21548
rect 46431 21508 47400 21536
rect 46431 21505 46443 21508
rect 46385 21499 46443 21505
rect 47394 21496 47400 21508
rect 47452 21496 47458 21548
rect 47578 21496 47584 21548
rect 47636 21536 47642 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47636 21508 47961 21536
rect 47636 21496 47642 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 49234 21496 49240 21548
rect 49292 21536 49298 21548
rect 49329 21539 49387 21545
rect 49329 21536 49341 21539
rect 49292 21508 49341 21536
rect 49292 21496 49298 21508
rect 49329 21505 49341 21508
rect 49375 21505 49387 21539
rect 49329 21499 49387 21505
rect 37001 21471 37059 21477
rect 37001 21437 37013 21471
rect 37047 21468 37059 21471
rect 37182 21468 37188 21480
rect 37047 21440 37188 21468
rect 37047 21437 37059 21440
rect 37001 21431 37059 21437
rect 37182 21428 37188 21440
rect 37240 21428 37246 21480
rect 37918 21428 37924 21480
rect 37976 21468 37982 21480
rect 38013 21471 38071 21477
rect 38013 21468 38025 21471
rect 37976 21440 38025 21468
rect 37976 21428 37982 21440
rect 38013 21437 38025 21440
rect 38059 21437 38071 21471
rect 38013 21431 38071 21437
rect 38286 21428 38292 21480
rect 38344 21468 38350 21480
rect 39574 21468 39580 21480
rect 38344 21440 39580 21468
rect 38344 21428 38350 21440
rect 39574 21428 39580 21440
rect 39632 21428 39638 21480
rect 39758 21428 39764 21480
rect 39816 21428 39822 21480
rect 41046 21428 41052 21480
rect 41104 21468 41110 21480
rect 41233 21471 41291 21477
rect 41233 21468 41245 21471
rect 41104 21440 41245 21468
rect 41104 21428 41110 21440
rect 41233 21437 41245 21440
rect 41279 21437 41291 21471
rect 41233 21431 41291 21437
rect 41506 21428 41512 21480
rect 41564 21428 41570 21480
rect 44177 21471 44235 21477
rect 44177 21437 44189 21471
rect 44223 21468 44235 21471
rect 44266 21468 44272 21480
rect 44223 21440 44272 21468
rect 44223 21437 44235 21440
rect 44177 21431 44235 21437
rect 44266 21428 44272 21440
rect 44324 21428 44330 21480
rect 46201 21471 46259 21477
rect 46201 21468 46213 21471
rect 44836 21440 46213 21468
rect 34238 21360 34244 21412
rect 34296 21400 34302 21412
rect 36538 21400 36544 21412
rect 34296 21372 36544 21400
rect 34296 21360 34302 21372
rect 36538 21360 36544 21372
rect 36596 21360 36602 21412
rect 36630 21360 36636 21412
rect 36688 21400 36694 21412
rect 36688 21372 38148 21400
rect 36688 21360 36694 21372
rect 33502 21332 33508 21344
rect 33336 21304 33508 21332
rect 30745 21295 30803 21301
rect 33502 21292 33508 21304
rect 33560 21292 33566 21344
rect 33965 21335 34023 21341
rect 33965 21301 33977 21335
rect 34011 21332 34023 21335
rect 34974 21332 34980 21344
rect 34011 21304 34980 21332
rect 34011 21301 34023 21304
rect 33965 21295 34023 21301
rect 34974 21292 34980 21304
rect 35032 21292 35038 21344
rect 35158 21292 35164 21344
rect 35216 21292 35222 21344
rect 35710 21292 35716 21344
rect 35768 21292 35774 21344
rect 35986 21292 35992 21344
rect 36044 21332 36050 21344
rect 36725 21335 36783 21341
rect 36725 21332 36737 21335
rect 36044 21304 36737 21332
rect 36044 21292 36050 21304
rect 36725 21301 36737 21304
rect 36771 21332 36783 21335
rect 36998 21332 37004 21344
rect 36771 21304 37004 21332
rect 36771 21301 36783 21304
rect 36725 21295 36783 21301
rect 36998 21292 37004 21304
rect 37056 21292 37062 21344
rect 37274 21292 37280 21344
rect 37332 21332 37338 21344
rect 37642 21332 37648 21344
rect 37332 21304 37648 21332
rect 37332 21292 37338 21304
rect 37642 21292 37648 21304
rect 37700 21292 37706 21344
rect 38120 21332 38148 21372
rect 39482 21360 39488 21412
rect 39540 21400 39546 21412
rect 40037 21403 40095 21409
rect 40037 21400 40049 21403
rect 39540 21372 40049 21400
rect 39540 21360 39546 21372
rect 40037 21369 40049 21372
rect 40083 21369 40095 21403
rect 40037 21363 40095 21369
rect 40862 21332 40868 21344
rect 38120 21304 40868 21332
rect 40862 21292 40868 21304
rect 40920 21292 40926 21344
rect 42794 21292 42800 21344
rect 42852 21332 42858 21344
rect 43257 21335 43315 21341
rect 43257 21332 43269 21335
rect 42852 21304 43269 21332
rect 42852 21292 42858 21304
rect 43257 21301 43269 21304
rect 43303 21301 43315 21335
rect 43257 21295 43315 21301
rect 43530 21292 43536 21344
rect 43588 21332 43594 21344
rect 44836 21332 44864 21440
rect 46201 21437 46213 21440
rect 46247 21437 46259 21471
rect 46201 21431 46259 21437
rect 47762 21428 47768 21480
rect 47820 21428 47826 21480
rect 46290 21360 46296 21412
rect 46348 21400 46354 21412
rect 46937 21403 46995 21409
rect 46937 21400 46949 21403
rect 46348 21372 46949 21400
rect 46348 21360 46354 21372
rect 46937 21369 46949 21372
rect 46983 21369 46995 21403
rect 46937 21363 46995 21369
rect 47210 21360 47216 21412
rect 47268 21400 47274 21412
rect 48685 21403 48743 21409
rect 48685 21400 48697 21403
rect 47268 21372 48697 21400
rect 47268 21360 47274 21372
rect 48685 21369 48697 21372
rect 48731 21369 48743 21403
rect 48685 21363 48743 21369
rect 43588 21304 44864 21332
rect 43588 21292 43594 21304
rect 47394 21292 47400 21344
rect 47452 21332 47458 21344
rect 48317 21335 48375 21341
rect 48317 21332 48329 21335
rect 47452 21304 48329 21332
rect 47452 21292 47458 21304
rect 48317 21301 48329 21304
rect 48363 21301 48375 21335
rect 48317 21295 48375 21301
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 12434 21128 12440 21140
rect 5368 21100 12440 21128
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 2866 20992 2872 21004
rect 2547 20964 2872 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 4154 20952 4160 21004
rect 4212 20952 4218 21004
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 5258 20924 5264 20936
rect 3007 20896 5264 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 5258 20884 5264 20896
rect 5316 20884 5322 20936
rect 5368 20933 5396 21100
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 14274 21088 14280 21140
rect 14332 21088 14338 21140
rect 19981 21131 20039 21137
rect 19981 21128 19993 21131
rect 14476 21100 19993 21128
rect 7834 21020 7840 21072
rect 7892 21060 7898 21072
rect 9217 21063 9275 21069
rect 9217 21060 9229 21063
rect 7892 21032 9229 21060
rect 7892 21020 7898 21032
rect 9217 21029 9229 21032
rect 9263 21029 9275 21063
rect 9217 21023 9275 21029
rect 10410 21020 10416 21072
rect 10468 21060 10474 21072
rect 11974 21060 11980 21072
rect 10468 21032 11980 21060
rect 10468 21020 10474 21032
rect 11974 21020 11980 21032
rect 12032 21020 12038 21072
rect 12158 21020 12164 21072
rect 12216 21060 12222 21072
rect 12713 21063 12771 21069
rect 12713 21060 12725 21063
rect 12216 21032 12725 21060
rect 12216 21020 12222 21032
rect 12713 21029 12725 21032
rect 12759 21029 12771 21063
rect 12713 21023 12771 21029
rect 5994 20952 6000 21004
rect 6052 20952 6058 21004
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 9950 20992 9956 21004
rect 6420 20964 9956 20992
rect 6420 20952 6426 20964
rect 9950 20952 9956 20964
rect 10008 20952 10014 21004
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 13354 20992 13360 21004
rect 10091 20964 13360 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 7193 20927 7251 20933
rect 7193 20893 7205 20927
rect 7239 20924 7251 20927
rect 8021 20927 8079 20933
rect 7239 20896 7880 20924
rect 7239 20893 7251 20896
rect 7193 20887 7251 20893
rect 7190 20748 7196 20800
rect 7248 20788 7254 20800
rect 7466 20788 7472 20800
rect 7248 20760 7472 20788
rect 7248 20748 7254 20760
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 7852 20797 7880 20896
rect 8021 20893 8033 20927
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20757 7895 20791
rect 8036 20788 8064 20887
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 8570 20924 8576 20936
rect 8444 20896 8576 20924
rect 8444 20884 8450 20896
rect 8570 20884 8576 20896
rect 8628 20884 8634 20936
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20924 9459 20927
rect 11146 20924 11152 20936
rect 9447 20896 11152 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 11146 20884 11152 20896
rect 11204 20884 11210 20936
rect 11330 20884 11336 20936
rect 11388 20884 11394 20936
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11848 20896 11989 20924
rect 11848 20884 11854 20896
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 12158 20884 12164 20936
rect 12216 20924 12222 20936
rect 13725 20927 13783 20933
rect 12216 20896 13584 20924
rect 12216 20884 12222 20896
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 8536 20828 11928 20856
rect 8536 20816 8542 20828
rect 10594 20788 10600 20800
rect 8036 20760 10600 20788
rect 7837 20751 7895 20757
rect 10594 20748 10600 20760
rect 10652 20748 10658 20800
rect 10689 20791 10747 20797
rect 10689 20757 10701 20791
rect 10735 20788 10747 20791
rect 11054 20788 11060 20800
rect 10735 20760 11060 20788
rect 10735 20757 10747 20760
rect 10689 20751 10747 20757
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11149 20791 11207 20797
rect 11149 20757 11161 20791
rect 11195 20788 11207 20791
rect 11238 20788 11244 20800
rect 11195 20760 11244 20788
rect 11195 20757 11207 20760
rect 11149 20751 11207 20757
rect 11238 20748 11244 20760
rect 11296 20748 11302 20800
rect 11900 20797 11928 20828
rect 12342 20816 12348 20868
rect 12400 20816 12406 20868
rect 12802 20816 12808 20868
rect 12860 20856 12866 20868
rect 12897 20859 12955 20865
rect 12897 20856 12909 20859
rect 12860 20828 12909 20856
rect 12860 20816 12866 20828
rect 12897 20825 12909 20828
rect 12943 20825 12955 20859
rect 12897 20819 12955 20825
rect 13556 20797 13584 20896
rect 13725 20893 13737 20927
rect 13771 20924 13783 20927
rect 14476 20924 14504 21100
rect 19981 21097 19993 21100
rect 20027 21097 20039 21131
rect 19981 21091 20039 21097
rect 24029 21131 24087 21137
rect 24029 21097 24041 21131
rect 24075 21128 24087 21131
rect 24302 21128 24308 21140
rect 24075 21100 24308 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 24302 21088 24308 21100
rect 24360 21088 24366 21140
rect 24762 21088 24768 21140
rect 24820 21088 24826 21140
rect 24946 21088 24952 21140
rect 25004 21128 25010 21140
rect 25004 21100 27384 21128
rect 25004 21088 25010 21100
rect 21177 21063 21235 21069
rect 21177 21060 21189 21063
rect 20548 21032 21189 21060
rect 14550 20952 14556 21004
rect 14608 20992 14614 21004
rect 16669 20995 16727 21001
rect 14608 20964 16068 20992
rect 14608 20952 14614 20964
rect 16040 20933 16068 20964
rect 16669 20961 16681 20995
rect 16715 20992 16727 20995
rect 18506 20992 18512 21004
rect 16715 20964 18512 20992
rect 16715 20961 16727 20964
rect 16669 20955 16727 20961
rect 18506 20952 18512 20964
rect 18564 20952 18570 21004
rect 18601 20995 18659 21001
rect 18601 20961 18613 20995
rect 18647 20992 18659 20995
rect 19702 20992 19708 21004
rect 18647 20964 19708 20992
rect 18647 20961 18659 20964
rect 18601 20955 18659 20961
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 19794 20952 19800 21004
rect 19852 20992 19858 21004
rect 20548 21001 20576 21032
rect 21177 21029 21189 21032
rect 21223 21029 21235 21063
rect 21177 21023 21235 21029
rect 23290 21020 23296 21072
rect 23348 21060 23354 21072
rect 23385 21063 23443 21069
rect 23385 21060 23397 21063
rect 23348 21032 23397 21060
rect 23348 21020 23354 21032
rect 23385 21029 23397 21032
rect 23431 21029 23443 21063
rect 23385 21023 23443 21029
rect 23474 21020 23480 21072
rect 23532 21060 23538 21072
rect 26050 21060 26056 21072
rect 23532 21032 26056 21060
rect 23532 21020 23538 21032
rect 26050 21020 26056 21032
rect 26108 21020 26114 21072
rect 27246 21060 27252 21072
rect 26160 21032 27252 21060
rect 20533 20995 20591 21001
rect 20533 20992 20545 20995
rect 19852 20964 20545 20992
rect 19852 20952 19858 20964
rect 20533 20961 20545 20964
rect 20579 20961 20591 20995
rect 22554 20992 22560 21004
rect 20533 20955 20591 20961
rect 21192 20964 22560 20992
rect 13771 20896 14504 20924
rect 16025 20927 16083 20933
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 16025 20893 16037 20927
rect 16071 20924 16083 20927
rect 17034 20924 17040 20936
rect 16071 20896 17040 20924
rect 16071 20893 16083 20896
rect 16025 20887 16083 20893
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20924 18935 20927
rect 19334 20924 19340 20936
rect 18923 20896 19340 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 19334 20884 19340 20896
rect 19392 20924 19398 20936
rect 20349 20927 20407 20933
rect 19392 20896 19564 20924
rect 19392 20884 19398 20896
rect 15749 20859 15807 20865
rect 15318 20828 15424 20856
rect 11885 20791 11943 20797
rect 11885 20757 11897 20791
rect 11931 20757 11943 20791
rect 11885 20751 11943 20757
rect 13541 20791 13599 20797
rect 13541 20757 13553 20791
rect 13587 20757 13599 20791
rect 13541 20751 13599 20757
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 15396 20788 15424 20828
rect 15749 20825 15761 20859
rect 15795 20856 15807 20859
rect 16114 20856 16120 20868
rect 15795 20828 16120 20856
rect 15795 20825 15807 20828
rect 15749 20819 15807 20825
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 18170 20828 19380 20856
rect 16206 20788 16212 20800
rect 13780 20760 16212 20788
rect 13780 20748 13786 20760
rect 16206 20748 16212 20760
rect 16264 20748 16270 20800
rect 16298 20748 16304 20800
rect 16356 20788 16362 20800
rect 17129 20791 17187 20797
rect 17129 20788 17141 20791
rect 16356 20760 17141 20788
rect 16356 20748 16362 20760
rect 17129 20757 17141 20760
rect 17175 20788 17187 20791
rect 18414 20788 18420 20800
rect 17175 20760 18420 20788
rect 17175 20757 17187 20760
rect 17129 20751 17187 20757
rect 18414 20748 18420 20760
rect 18472 20748 18478 20800
rect 19352 20797 19380 20828
rect 19337 20791 19395 20797
rect 19337 20757 19349 20791
rect 19383 20788 19395 20791
rect 19426 20788 19432 20800
rect 19383 20760 19432 20788
rect 19383 20757 19395 20760
rect 19337 20751 19395 20757
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 19536 20797 19564 20896
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 21192 20924 21220 20964
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 22646 20952 22652 21004
rect 22704 20952 22710 21004
rect 26160 21001 26188 21032
rect 27246 21020 27252 21032
rect 27304 21020 27310 21072
rect 25317 20995 25375 21001
rect 25317 20992 25329 20995
rect 24688 20964 25329 20992
rect 20395 20896 21220 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 22922 20884 22928 20936
rect 22980 20884 22986 20936
rect 23492 20896 24164 20924
rect 20441 20859 20499 20865
rect 20441 20825 20453 20859
rect 20487 20856 20499 20859
rect 20487 20828 21312 20856
rect 20487 20825 20499 20828
rect 20441 20819 20499 20825
rect 19521 20791 19579 20797
rect 19521 20757 19533 20791
rect 19567 20788 19579 20791
rect 19610 20788 19616 20800
rect 19567 20760 19616 20788
rect 19567 20757 19579 20760
rect 19521 20751 19579 20757
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 21284 20788 21312 20828
rect 22186 20816 22192 20868
rect 22244 20856 22250 20868
rect 23492 20856 23520 20896
rect 24136 20868 24164 20896
rect 24302 20884 24308 20936
rect 24360 20924 24366 20936
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24360 20896 24593 20924
rect 24360 20884 24366 20896
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24688 20868 24716 20964
rect 25317 20961 25329 20964
rect 25363 20961 25375 20995
rect 25317 20955 25375 20961
rect 26145 20995 26203 21001
rect 26145 20961 26157 20995
rect 26191 20961 26203 20995
rect 26145 20955 26203 20961
rect 26234 20952 26240 21004
rect 26292 20952 26298 21004
rect 26418 20952 26424 21004
rect 26476 20992 26482 21004
rect 26697 20995 26755 21001
rect 26697 20992 26709 20995
rect 26476 20964 26709 20992
rect 26476 20952 26482 20964
rect 26697 20961 26709 20964
rect 26743 20992 26755 20995
rect 27154 20992 27160 21004
rect 26743 20964 27160 20992
rect 26743 20961 26755 20964
rect 26697 20955 26755 20961
rect 27154 20952 27160 20964
rect 27212 20952 27218 21004
rect 24762 20884 24768 20936
rect 24820 20924 24826 20936
rect 26053 20927 26111 20933
rect 24820 20896 25912 20924
rect 24820 20884 24826 20896
rect 22244 20828 23520 20856
rect 22244 20816 22250 20828
rect 23566 20816 23572 20868
rect 23624 20816 23630 20868
rect 24118 20816 24124 20868
rect 24176 20856 24182 20868
rect 24213 20859 24271 20865
rect 24213 20856 24225 20859
rect 24176 20828 24225 20856
rect 24176 20816 24182 20828
rect 24213 20825 24225 20828
rect 24259 20856 24271 20859
rect 24670 20856 24676 20868
rect 24259 20828 24676 20856
rect 24259 20825 24271 20828
rect 24213 20819 24271 20825
rect 24670 20816 24676 20828
rect 24728 20856 24734 20868
rect 25133 20859 25191 20865
rect 25133 20856 25145 20859
rect 24728 20828 25145 20856
rect 24728 20816 24734 20828
rect 25133 20825 25145 20828
rect 25179 20825 25191 20859
rect 25774 20856 25780 20868
rect 25133 20819 25191 20825
rect 25332 20828 25780 20856
rect 25332 20788 25360 20828
rect 25774 20816 25780 20828
rect 25832 20816 25838 20868
rect 21284 20760 25360 20788
rect 25406 20748 25412 20800
rect 25464 20788 25470 20800
rect 25685 20791 25743 20797
rect 25685 20788 25697 20791
rect 25464 20760 25697 20788
rect 25464 20748 25470 20760
rect 25685 20757 25697 20760
rect 25731 20757 25743 20791
rect 25884 20788 25912 20896
rect 26053 20893 26065 20927
rect 26099 20893 26111 20927
rect 26053 20887 26111 20893
rect 26068 20856 26096 20887
rect 26510 20884 26516 20936
rect 26568 20924 26574 20936
rect 26881 20927 26939 20933
rect 26881 20924 26893 20927
rect 26568 20896 26893 20924
rect 26568 20884 26574 20896
rect 26881 20893 26893 20896
rect 26927 20893 26939 20927
rect 27356 20924 27384 21100
rect 29730 21088 29736 21140
rect 29788 21088 29794 21140
rect 30650 21088 30656 21140
rect 30708 21128 30714 21140
rect 30837 21131 30895 21137
rect 30837 21128 30849 21131
rect 30708 21100 30849 21128
rect 30708 21088 30714 21100
rect 30837 21097 30849 21100
rect 30883 21097 30895 21131
rect 30837 21091 30895 21097
rect 31018 21088 31024 21140
rect 31076 21088 31082 21140
rect 35710 21128 35716 21140
rect 31312 21100 35716 21128
rect 29089 21063 29147 21069
rect 29089 21029 29101 21063
rect 29135 21060 29147 21063
rect 30098 21060 30104 21072
rect 29135 21032 30104 21060
rect 29135 21029 29147 21032
rect 29089 21023 29147 21029
rect 30098 21020 30104 21032
rect 30156 21020 30162 21072
rect 30285 21063 30343 21069
rect 30285 21029 30297 21063
rect 30331 21060 30343 21063
rect 31036 21060 31064 21088
rect 30331 21032 31064 21060
rect 30331 21029 30343 21032
rect 30285 21023 30343 21029
rect 27890 20952 27896 21004
rect 27948 20952 27954 21004
rect 31312 21001 31340 21100
rect 35710 21088 35716 21100
rect 35768 21088 35774 21140
rect 36722 21088 36728 21140
rect 36780 21128 36786 21140
rect 37642 21128 37648 21140
rect 36780 21100 37648 21128
rect 36780 21088 36786 21100
rect 37642 21088 37648 21100
rect 37700 21088 37706 21140
rect 37734 21088 37740 21140
rect 37792 21128 37798 21140
rect 37792 21100 39344 21128
rect 37792 21088 37798 21100
rect 34054 21020 34060 21072
rect 34112 21060 34118 21072
rect 35066 21060 35072 21072
rect 34112 21032 35072 21060
rect 34112 21020 34118 21032
rect 35066 21020 35072 21032
rect 35124 21020 35130 21072
rect 37366 21020 37372 21072
rect 37424 21060 37430 21072
rect 38102 21060 38108 21072
rect 37424 21032 38108 21060
rect 37424 21020 37430 21032
rect 38102 21020 38108 21032
rect 38160 21020 38166 21072
rect 39316 21060 39344 21100
rect 39574 21088 39580 21140
rect 39632 21128 39638 21140
rect 39632 21100 40816 21128
rect 39632 21088 39638 21100
rect 39316 21032 40724 21060
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20992 28595 20995
rect 31297 20995 31355 21001
rect 28583 20964 30144 20992
rect 28583 20961 28595 20964
rect 28537 20955 28595 20961
rect 28629 20927 28687 20933
rect 28629 20924 28641 20927
rect 27356 20896 28641 20924
rect 26881 20887 26939 20893
rect 28629 20893 28641 20896
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28718 20884 28724 20936
rect 28776 20884 28782 20936
rect 29914 20884 29920 20936
rect 29972 20884 29978 20936
rect 30116 20924 30144 20964
rect 31297 20961 31309 20995
rect 31343 20961 31355 20995
rect 31297 20955 31355 20961
rect 31481 20995 31539 21001
rect 31481 20961 31493 20995
rect 31527 20992 31539 20995
rect 32306 20992 32312 21004
rect 31527 20964 32312 20992
rect 31527 20961 31539 20964
rect 31481 20955 31539 20961
rect 32306 20952 32312 20964
rect 32364 20992 32370 21004
rect 32769 20995 32827 21001
rect 32769 20992 32781 20995
rect 32364 20964 32781 20992
rect 32364 20952 32370 20964
rect 32769 20961 32781 20964
rect 32815 20961 32827 20995
rect 32769 20955 32827 20961
rect 33962 20952 33968 21004
rect 34020 20992 34026 21004
rect 34238 20992 34244 21004
rect 34020 20964 34244 20992
rect 34020 20952 34026 20964
rect 34238 20952 34244 20964
rect 34296 20952 34302 21004
rect 35894 20952 35900 21004
rect 35952 20992 35958 21004
rect 36357 20995 36415 21001
rect 36357 20992 36369 20995
rect 35952 20964 36369 20992
rect 35952 20952 35958 20964
rect 36357 20961 36369 20964
rect 36403 20992 36415 20995
rect 36906 20992 36912 21004
rect 36403 20964 36912 20992
rect 36403 20961 36415 20964
rect 36357 20955 36415 20961
rect 36906 20952 36912 20964
rect 36964 20952 36970 21004
rect 37918 20992 37924 21004
rect 37568 20964 37924 20992
rect 32398 20924 32404 20936
rect 30116 20896 32404 20924
rect 32398 20884 32404 20896
rect 32456 20884 32462 20936
rect 32490 20884 32496 20936
rect 32548 20884 32554 20936
rect 34606 20884 34612 20936
rect 34664 20924 34670 20936
rect 35250 20924 35256 20936
rect 34664 20896 35256 20924
rect 34664 20884 34670 20896
rect 35250 20884 35256 20896
rect 35308 20884 35314 20936
rect 36633 20927 36691 20933
rect 36633 20893 36645 20927
rect 36679 20924 36691 20927
rect 36679 20896 37228 20924
rect 36679 20893 36691 20896
rect 36633 20887 36691 20893
rect 26786 20856 26792 20868
rect 26068 20828 26792 20856
rect 26786 20816 26792 20828
rect 26844 20816 26850 20868
rect 27338 20816 27344 20868
rect 27396 20816 27402 20868
rect 28810 20816 28816 20868
rect 28868 20856 28874 20868
rect 30466 20856 30472 20868
rect 28868 20828 30472 20856
rect 28868 20816 28874 20828
rect 30466 20816 30472 20828
rect 30524 20816 30530 20868
rect 30926 20816 30932 20868
rect 30984 20856 30990 20868
rect 31754 20856 31760 20868
rect 30984 20828 31760 20856
rect 30984 20816 30990 20828
rect 31754 20816 31760 20828
rect 31812 20816 31818 20868
rect 31846 20816 31852 20868
rect 31904 20856 31910 20868
rect 31941 20859 31999 20865
rect 31941 20856 31953 20859
rect 31904 20828 31953 20856
rect 31904 20816 31910 20828
rect 31941 20825 31953 20828
rect 31987 20856 31999 20859
rect 32858 20856 32864 20868
rect 31987 20828 32864 20856
rect 31987 20825 31999 20828
rect 31941 20819 31999 20825
rect 32858 20816 32864 20828
rect 32916 20816 32922 20868
rect 37200 20865 37228 20896
rect 37568 20868 37596 20964
rect 37918 20952 37924 20964
rect 37976 20992 37982 21004
rect 39393 20995 39451 21001
rect 39393 20992 39405 20995
rect 37976 20964 39405 20992
rect 37976 20952 37982 20964
rect 39393 20961 39405 20964
rect 39439 20992 39451 20995
rect 39482 20992 39488 21004
rect 39439 20964 39488 20992
rect 39439 20961 39451 20964
rect 39393 20955 39451 20961
rect 39482 20952 39488 20964
rect 39540 20952 39546 21004
rect 39758 20952 39764 21004
rect 39816 20992 39822 21004
rect 40589 20995 40647 21001
rect 40589 20992 40601 20995
rect 39816 20964 40601 20992
rect 39816 20952 39822 20964
rect 40589 20961 40601 20964
rect 40635 20961 40647 20995
rect 40589 20955 40647 20961
rect 40497 20927 40555 20933
rect 40497 20924 40509 20927
rect 39868 20896 40509 20924
rect 37185 20859 37243 20865
rect 33152 20828 33258 20856
rect 34164 20828 34928 20856
rect 30006 20788 30012 20800
rect 25884 20760 30012 20788
rect 25685 20751 25743 20757
rect 30006 20748 30012 20760
rect 30064 20748 30070 20800
rect 30098 20748 30104 20800
rect 30156 20788 30162 20800
rect 30377 20791 30435 20797
rect 30377 20788 30389 20791
rect 30156 20760 30389 20788
rect 30156 20748 30162 20760
rect 30377 20757 30389 20760
rect 30423 20757 30435 20791
rect 30377 20751 30435 20757
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 32214 20748 32220 20800
rect 32272 20788 32278 20800
rect 33152 20788 33180 20828
rect 32272 20760 33180 20788
rect 32272 20748 32278 20760
rect 33686 20748 33692 20800
rect 33744 20788 33750 20800
rect 34164 20788 34192 20828
rect 34900 20797 34928 20828
rect 37185 20825 37197 20859
rect 37231 20856 37243 20859
rect 37550 20856 37556 20868
rect 37231 20828 37556 20856
rect 37231 20825 37243 20828
rect 37185 20819 37243 20825
rect 37550 20816 37556 20828
rect 37608 20816 37614 20868
rect 37752 20828 37950 20856
rect 37752 20800 37780 20828
rect 39114 20816 39120 20868
rect 39172 20856 39178 20868
rect 39758 20856 39764 20868
rect 39172 20828 39764 20856
rect 39172 20816 39178 20828
rect 39758 20816 39764 20828
rect 39816 20816 39822 20868
rect 33744 20760 34192 20788
rect 34885 20791 34943 20797
rect 33744 20748 33750 20760
rect 34885 20757 34897 20791
rect 34931 20788 34943 20791
rect 36262 20788 36268 20800
rect 34931 20760 36268 20788
rect 34931 20757 34943 20760
rect 34885 20751 34943 20757
rect 36262 20748 36268 20760
rect 36320 20748 36326 20800
rect 36906 20748 36912 20800
rect 36964 20748 36970 20800
rect 37274 20748 37280 20800
rect 37332 20788 37338 20800
rect 37734 20788 37740 20800
rect 37332 20760 37740 20788
rect 37332 20748 37338 20760
rect 37734 20748 37740 20760
rect 37792 20748 37798 20800
rect 38746 20748 38752 20800
rect 38804 20788 38810 20800
rect 39868 20788 39896 20896
rect 40497 20893 40509 20896
rect 40543 20893 40555 20927
rect 40696 20924 40724 21032
rect 40788 20992 40816 21100
rect 41690 21088 41696 21140
rect 41748 21128 41754 21140
rect 42797 21131 42855 21137
rect 42797 21128 42809 21131
rect 41748 21100 42809 21128
rect 41748 21088 41754 21100
rect 42797 21097 42809 21100
rect 42843 21128 42855 21131
rect 43530 21128 43536 21140
rect 42843 21100 43536 21128
rect 42843 21097 42855 21100
rect 42797 21091 42855 21097
rect 43530 21088 43536 21100
rect 43588 21088 43594 21140
rect 43806 21088 43812 21140
rect 43864 21128 43870 21140
rect 44085 21131 44143 21137
rect 44085 21128 44097 21131
rect 43864 21100 44097 21128
rect 43864 21088 43870 21100
rect 44085 21097 44097 21100
rect 44131 21097 44143 21131
rect 44085 21091 44143 21097
rect 44450 21088 44456 21140
rect 44508 21088 44514 21140
rect 45186 21088 45192 21140
rect 45244 21088 45250 21140
rect 45830 21088 45836 21140
rect 45888 21088 45894 21140
rect 40862 21020 40868 21072
rect 40920 21060 40926 21072
rect 42613 21063 42671 21069
rect 42613 21060 42625 21063
rect 40920 21032 42625 21060
rect 40920 21020 40926 21032
rect 42613 21029 42625 21032
rect 42659 21029 42671 21063
rect 42613 21023 42671 21029
rect 41785 20995 41843 21001
rect 41785 20992 41797 20995
rect 40788 20964 41797 20992
rect 41785 20961 41797 20964
rect 41831 20961 41843 20995
rect 41785 20955 41843 20961
rect 42426 20952 42432 21004
rect 42484 20952 42490 21004
rect 42628 20992 42656 21023
rect 43346 21020 43352 21072
rect 43404 21060 43410 21072
rect 43901 21063 43959 21069
rect 43901 21060 43913 21063
rect 43404 21032 43913 21060
rect 43404 21020 43410 21032
rect 43901 21029 43913 21032
rect 43947 21029 43959 21063
rect 43901 21023 43959 21029
rect 44358 21020 44364 21072
rect 44416 21060 44422 21072
rect 44729 21063 44787 21069
rect 44729 21060 44741 21063
rect 44416 21032 44741 21060
rect 44416 21020 44422 21032
rect 44729 21029 44741 21032
rect 44775 21060 44787 21063
rect 45370 21060 45376 21072
rect 44775 21032 45376 21060
rect 44775 21029 44787 21032
rect 44729 21023 44787 21029
rect 45370 21020 45376 21032
rect 45428 21020 45434 21072
rect 46569 21063 46627 21069
rect 46569 21060 46581 21063
rect 45526 21032 46581 21060
rect 45526 20992 45554 21032
rect 46569 21029 46581 21032
rect 46615 21029 46627 21063
rect 46842 21060 46848 21072
rect 46569 21023 46627 21029
rect 46676 21032 46848 21060
rect 42628 20964 45554 20992
rect 43441 20927 43499 20933
rect 43441 20924 43453 20927
rect 40696 20896 43453 20924
rect 40497 20887 40555 20893
rect 43441 20893 43453 20896
rect 43487 20924 43499 20927
rect 43717 20927 43775 20933
rect 43717 20924 43729 20927
rect 43487 20896 43729 20924
rect 43487 20893 43499 20896
rect 43441 20887 43499 20893
rect 43717 20893 43729 20896
rect 43763 20893 43775 20927
rect 43717 20887 43775 20893
rect 45370 20884 45376 20936
rect 45428 20884 45434 20936
rect 46017 20927 46075 20933
rect 46017 20893 46029 20927
rect 46063 20924 46075 20927
rect 46676 20924 46704 21032
rect 46842 21020 46848 21032
rect 46900 21020 46906 21072
rect 48314 20992 48320 21004
rect 46768 20964 48320 20992
rect 46768 20933 46796 20964
rect 48314 20952 48320 20964
rect 48372 20952 48378 21004
rect 46063 20896 46704 20924
rect 46753 20927 46811 20933
rect 46063 20893 46075 20896
rect 46017 20887 46075 20893
rect 46753 20893 46765 20927
rect 46799 20893 46811 20927
rect 46753 20887 46811 20893
rect 47489 20927 47547 20933
rect 47489 20893 47501 20927
rect 47535 20924 47547 20927
rect 47854 20924 47860 20936
rect 47535 20896 47860 20924
rect 47535 20893 47547 20896
rect 47489 20887 47547 20893
rect 47854 20884 47860 20896
rect 47912 20884 47918 20936
rect 48225 20927 48283 20933
rect 48225 20893 48237 20927
rect 48271 20924 48283 20927
rect 48685 20927 48743 20933
rect 48685 20924 48697 20927
rect 48271 20896 48697 20924
rect 48271 20893 48283 20896
rect 48225 20887 48283 20893
rect 48685 20893 48697 20896
rect 48731 20893 48743 20927
rect 48685 20887 48743 20893
rect 49326 20884 49332 20936
rect 49384 20884 49390 20936
rect 40126 20856 40132 20868
rect 40052 20828 40132 20856
rect 40052 20797 40080 20828
rect 40126 20816 40132 20828
rect 40184 20816 40190 20868
rect 40405 20859 40463 20865
rect 40405 20825 40417 20859
rect 40451 20856 40463 20859
rect 41601 20859 41659 20865
rect 40451 20828 41276 20856
rect 40451 20825 40463 20828
rect 40405 20819 40463 20825
rect 41248 20797 41276 20828
rect 41601 20825 41613 20859
rect 41647 20856 41659 20859
rect 44174 20856 44180 20868
rect 41647 20828 44180 20856
rect 41647 20825 41659 20828
rect 41601 20819 41659 20825
rect 44174 20816 44180 20828
rect 44232 20816 44238 20868
rect 44637 20859 44695 20865
rect 44637 20825 44649 20859
rect 44683 20856 44695 20859
rect 49344 20856 49372 20884
rect 44683 20828 49372 20856
rect 44683 20825 44695 20828
rect 44637 20819 44695 20825
rect 38804 20760 39896 20788
rect 40037 20791 40095 20797
rect 38804 20748 38810 20760
rect 40037 20757 40049 20791
rect 40083 20757 40095 20791
rect 40037 20751 40095 20757
rect 41233 20791 41291 20797
rect 41233 20757 41245 20791
rect 41279 20757 41291 20791
rect 41233 20751 41291 20757
rect 41322 20748 41328 20800
rect 41380 20788 41386 20800
rect 41693 20791 41751 20797
rect 41693 20788 41705 20791
rect 41380 20760 41705 20788
rect 41380 20748 41386 20760
rect 41693 20757 41705 20760
rect 41739 20788 41751 20791
rect 42245 20791 42303 20797
rect 42245 20788 42257 20791
rect 41739 20760 42257 20788
rect 41739 20757 41751 20760
rect 41693 20751 41751 20757
rect 42245 20757 42257 20760
rect 42291 20757 42303 20791
rect 42245 20751 42303 20757
rect 43257 20791 43315 20797
rect 43257 20757 43269 20791
rect 43303 20788 43315 20791
rect 43346 20788 43352 20800
rect 43303 20760 43352 20788
rect 43303 20757 43315 20760
rect 43257 20751 43315 20757
rect 43346 20748 43352 20760
rect 43404 20748 43410 20800
rect 47302 20748 47308 20800
rect 47360 20748 47366 20800
rect 47394 20748 47400 20800
rect 47452 20788 47458 20800
rect 48041 20791 48099 20797
rect 48041 20788 48053 20791
rect 47452 20760 48053 20788
rect 47452 20748 47458 20760
rect 48041 20757 48053 20760
rect 48087 20757 48099 20791
rect 48041 20751 48099 20757
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5445 20587 5503 20593
rect 5445 20553 5457 20587
rect 5491 20584 5503 20587
rect 6546 20584 6552 20596
rect 5491 20556 6552 20584
rect 5491 20553 5503 20556
rect 5445 20547 5503 20553
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 14093 20587 14151 20593
rect 14093 20584 14105 20587
rect 11112 20556 14105 20584
rect 11112 20544 11118 20556
rect 14093 20553 14105 20556
rect 14139 20553 14151 20587
rect 14093 20547 14151 20553
rect 14921 20587 14979 20593
rect 14921 20553 14933 20587
rect 14967 20553 14979 20587
rect 14921 20547 14979 20553
rect 1302 20476 1308 20528
rect 1360 20516 1366 20528
rect 3605 20519 3663 20525
rect 3605 20516 3617 20519
rect 1360 20488 3617 20516
rect 1360 20476 1366 20488
rect 3605 20485 3617 20488
rect 3651 20485 3663 20519
rect 8294 20516 8300 20528
rect 3605 20479 3663 20485
rect 5276 20488 8300 20516
rect 5276 20457 5304 20488
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 11149 20519 11207 20525
rect 11149 20485 11161 20519
rect 11195 20516 11207 20519
rect 13538 20516 13544 20528
rect 11195 20488 13544 20516
rect 11195 20485 11207 20488
rect 11149 20479 11207 20485
rect 13538 20476 13544 20488
rect 13596 20476 13602 20528
rect 13630 20476 13636 20528
rect 13688 20516 13694 20528
rect 14936 20516 14964 20547
rect 15562 20544 15568 20596
rect 15620 20544 15626 20596
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15896 20556 15945 20584
rect 15896 20544 15902 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 16022 20544 16028 20596
rect 16080 20544 16086 20596
rect 17126 20544 17132 20596
rect 17184 20544 17190 20596
rect 18785 20587 18843 20593
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 18874 20584 18880 20596
rect 18831 20556 18880 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 19702 20544 19708 20596
rect 19760 20544 19766 20596
rect 19886 20544 19892 20596
rect 19944 20584 19950 20596
rect 19944 20556 22094 20584
rect 19944 20544 19950 20556
rect 16206 20516 16212 20528
rect 13688 20488 14964 20516
rect 15028 20488 16212 20516
rect 13688 20476 13694 20488
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 4801 20451 4859 20457
rect 3007 20420 4752 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 2547 20352 2774 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 2746 20324 2774 20352
rect 2746 20284 2780 20324
rect 2774 20272 2780 20284
rect 2832 20272 2838 20324
rect 4724 20312 4752 20420
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 5261 20451 5319 20457
rect 5261 20417 5273 20451
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 4816 20380 4844 20411
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6512 20420 6561 20448
rect 6512 20408 6518 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9766 20448 9772 20460
rect 9263 20420 9772 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10410 20448 10416 20460
rect 9907 20420 10416 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10410 20408 10416 20420
rect 10468 20408 10474 20460
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 11514 20448 11520 20460
rect 10551 20420 11520 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 11514 20408 11520 20420
rect 11572 20408 11578 20460
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11756 20420 11897 20448
rect 11756 20408 11762 20420
rect 11885 20417 11897 20420
rect 11931 20448 11943 20451
rect 12434 20448 12440 20460
rect 11931 20420 12440 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 12434 20408 12440 20420
rect 12492 20408 12498 20460
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20448 12679 20451
rect 12894 20448 12900 20460
rect 12667 20420 12900 20448
rect 12667 20417 12679 20420
rect 12621 20411 12679 20417
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20448 13139 20451
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 13127 20420 13277 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13265 20417 13277 20420
rect 13311 20448 13323 20451
rect 13354 20448 13360 20460
rect 13311 20420 13360 20448
rect 13311 20417 13323 20420
rect 13265 20411 13323 20417
rect 13354 20408 13360 20420
rect 13412 20448 13418 20460
rect 13722 20448 13728 20460
rect 13412 20420 13728 20448
rect 13412 20408 13418 20420
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 15028 20448 15056 20488
rect 16206 20476 16212 20488
rect 16264 20476 16270 20528
rect 17144 20516 17172 20544
rect 16960 20488 17172 20516
rect 22066 20516 22094 20556
rect 22278 20544 22284 20596
rect 22336 20584 22342 20596
rect 22922 20584 22928 20596
rect 22336 20556 22928 20584
rect 22336 20544 22342 20556
rect 22922 20544 22928 20556
rect 22980 20584 22986 20596
rect 25682 20584 25688 20596
rect 22980 20556 25688 20584
rect 22980 20544 22986 20556
rect 22373 20519 22431 20525
rect 22066 20488 22324 20516
rect 13872 20420 15056 20448
rect 13872 20408 13878 20420
rect 15102 20408 15108 20460
rect 15160 20408 15166 20460
rect 6362 20380 6368 20392
rect 4816 20352 6368 20380
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 6638 20340 6644 20392
rect 6696 20380 6702 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 6696 20352 7021 20380
rect 6696 20340 6702 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 8386 20340 8392 20392
rect 8444 20380 8450 20392
rect 11054 20380 11060 20392
rect 8444 20352 11060 20380
rect 8444 20340 8450 20352
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 14185 20383 14243 20389
rect 11204 20352 13768 20380
rect 11204 20340 11210 20352
rect 4724 20284 9168 20312
rect 4522 20204 4528 20256
rect 4580 20244 4586 20256
rect 9033 20247 9091 20253
rect 9033 20244 9045 20247
rect 4580 20216 9045 20244
rect 4580 20204 4586 20216
rect 9033 20213 9045 20216
rect 9079 20213 9091 20247
rect 9140 20244 9168 20284
rect 10134 20272 10140 20324
rect 10192 20312 10198 20324
rect 13740 20321 13768 20352
rect 14185 20349 14197 20383
rect 14231 20349 14243 20383
rect 14185 20343 14243 20349
rect 13725 20315 13783 20321
rect 10192 20284 13676 20312
rect 10192 20272 10198 20284
rect 11054 20244 11060 20256
rect 9140 20216 11060 20244
rect 9033 20207 9091 20213
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11606 20204 11612 20256
rect 11664 20244 11670 20256
rect 11793 20247 11851 20253
rect 11793 20244 11805 20247
rect 11664 20216 11805 20244
rect 11664 20204 11670 20216
rect 11793 20213 11805 20216
rect 11839 20213 11851 20247
rect 11793 20207 11851 20213
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 12529 20247 12587 20253
rect 12529 20244 12541 20247
rect 11940 20216 12541 20244
rect 11940 20204 11946 20216
rect 12529 20213 12541 20216
rect 12575 20213 12587 20247
rect 12529 20207 12587 20213
rect 13446 20204 13452 20256
rect 13504 20204 13510 20256
rect 13648 20244 13676 20284
rect 13725 20281 13737 20315
rect 13771 20281 13783 20315
rect 14200 20312 14228 20343
rect 14274 20340 14280 20392
rect 14332 20340 14338 20392
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20380 16267 20383
rect 16960 20380 16988 20488
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 19061 20451 19119 20457
rect 19061 20448 19073 20451
rect 18446 20420 19073 20448
rect 19061 20417 19073 20420
rect 19107 20448 19119 20451
rect 19426 20448 19432 20460
rect 19107 20420 19432 20448
rect 19107 20417 19119 20420
rect 19061 20411 19119 20417
rect 19426 20408 19432 20420
rect 19484 20448 19490 20460
rect 21453 20451 21511 20457
rect 19484 20420 20102 20448
rect 19484 20408 19490 20420
rect 21453 20417 21465 20451
rect 21499 20448 21511 20451
rect 22094 20448 22100 20460
rect 21499 20420 22100 20448
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 22094 20408 22100 20420
rect 22152 20408 22158 20460
rect 22296 20448 22324 20488
rect 22373 20485 22385 20519
rect 22419 20516 22431 20519
rect 23658 20516 23664 20528
rect 22419 20488 23664 20516
rect 22419 20485 22431 20488
rect 22373 20479 22431 20485
rect 23658 20476 23664 20488
rect 23716 20476 23722 20528
rect 23385 20451 23443 20457
rect 22296 20420 23336 20448
rect 16255 20352 16988 20380
rect 17313 20383 17371 20389
rect 16255 20349 16267 20352
rect 16209 20343 16267 20349
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17402 20380 17408 20392
rect 17359 20352 17408 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 17402 20340 17408 20352
rect 17460 20380 17466 20392
rect 20438 20380 20444 20392
rect 17460 20352 20444 20380
rect 17460 20340 17466 20352
rect 20438 20340 20444 20352
rect 20496 20340 20502 20392
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21542 20380 21548 20392
rect 21223 20352 21548 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 21542 20340 21548 20352
rect 21600 20340 21606 20392
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20349 22523 20383
rect 22465 20343 22523 20349
rect 16850 20312 16856 20324
rect 14200 20284 16856 20312
rect 13725 20275 13783 20281
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 20070 20312 20076 20324
rect 18340 20284 20076 20312
rect 16482 20244 16488 20256
rect 13648 20216 16488 20244
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 16761 20247 16819 20253
rect 16761 20213 16773 20247
rect 16807 20244 16819 20247
rect 17126 20244 17132 20256
rect 16807 20216 17132 20244
rect 16807 20213 16819 20216
rect 16761 20207 16819 20213
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 17310 20204 17316 20256
rect 17368 20244 17374 20256
rect 18340 20244 18368 20284
rect 20070 20272 20076 20284
rect 20128 20272 20134 20324
rect 17368 20216 18368 20244
rect 19337 20247 19395 20253
rect 17368 20204 17374 20216
rect 19337 20213 19349 20247
rect 19383 20244 19395 20247
rect 19610 20244 19616 20256
rect 19383 20216 19616 20244
rect 19383 20213 19395 20216
rect 19337 20207 19395 20213
rect 19610 20204 19616 20216
rect 19668 20204 19674 20256
rect 19978 20204 19984 20256
rect 20036 20244 20042 20256
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 20036 20216 22017 20244
rect 20036 20204 20042 20216
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22480 20244 22508 20343
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 23308 20380 23336 20420
rect 23385 20417 23397 20451
rect 23431 20448 23443 20451
rect 23750 20448 23756 20460
rect 23431 20420 23756 20448
rect 23431 20417 23443 20420
rect 23385 20411 23443 20417
rect 23750 20408 23756 20420
rect 23808 20408 23814 20460
rect 23860 20457 23888 20556
rect 25682 20544 25688 20556
rect 25740 20544 25746 20596
rect 30834 20584 30840 20596
rect 27264 20556 30840 20584
rect 24026 20476 24032 20528
rect 24084 20516 24090 20528
rect 24121 20519 24179 20525
rect 24121 20516 24133 20519
rect 24084 20488 24133 20516
rect 24084 20476 24090 20488
rect 24121 20485 24133 20488
rect 24167 20516 24179 20519
rect 24210 20516 24216 20528
rect 24167 20488 24216 20516
rect 24167 20485 24179 20488
rect 24121 20479 24179 20485
rect 24210 20476 24216 20488
rect 24268 20476 24274 20528
rect 24578 20476 24584 20528
rect 24636 20476 24642 20528
rect 25866 20476 25872 20528
rect 25924 20516 25930 20528
rect 25924 20488 26188 20516
rect 25924 20476 25930 20488
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 25958 20408 25964 20460
rect 26016 20448 26022 20460
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 26016 20420 26065 20448
rect 26016 20408 26022 20420
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 23308 20352 25176 20380
rect 22738 20272 22744 20324
rect 22796 20312 22802 20324
rect 23201 20315 23259 20321
rect 23201 20312 23213 20315
rect 22796 20284 23213 20312
rect 22796 20272 22802 20284
rect 23201 20281 23213 20284
rect 23247 20281 23259 20315
rect 25148 20312 25176 20352
rect 25590 20340 25596 20392
rect 25648 20340 25654 20392
rect 26160 20380 26188 20488
rect 27264 20457 27292 20556
rect 30834 20544 30840 20556
rect 30892 20584 30898 20596
rect 31478 20584 31484 20596
rect 30892 20556 31484 20584
rect 30892 20544 30898 20556
rect 31478 20544 31484 20556
rect 31536 20584 31542 20596
rect 32490 20584 32496 20596
rect 31536 20556 32496 20584
rect 31536 20544 31542 20556
rect 32490 20544 32496 20556
rect 32548 20584 32554 20596
rect 35253 20587 35311 20593
rect 32548 20556 34100 20584
rect 32548 20544 32554 20556
rect 28258 20476 28264 20528
rect 28316 20476 28322 20528
rect 29638 20476 29644 20528
rect 29696 20516 29702 20528
rect 29733 20519 29791 20525
rect 29733 20516 29745 20519
rect 29696 20488 29745 20516
rect 29696 20476 29702 20488
rect 29733 20485 29745 20488
rect 29779 20516 29791 20519
rect 31021 20519 31079 20525
rect 29779 20488 30604 20516
rect 29779 20485 29791 20488
rect 29733 20479 29791 20485
rect 27249 20451 27307 20457
rect 27249 20417 27261 20451
rect 27295 20417 27307 20451
rect 29825 20451 29883 20457
rect 29825 20448 29837 20451
rect 27249 20411 27307 20417
rect 28736 20420 29837 20448
rect 27525 20383 27583 20389
rect 27525 20380 27537 20383
rect 26160 20352 27537 20380
rect 27525 20349 27537 20352
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 28534 20340 28540 20392
rect 28592 20380 28598 20392
rect 28736 20380 28764 20420
rect 29825 20417 29837 20420
rect 29871 20417 29883 20451
rect 29825 20411 29883 20417
rect 28592 20352 28764 20380
rect 28592 20340 28598 20352
rect 29086 20340 29092 20392
rect 29144 20380 29150 20392
rect 29454 20380 29460 20392
rect 29144 20352 29460 20380
rect 29144 20340 29150 20352
rect 29454 20340 29460 20352
rect 29512 20380 29518 20392
rect 29549 20383 29607 20389
rect 29549 20380 29561 20383
rect 29512 20352 29561 20380
rect 29512 20340 29518 20352
rect 29549 20349 29561 20352
rect 29595 20380 29607 20383
rect 30098 20380 30104 20392
rect 29595 20352 30104 20380
rect 29595 20349 29607 20352
rect 29549 20343 29607 20349
rect 30098 20340 30104 20352
rect 30156 20340 30162 20392
rect 26050 20312 26056 20324
rect 25148 20284 26056 20312
rect 23201 20275 23259 20281
rect 26050 20272 26056 20284
rect 26108 20272 26114 20324
rect 26142 20272 26148 20324
rect 26200 20312 26206 20324
rect 26605 20315 26663 20321
rect 26605 20312 26617 20315
rect 26200 20284 26617 20312
rect 26200 20272 26206 20284
rect 26605 20281 26617 20284
rect 26651 20281 26663 20315
rect 26605 20275 26663 20281
rect 28997 20315 29055 20321
rect 28997 20281 29009 20315
rect 29043 20312 29055 20315
rect 29362 20312 29368 20324
rect 29043 20284 29368 20312
rect 29043 20281 29055 20284
rect 28997 20275 29055 20281
rect 29362 20272 29368 20284
rect 29420 20272 29426 20324
rect 30282 20312 30288 20324
rect 30024 20284 30288 20312
rect 25498 20244 25504 20256
rect 22480 20216 25504 20244
rect 22005 20207 22063 20213
rect 25498 20204 25504 20216
rect 25556 20204 25562 20256
rect 26237 20247 26295 20253
rect 26237 20213 26249 20247
rect 26283 20244 26295 20247
rect 26418 20244 26424 20256
rect 26283 20216 26424 20244
rect 26283 20213 26295 20216
rect 26237 20207 26295 20213
rect 26418 20204 26424 20216
rect 26476 20204 26482 20256
rect 27338 20204 27344 20256
rect 27396 20244 27402 20256
rect 30024 20244 30052 20284
rect 30282 20272 30288 20284
rect 30340 20272 30346 20324
rect 30576 20312 30604 20488
rect 31021 20485 31033 20519
rect 31067 20516 31079 20519
rect 31570 20516 31576 20528
rect 31067 20488 31576 20516
rect 31067 20485 31079 20488
rect 31021 20479 31079 20485
rect 31570 20476 31576 20488
rect 31628 20476 31634 20528
rect 31662 20476 31668 20528
rect 31720 20516 31726 20528
rect 31720 20488 31984 20516
rect 31720 20476 31726 20488
rect 31113 20451 31171 20457
rect 31113 20417 31125 20451
rect 31159 20448 31171 20451
rect 31159 20420 31754 20448
rect 31159 20417 31171 20420
rect 31113 20411 31171 20417
rect 30650 20340 30656 20392
rect 30708 20380 30714 20392
rect 31205 20383 31263 20389
rect 31205 20380 31217 20383
rect 30708 20352 31217 20380
rect 30708 20340 30714 20352
rect 31205 20349 31217 20352
rect 31251 20349 31263 20383
rect 31726 20380 31754 20420
rect 31956 20392 31984 20488
rect 32214 20476 32220 20528
rect 32272 20516 32278 20528
rect 32272 20488 32614 20516
rect 32272 20476 32278 20488
rect 31846 20380 31852 20392
rect 31726 20352 31852 20380
rect 31205 20343 31263 20349
rect 31846 20340 31852 20352
rect 31904 20340 31910 20392
rect 31938 20340 31944 20392
rect 31996 20340 32002 20392
rect 32306 20340 32312 20392
rect 32364 20340 32370 20392
rect 32582 20340 32588 20392
rect 32640 20380 32646 20392
rect 33410 20380 33416 20392
rect 32640 20352 33416 20380
rect 32640 20340 32646 20352
rect 33410 20340 33416 20352
rect 33468 20340 33474 20392
rect 33686 20340 33692 20392
rect 33744 20380 33750 20392
rect 34072 20389 34100 20556
rect 35253 20553 35265 20587
rect 35299 20584 35311 20587
rect 36170 20584 36176 20596
rect 35299 20556 36176 20584
rect 35299 20553 35311 20556
rect 35253 20547 35311 20553
rect 36170 20544 36176 20556
rect 36228 20544 36234 20596
rect 36906 20584 36912 20596
rect 36372 20556 36912 20584
rect 35894 20516 35900 20528
rect 34716 20488 35900 20516
rect 33781 20383 33839 20389
rect 33781 20380 33793 20383
rect 33744 20352 33793 20380
rect 33744 20340 33750 20352
rect 33781 20349 33793 20352
rect 33827 20349 33839 20383
rect 33781 20343 33839 20349
rect 34057 20383 34115 20389
rect 34057 20349 34069 20383
rect 34103 20380 34115 20383
rect 34514 20380 34520 20392
rect 34103 20352 34520 20380
rect 34103 20349 34115 20352
rect 34057 20343 34115 20349
rect 34514 20340 34520 20352
rect 34572 20340 34578 20392
rect 34716 20389 34744 20488
rect 35894 20476 35900 20488
rect 35952 20476 35958 20528
rect 34882 20408 34888 20460
rect 34940 20448 34946 20460
rect 36372 20448 36400 20556
rect 36906 20544 36912 20556
rect 36964 20544 36970 20596
rect 37090 20544 37096 20596
rect 37148 20584 37154 20596
rect 40221 20587 40279 20593
rect 37148 20556 38884 20584
rect 37148 20544 37154 20556
rect 36541 20519 36599 20525
rect 36541 20485 36553 20519
rect 36587 20516 36599 20519
rect 37182 20516 37188 20528
rect 36587 20488 37188 20516
rect 36587 20485 36599 20488
rect 36541 20479 36599 20485
rect 37182 20476 37188 20488
rect 37240 20476 37246 20528
rect 37734 20476 37740 20528
rect 37792 20516 37798 20528
rect 37918 20516 37924 20528
rect 37792 20488 37924 20516
rect 37792 20476 37798 20488
rect 37918 20476 37924 20488
rect 37976 20516 37982 20528
rect 38856 20516 38884 20556
rect 40221 20553 40233 20587
rect 40267 20584 40279 20587
rect 41785 20587 41843 20593
rect 41785 20584 41797 20587
rect 40267 20556 41797 20584
rect 40267 20553 40279 20556
rect 40221 20547 40279 20553
rect 41785 20553 41797 20556
rect 41831 20584 41843 20587
rect 43622 20584 43628 20596
rect 41831 20556 43628 20584
rect 41831 20553 41843 20556
rect 41785 20547 41843 20553
rect 43622 20544 43628 20556
rect 43680 20544 43686 20596
rect 43898 20544 43904 20596
rect 43956 20584 43962 20596
rect 45189 20587 45247 20593
rect 45189 20584 45201 20587
rect 43956 20556 45201 20584
rect 43956 20544 43962 20556
rect 45189 20553 45201 20556
rect 45235 20553 45247 20587
rect 45189 20547 45247 20553
rect 46198 20544 46204 20596
rect 46256 20584 46262 20596
rect 46293 20587 46351 20593
rect 46293 20584 46305 20587
rect 46256 20556 46305 20584
rect 46256 20544 46262 20556
rect 46293 20553 46305 20556
rect 46339 20553 46351 20587
rect 46293 20547 46351 20553
rect 46474 20544 46480 20596
rect 46532 20544 46538 20596
rect 46842 20544 46848 20596
rect 46900 20584 46906 20596
rect 47670 20584 47676 20596
rect 46900 20556 47676 20584
rect 46900 20544 46906 20556
rect 47670 20544 47676 20556
rect 47728 20544 47734 20596
rect 41141 20519 41199 20525
rect 41141 20516 41153 20519
rect 37976 20488 38042 20516
rect 38856 20488 41153 20516
rect 37976 20476 37982 20488
rect 41141 20485 41153 20488
rect 41187 20485 41199 20519
rect 47949 20519 48007 20525
rect 47949 20516 47961 20519
rect 41141 20479 41199 20485
rect 41616 20488 47961 20516
rect 34940 20420 36400 20448
rect 36449 20451 36507 20457
rect 34940 20408 34946 20420
rect 36449 20417 36461 20451
rect 36495 20448 36507 20451
rect 37458 20448 37464 20460
rect 36495 20420 37464 20448
rect 36495 20417 36507 20420
rect 36449 20411 36507 20417
rect 37458 20408 37464 20420
rect 37516 20408 37522 20460
rect 39482 20408 39488 20460
rect 39540 20408 39546 20460
rect 39758 20408 39764 20460
rect 39816 20448 39822 20460
rect 41616 20457 41644 20488
rect 47949 20485 47961 20488
rect 47995 20485 48007 20519
rect 47949 20479 48007 20485
rect 40313 20451 40371 20457
rect 40313 20448 40325 20451
rect 39816 20420 40325 20448
rect 39816 20408 39822 20420
rect 40313 20417 40325 20420
rect 40359 20448 40371 20451
rect 41601 20451 41659 20457
rect 41601 20448 41613 20451
rect 40359 20420 41613 20448
rect 40359 20417 40371 20420
rect 40313 20411 40371 20417
rect 41601 20417 41613 20420
rect 41647 20417 41659 20451
rect 41601 20411 41659 20417
rect 45373 20451 45431 20457
rect 45373 20417 45385 20451
rect 45419 20448 45431 20451
rect 46017 20451 46075 20457
rect 45419 20420 45554 20448
rect 45419 20417 45431 20420
rect 45373 20411 45431 20417
rect 34701 20383 34759 20389
rect 34701 20349 34713 20383
rect 34747 20349 34759 20383
rect 34701 20343 34759 20349
rect 34790 20340 34796 20392
rect 34848 20340 34854 20392
rect 35066 20340 35072 20392
rect 35124 20380 35130 20392
rect 35713 20383 35771 20389
rect 35713 20380 35725 20383
rect 35124 20352 35725 20380
rect 35124 20340 35130 20352
rect 35713 20349 35725 20352
rect 35759 20349 35771 20383
rect 35713 20343 35771 20349
rect 36725 20383 36783 20389
rect 36725 20349 36737 20383
rect 36771 20380 36783 20383
rect 37274 20380 37280 20392
rect 36771 20352 37280 20380
rect 36771 20349 36783 20352
rect 36725 20343 36783 20349
rect 37274 20340 37280 20352
rect 37332 20340 37338 20392
rect 37642 20340 37648 20392
rect 37700 20380 37706 20392
rect 39209 20383 39267 20389
rect 39209 20380 39221 20383
rect 37700 20352 39221 20380
rect 37700 20340 37706 20352
rect 39209 20349 39221 20352
rect 39255 20349 39267 20383
rect 39209 20343 39267 20349
rect 40126 20340 40132 20392
rect 40184 20340 40190 20392
rect 45526 20380 45554 20420
rect 46017 20417 46029 20451
rect 46063 20448 46075 20451
rect 46474 20448 46480 20460
rect 46063 20420 46480 20448
rect 46063 20417 46075 20420
rect 46017 20411 46075 20417
rect 46474 20408 46480 20420
rect 46532 20408 46538 20460
rect 47210 20408 47216 20460
rect 47268 20408 47274 20460
rect 48133 20451 48191 20457
rect 48133 20417 48145 20451
rect 48179 20448 48191 20451
rect 48685 20451 48743 20457
rect 48685 20448 48697 20451
rect 48179 20420 48697 20448
rect 48179 20417 48191 20420
rect 48133 20411 48191 20417
rect 48685 20417 48697 20420
rect 48731 20417 48743 20451
rect 48685 20411 48743 20417
rect 49326 20408 49332 20460
rect 49384 20408 49390 20460
rect 46198 20380 46204 20392
rect 45526 20352 46204 20380
rect 46198 20340 46204 20352
rect 46256 20340 46262 20392
rect 42794 20312 42800 20324
rect 30576 20284 30972 20312
rect 27396 20216 30052 20244
rect 30193 20247 30251 20253
rect 27396 20204 27402 20216
rect 30193 20213 30205 20247
rect 30239 20244 30251 20247
rect 30558 20244 30564 20256
rect 30239 20216 30564 20244
rect 30239 20213 30251 20216
rect 30193 20207 30251 20213
rect 30558 20204 30564 20216
rect 30616 20204 30622 20256
rect 30653 20247 30711 20253
rect 30653 20213 30665 20247
rect 30699 20244 30711 20247
rect 30834 20244 30840 20256
rect 30699 20216 30840 20244
rect 30699 20213 30711 20216
rect 30653 20207 30711 20213
rect 30834 20204 30840 20216
rect 30892 20204 30898 20256
rect 30944 20244 30972 20284
rect 33980 20284 37872 20312
rect 31757 20247 31815 20253
rect 31757 20244 31769 20247
rect 30944 20216 31769 20244
rect 31757 20213 31769 20216
rect 31803 20244 31815 20247
rect 33980 20244 34008 20284
rect 31803 20216 34008 20244
rect 31803 20213 31815 20216
rect 31757 20207 31815 20213
rect 35250 20204 35256 20256
rect 35308 20244 35314 20256
rect 35529 20247 35587 20253
rect 35529 20244 35541 20247
rect 35308 20216 35541 20244
rect 35308 20204 35314 20216
rect 35529 20213 35541 20216
rect 35575 20213 35587 20247
rect 35529 20207 35587 20213
rect 36078 20204 36084 20256
rect 36136 20204 36142 20256
rect 37369 20247 37427 20253
rect 37369 20213 37381 20247
rect 37415 20244 37427 20247
rect 37642 20244 37648 20256
rect 37415 20216 37648 20244
rect 37415 20213 37427 20216
rect 37369 20207 37427 20213
rect 37642 20204 37648 20216
rect 37700 20204 37706 20256
rect 37734 20204 37740 20256
rect 37792 20204 37798 20256
rect 37844 20244 37872 20284
rect 39408 20284 42800 20312
rect 39408 20244 39436 20284
rect 42794 20272 42800 20284
rect 42852 20272 42858 20324
rect 44913 20315 44971 20321
rect 44913 20281 44925 20315
rect 44959 20312 44971 20315
rect 49326 20312 49332 20324
rect 44959 20284 49332 20312
rect 44959 20281 44971 20284
rect 44913 20275 44971 20281
rect 49326 20272 49332 20284
rect 49384 20272 49390 20324
rect 37844 20216 39436 20244
rect 40678 20204 40684 20256
rect 40736 20204 40742 20256
rect 41138 20204 41144 20256
rect 41196 20244 41202 20256
rect 45833 20247 45891 20253
rect 45833 20244 45845 20247
rect 41196 20216 45845 20244
rect 41196 20204 41202 20216
rect 45833 20213 45845 20216
rect 45879 20213 45891 20247
rect 45833 20207 45891 20213
rect 47026 20204 47032 20256
rect 47084 20204 47090 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 5276 20012 13768 20040
rect 4246 19864 4252 19916
rect 4304 19864 4310 19916
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 5276 19836 5304 20012
rect 6362 19932 6368 19984
rect 6420 19972 6426 19984
rect 11241 19975 11299 19981
rect 11241 19972 11253 19975
rect 6420 19944 11253 19972
rect 6420 19932 6426 19944
rect 11241 19941 11253 19944
rect 11287 19941 11299 19975
rect 13740 19972 13768 20012
rect 14458 20000 14464 20052
rect 14516 20000 14522 20052
rect 15010 20000 15016 20052
rect 15068 20040 15074 20052
rect 15068 20012 15792 20040
rect 15068 20000 15074 20012
rect 14921 19975 14979 19981
rect 14921 19972 14933 19975
rect 13740 19944 14933 19972
rect 11241 19935 11299 19941
rect 14921 19941 14933 19944
rect 14967 19941 14979 19975
rect 15764 19972 15792 20012
rect 16482 20000 16488 20052
rect 16540 20040 16546 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16540 20012 16865 20040
rect 16540 20000 16546 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 18322 20040 18328 20052
rect 18187 20012 18328 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 19337 20043 19395 20049
rect 19337 20040 19349 20043
rect 18472 20012 19349 20040
rect 18472 20000 18478 20012
rect 19337 20009 19349 20012
rect 19383 20040 19395 20043
rect 19886 20040 19892 20052
rect 19383 20012 19892 20040
rect 19383 20009 19395 20012
rect 19337 20003 19395 20009
rect 19886 20000 19892 20012
rect 19944 20000 19950 20052
rect 20070 20000 20076 20052
rect 20128 20040 20134 20052
rect 20257 20043 20315 20049
rect 20257 20040 20269 20043
rect 20128 20012 20269 20040
rect 20128 20000 20134 20012
rect 20257 20009 20269 20012
rect 20303 20040 20315 20043
rect 24029 20043 24087 20049
rect 20303 20012 22692 20040
rect 20303 20009 20315 20012
rect 20257 20003 20315 20009
rect 17310 19972 17316 19984
rect 15764 19944 17316 19972
rect 14921 19935 14979 19941
rect 17310 19932 17316 19944
rect 17368 19932 17374 19984
rect 18874 19972 18880 19984
rect 17512 19944 18880 19972
rect 5718 19864 5724 19916
rect 5776 19904 5782 19916
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5776 19876 6009 19904
rect 5776 19864 5782 19876
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 10962 19904 10968 19916
rect 5997 19867 6055 19873
rect 7944 19876 10968 19904
rect 3007 19808 5304 19836
rect 5353 19839 5411 19845
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 5353 19805 5365 19839
rect 5399 19836 5411 19839
rect 5442 19836 5448 19848
rect 5399 19808 5448 19836
rect 5399 19805 5411 19808
rect 5353 19799 5411 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 7944 19845 7972 19876
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19904 12035 19907
rect 12342 19904 12348 19916
rect 12023 19876 12348 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 13446 19864 13452 19916
rect 13504 19864 13510 19916
rect 16298 19864 16304 19916
rect 16356 19864 16362 19916
rect 17512 19913 17540 19944
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19873 17555 19907
rect 18785 19907 18843 19913
rect 17497 19867 17555 19873
rect 18432 19876 18736 19904
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 1486 19728 1492 19780
rect 1544 19768 1550 19780
rect 1765 19771 1823 19777
rect 1765 19768 1777 19771
rect 1544 19740 1777 19768
rect 1544 19728 1550 19740
rect 1765 19737 1777 19740
rect 1811 19737 1823 19771
rect 1765 19731 1823 19737
rect 7208 19700 7236 19799
rect 10134 19796 10140 19848
rect 10192 19796 10198 19848
rect 10778 19796 10784 19848
rect 10836 19796 10842 19848
rect 13354 19796 13360 19848
rect 13412 19796 13418 19848
rect 13464 19836 13492 19864
rect 14277 19839 14335 19845
rect 13464 19808 13584 19836
rect 9677 19771 9735 19777
rect 9677 19737 9689 19771
rect 9723 19768 9735 19771
rect 11422 19768 11428 19780
rect 9723 19740 11428 19768
rect 9723 19737 9735 19740
rect 9677 19731 9735 19737
rect 11422 19728 11428 19740
rect 11480 19728 11486 19780
rect 11698 19728 11704 19780
rect 11756 19768 11762 19780
rect 12253 19771 12311 19777
rect 12253 19768 12265 19771
rect 11756 19740 12265 19768
rect 11756 19728 11762 19740
rect 12253 19737 12265 19740
rect 12299 19737 12311 19771
rect 13556 19768 13584 19808
rect 14277 19805 14289 19839
rect 14323 19836 14335 19839
rect 16117 19839 16175 19845
rect 14323 19808 15976 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 15105 19771 15163 19777
rect 15105 19768 15117 19771
rect 13556 19740 15117 19768
rect 12253 19731 12311 19737
rect 15105 19737 15117 19740
rect 15151 19768 15163 19771
rect 15194 19768 15200 19780
rect 15151 19740 15200 19768
rect 15151 19737 15163 19740
rect 15105 19731 15163 19737
rect 15194 19728 15200 19740
rect 15252 19728 15258 19780
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7208 19672 7757 19700
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 9950 19660 9956 19712
rect 10008 19660 10014 19712
rect 10594 19660 10600 19712
rect 10652 19700 10658 19712
rect 10778 19700 10784 19712
rect 10652 19672 10784 19700
rect 10652 19660 10658 19672
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 13725 19703 13783 19709
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 15470 19700 15476 19712
rect 13771 19672 15476 19700
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 15470 19660 15476 19672
rect 15528 19660 15534 19712
rect 15654 19660 15660 19712
rect 15712 19660 15718 19712
rect 15948 19700 15976 19808
rect 16117 19805 16129 19839
rect 16163 19836 16175 19839
rect 18432 19836 18460 19876
rect 16163 19808 18460 19836
rect 18509 19839 18567 19845
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 18509 19805 18521 19839
rect 18555 19836 18567 19839
rect 18598 19836 18604 19848
rect 18555 19808 18604 19836
rect 18555 19805 18567 19808
rect 18509 19799 18567 19805
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 18708 19836 18736 19876
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 19334 19904 19340 19916
rect 18831 19876 19340 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 21450 19904 21456 19916
rect 19628 19876 21456 19904
rect 19628 19836 19656 19876
rect 21450 19864 21456 19876
rect 21508 19864 21514 19916
rect 22278 19864 22284 19916
rect 22336 19864 22342 19916
rect 20714 19836 20720 19848
rect 18708 19808 19656 19836
rect 19720 19808 20720 19836
rect 16025 19771 16083 19777
rect 16025 19737 16037 19771
rect 16071 19768 16083 19771
rect 16482 19768 16488 19780
rect 16071 19740 16488 19768
rect 16071 19737 16083 19740
rect 16025 19731 16083 19737
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 17678 19768 17684 19780
rect 17144 19740 17684 19768
rect 17144 19700 17172 19740
rect 17678 19728 17684 19740
rect 17736 19728 17742 19780
rect 19720 19768 19748 19808
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 20898 19796 20904 19848
rect 20956 19796 20962 19848
rect 22664 19836 22692 20012
rect 24029 20009 24041 20043
rect 24075 20040 24087 20043
rect 24946 20040 24952 20052
rect 24075 20012 24952 20040
rect 24075 20009 24087 20012
rect 24029 20003 24087 20009
rect 24946 20000 24952 20012
rect 25004 20000 25010 20052
rect 25038 20000 25044 20052
rect 25096 20040 25102 20052
rect 25222 20040 25228 20052
rect 25096 20012 25228 20040
rect 25096 20000 25102 20012
rect 25222 20000 25228 20012
rect 25280 20000 25286 20052
rect 25498 20000 25504 20052
rect 25556 20040 25562 20052
rect 25593 20043 25651 20049
rect 25593 20040 25605 20043
rect 25556 20012 25605 20040
rect 25556 20000 25562 20012
rect 25593 20009 25605 20012
rect 25639 20009 25651 20043
rect 25958 20040 25964 20052
rect 25593 20003 25651 20009
rect 25884 20012 25964 20040
rect 22741 19975 22799 19981
rect 22741 19941 22753 19975
rect 22787 19972 22799 19975
rect 25133 19975 25191 19981
rect 22787 19944 23520 19972
rect 22787 19941 22799 19944
rect 22741 19935 22799 19941
rect 23492 19913 23520 19944
rect 25133 19941 25145 19975
rect 25179 19972 25191 19975
rect 25884 19972 25912 20012
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 26050 20000 26056 20052
rect 26108 20040 26114 20052
rect 28534 20040 28540 20052
rect 26108 20012 28540 20040
rect 26108 20000 26114 20012
rect 28534 20000 28540 20012
rect 28592 20000 28598 20052
rect 30926 20040 30932 20052
rect 29012 20012 30932 20040
rect 27798 19972 27804 19984
rect 25179 19944 25912 19972
rect 25976 19944 27804 19972
rect 25179 19941 25191 19944
rect 25133 19935 25191 19941
rect 23477 19907 23535 19913
rect 23477 19873 23489 19907
rect 23523 19904 23535 19907
rect 23523 19876 23888 19904
rect 23523 19873 23535 19876
rect 23477 19867 23535 19873
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 22664 19808 23673 19836
rect 23661 19805 23673 19808
rect 23707 19805 23719 19839
rect 23860 19836 23888 19876
rect 23934 19864 23940 19916
rect 23992 19904 23998 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 23992 19876 24593 19904
rect 23992 19864 23998 19876
rect 24581 19873 24593 19876
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 25498 19836 25504 19848
rect 23860 19808 25504 19836
rect 23661 19799 23719 19805
rect 25498 19796 25504 19808
rect 25556 19796 25562 19848
rect 25976 19845 26004 19944
rect 27798 19932 27804 19944
rect 27856 19972 27862 19984
rect 28626 19972 28632 19984
rect 27856 19944 28632 19972
rect 27856 19932 27862 19944
rect 28626 19932 28632 19944
rect 28684 19932 28690 19984
rect 26050 19864 26056 19916
rect 26108 19864 26114 19916
rect 26237 19907 26295 19913
rect 26237 19873 26249 19907
rect 26283 19873 26295 19907
rect 27338 19904 27344 19916
rect 26237 19867 26295 19873
rect 26344 19876 27344 19904
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19805 26019 19839
rect 25961 19799 26019 19805
rect 18616 19740 19748 19768
rect 19797 19771 19855 19777
rect 15948 19672 17172 19700
rect 17218 19660 17224 19712
rect 17276 19660 17282 19712
rect 17310 19660 17316 19712
rect 17368 19660 17374 19712
rect 18616 19709 18644 19740
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 20622 19768 20628 19780
rect 19843 19740 20628 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 20622 19728 20628 19740
rect 20680 19728 20686 19780
rect 22005 19771 22063 19777
rect 22005 19737 22017 19771
rect 22051 19768 22063 19771
rect 22278 19768 22284 19780
rect 22051 19740 22284 19768
rect 22051 19737 22063 19740
rect 22005 19731 22063 19737
rect 22278 19728 22284 19740
rect 22336 19728 22342 19780
rect 25314 19768 25320 19780
rect 22572 19740 25320 19768
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19669 18659 19703
rect 18601 19663 18659 19669
rect 19518 19660 19524 19712
rect 19576 19700 19582 19712
rect 19705 19703 19763 19709
rect 19705 19700 19717 19703
rect 19576 19672 19717 19700
rect 19576 19660 19582 19672
rect 19705 19669 19717 19672
rect 19751 19669 19763 19703
rect 19705 19663 19763 19669
rect 20438 19660 20444 19712
rect 20496 19700 20502 19712
rect 20533 19703 20591 19709
rect 20533 19700 20545 19703
rect 20496 19672 20545 19700
rect 20496 19660 20502 19672
rect 20533 19669 20545 19672
rect 20579 19669 20591 19703
rect 20533 19663 20591 19669
rect 21358 19660 21364 19712
rect 21416 19700 21422 19712
rect 21726 19700 21732 19712
rect 21416 19672 21732 19700
rect 21416 19660 21422 19672
rect 21726 19660 21732 19672
rect 21784 19700 21790 19712
rect 22572 19700 22600 19740
rect 25314 19728 25320 19740
rect 25372 19768 25378 19780
rect 26252 19768 26280 19867
rect 25372 19740 26280 19768
rect 25372 19728 25378 19740
rect 21784 19672 22600 19700
rect 21784 19660 21790 19672
rect 22646 19660 22652 19712
rect 22704 19660 22710 19712
rect 22738 19660 22744 19712
rect 22796 19700 22802 19712
rect 23017 19703 23075 19709
rect 23017 19700 23029 19703
rect 22796 19672 23029 19700
rect 22796 19660 22802 19672
rect 23017 19669 23029 19672
rect 23063 19700 23075 19703
rect 23569 19703 23627 19709
rect 23569 19700 23581 19703
rect 23063 19672 23581 19700
rect 23063 19669 23075 19672
rect 23017 19663 23075 19669
rect 23569 19669 23581 19672
rect 23615 19700 23627 19703
rect 23750 19700 23756 19712
rect 23615 19672 23756 19700
rect 23615 19669 23627 19672
rect 23569 19663 23627 19669
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 24210 19660 24216 19712
rect 24268 19700 24274 19712
rect 26344 19700 26372 19876
rect 27338 19864 27344 19876
rect 27396 19864 27402 19916
rect 27522 19864 27528 19916
rect 27580 19904 27586 19916
rect 28537 19907 28595 19913
rect 28537 19904 28549 19907
rect 27580 19876 28549 19904
rect 27580 19864 27586 19876
rect 28537 19873 28549 19876
rect 28583 19873 28595 19907
rect 28537 19867 28595 19873
rect 27154 19796 27160 19848
rect 27212 19836 27218 19848
rect 27249 19839 27307 19845
rect 27249 19836 27261 19839
rect 27212 19808 27261 19836
rect 27212 19796 27218 19808
rect 27249 19805 27261 19808
rect 27295 19805 27307 19839
rect 27249 19799 27307 19805
rect 28353 19839 28411 19845
rect 28353 19805 28365 19839
rect 28399 19836 28411 19839
rect 29012 19836 29040 20012
rect 30926 20000 30932 20012
rect 30984 20040 30990 20052
rect 31570 20040 31576 20052
rect 30984 20012 31576 20040
rect 30984 20000 30990 20012
rect 31570 20000 31576 20012
rect 31628 20000 31634 20052
rect 31665 20043 31723 20049
rect 31665 20009 31677 20043
rect 31711 20040 31723 20043
rect 32766 20040 32772 20052
rect 31711 20012 32772 20040
rect 31711 20009 31723 20012
rect 31665 20003 31723 20009
rect 32766 20000 32772 20012
rect 32824 20000 32830 20052
rect 38194 20040 38200 20052
rect 34072 20012 38200 20040
rect 29365 19975 29423 19981
rect 29365 19941 29377 19975
rect 29411 19972 29423 19975
rect 29454 19972 29460 19984
rect 29411 19944 29460 19972
rect 29411 19941 29423 19944
rect 29365 19935 29423 19941
rect 29454 19932 29460 19944
rect 29512 19932 29518 19984
rect 34072 19972 34100 20012
rect 38194 20000 38200 20012
rect 38252 20000 38258 20052
rect 38286 20000 38292 20052
rect 38344 20040 38350 20052
rect 39577 20043 39635 20049
rect 39577 20040 39589 20043
rect 38344 20012 39589 20040
rect 38344 20000 38350 20012
rect 39577 20009 39589 20012
rect 39623 20009 39635 20043
rect 39577 20003 39635 20009
rect 41046 20000 41052 20052
rect 41104 20000 41110 20052
rect 46201 20043 46259 20049
rect 46201 20009 46213 20043
rect 46247 20040 46259 20043
rect 46382 20040 46388 20052
rect 46247 20012 46388 20040
rect 46247 20009 46259 20012
rect 46201 20003 46259 20009
rect 46382 20000 46388 20012
rect 46440 20000 46446 20052
rect 47118 20000 47124 20052
rect 47176 20040 47182 20052
rect 47305 20043 47363 20049
rect 47305 20040 47317 20043
rect 47176 20012 47317 20040
rect 47176 20000 47182 20012
rect 47305 20009 47317 20012
rect 47351 20009 47363 20043
rect 47305 20003 47363 20009
rect 30300 19944 32720 19972
rect 29086 19864 29092 19916
rect 29144 19904 29150 19916
rect 30300 19913 30328 19944
rect 32692 19913 32720 19944
rect 32784 19944 34100 19972
rect 34149 19975 34207 19981
rect 32784 19916 32812 19944
rect 34149 19941 34161 19975
rect 34195 19972 34207 19975
rect 34698 19972 34704 19984
rect 34195 19944 34704 19972
rect 34195 19941 34207 19944
rect 34149 19935 34207 19941
rect 34698 19932 34704 19944
rect 34756 19932 34762 19984
rect 43346 19972 43352 19984
rect 34900 19944 43352 19972
rect 30285 19907 30343 19913
rect 30285 19904 30297 19907
rect 29144 19876 30297 19904
rect 29144 19864 29150 19876
rect 30285 19873 30297 19876
rect 30331 19873 30343 19907
rect 30285 19867 30343 19873
rect 31113 19907 31171 19913
rect 31113 19873 31125 19907
rect 31159 19904 31171 19907
rect 32677 19907 32735 19913
rect 31159 19876 32444 19904
rect 31159 19873 31171 19876
rect 31113 19867 31171 19873
rect 28399 19808 29040 19836
rect 28399 19805 28411 19808
rect 28353 19799 28411 19805
rect 30098 19796 30104 19848
rect 30156 19836 30162 19848
rect 30926 19836 30932 19848
rect 30156 19808 30932 19836
rect 30156 19796 30162 19808
rect 30926 19796 30932 19808
rect 30984 19796 30990 19848
rect 31018 19796 31024 19848
rect 31076 19836 31082 19848
rect 31205 19839 31263 19845
rect 31205 19836 31217 19839
rect 31076 19808 31217 19836
rect 31076 19796 31082 19808
rect 31205 19805 31217 19808
rect 31251 19805 31263 19839
rect 31205 19799 31263 19805
rect 28997 19771 29055 19777
rect 28997 19768 29009 19771
rect 27172 19740 29009 19768
rect 27172 19712 27200 19740
rect 28997 19737 29009 19740
rect 29043 19768 29055 19771
rect 30374 19768 30380 19780
rect 29043 19740 30380 19768
rect 29043 19737 29055 19740
rect 28997 19731 29055 19737
rect 30374 19728 30380 19740
rect 30432 19728 30438 19780
rect 30466 19728 30472 19780
rect 30524 19768 30530 19780
rect 32306 19768 32312 19780
rect 30524 19740 32312 19768
rect 30524 19728 30530 19740
rect 32306 19728 32312 19740
rect 32364 19728 32370 19780
rect 24268 19672 26372 19700
rect 24268 19660 24274 19672
rect 26786 19660 26792 19712
rect 26844 19660 26850 19712
rect 27154 19660 27160 19712
rect 27212 19660 27218 19712
rect 27614 19660 27620 19712
rect 27672 19700 27678 19712
rect 27985 19703 28043 19709
rect 27985 19700 27997 19703
rect 27672 19672 27997 19700
rect 27672 19660 27678 19672
rect 27985 19669 27997 19672
rect 28031 19669 28043 19703
rect 27985 19663 28043 19669
rect 28445 19703 28503 19709
rect 28445 19669 28457 19703
rect 28491 19700 28503 19703
rect 29638 19700 29644 19712
rect 28491 19672 29644 19700
rect 28491 19669 28503 19672
rect 28445 19663 28503 19669
rect 29638 19660 29644 19672
rect 29696 19660 29702 19712
rect 29730 19660 29736 19712
rect 29788 19660 29794 19712
rect 30006 19660 30012 19712
rect 30064 19700 30070 19712
rect 30193 19703 30251 19709
rect 30193 19700 30205 19703
rect 30064 19672 30205 19700
rect 30064 19660 30070 19672
rect 30193 19669 30205 19672
rect 30239 19700 30251 19703
rect 30282 19700 30288 19712
rect 30239 19672 30288 19700
rect 30239 19669 30251 19672
rect 30193 19663 30251 19669
rect 30282 19660 30288 19672
rect 30340 19660 30346 19712
rect 31294 19660 31300 19712
rect 31352 19660 31358 19712
rect 32122 19660 32128 19712
rect 32180 19660 32186 19712
rect 32416 19700 32444 19876
rect 32677 19873 32689 19907
rect 32723 19873 32735 19907
rect 32677 19867 32735 19873
rect 32766 19864 32772 19916
rect 32824 19864 32830 19916
rect 33594 19864 33600 19916
rect 33652 19864 33658 19916
rect 33689 19907 33747 19913
rect 33689 19873 33701 19907
rect 33735 19904 33747 19907
rect 34900 19904 34928 19944
rect 43346 19932 43352 19944
rect 43404 19932 43410 19984
rect 44174 19932 44180 19984
rect 44232 19972 44238 19984
rect 46661 19975 46719 19981
rect 46661 19972 46673 19975
rect 44232 19944 46673 19972
rect 44232 19932 44238 19944
rect 46661 19941 46673 19944
rect 46707 19941 46719 19975
rect 46661 19935 46719 19941
rect 33735 19876 34928 19904
rect 33735 19873 33747 19876
rect 33689 19867 33747 19873
rect 32493 19839 32551 19845
rect 32493 19805 32505 19839
rect 32539 19836 32551 19839
rect 33778 19836 33784 19848
rect 32539 19808 33784 19836
rect 32539 19805 32551 19808
rect 32493 19799 32551 19805
rect 33778 19796 33784 19808
rect 33836 19796 33842 19848
rect 32585 19771 32643 19777
rect 32585 19737 32597 19771
rect 32631 19768 32643 19771
rect 33888 19768 33916 19876
rect 35066 19864 35072 19916
rect 35124 19864 35130 19916
rect 35161 19907 35219 19913
rect 35161 19873 35173 19907
rect 35207 19904 35219 19907
rect 35342 19904 35348 19916
rect 35207 19876 35348 19904
rect 35207 19873 35219 19876
rect 35161 19867 35219 19873
rect 35342 19864 35348 19876
rect 35400 19864 35406 19916
rect 36170 19864 36176 19916
rect 36228 19904 36234 19916
rect 36633 19907 36691 19913
rect 36633 19904 36645 19907
rect 36228 19876 36645 19904
rect 36228 19864 36234 19876
rect 36633 19873 36645 19876
rect 36679 19873 36691 19907
rect 36633 19867 36691 19873
rect 37366 19864 37372 19916
rect 37424 19904 37430 19916
rect 37921 19907 37979 19913
rect 37921 19904 37933 19907
rect 37424 19876 37933 19904
rect 37424 19864 37430 19876
rect 37921 19873 37933 19876
rect 37967 19873 37979 19907
rect 39025 19907 39083 19913
rect 39025 19904 39037 19907
rect 37921 19867 37979 19873
rect 38120 19876 39037 19904
rect 35253 19839 35311 19845
rect 35253 19805 35265 19839
rect 35299 19836 35311 19839
rect 35710 19836 35716 19848
rect 35299 19808 35716 19836
rect 35299 19805 35311 19808
rect 35253 19799 35311 19805
rect 35710 19796 35716 19808
rect 35768 19796 35774 19848
rect 37826 19796 37832 19848
rect 37884 19836 37890 19848
rect 38120 19845 38148 19876
rect 39025 19873 39037 19876
rect 39071 19873 39083 19907
rect 39025 19867 39083 19873
rect 39390 19864 39396 19916
rect 39448 19904 39454 19916
rect 40129 19907 40187 19913
rect 40129 19904 40141 19907
rect 39448 19876 40141 19904
rect 39448 19864 39454 19876
rect 40129 19873 40141 19876
rect 40175 19873 40187 19907
rect 40129 19867 40187 19873
rect 40310 19864 40316 19916
rect 40368 19904 40374 19916
rect 41233 19907 41291 19913
rect 41233 19904 41245 19907
rect 40368 19876 41245 19904
rect 40368 19864 40374 19876
rect 41233 19873 41245 19876
rect 41279 19873 41291 19907
rect 41233 19867 41291 19873
rect 45741 19907 45799 19913
rect 45741 19873 45753 19907
rect 45787 19904 45799 19907
rect 49234 19904 49240 19916
rect 45787 19876 49240 19904
rect 45787 19873 45799 19876
rect 45741 19867 45799 19873
rect 49234 19864 49240 19876
rect 49292 19864 49298 19916
rect 38105 19839 38163 19845
rect 38105 19836 38117 19839
rect 37884 19808 38117 19836
rect 37884 19796 37890 19808
rect 38105 19805 38117 19808
rect 38151 19805 38163 19839
rect 38105 19799 38163 19805
rect 38194 19796 38200 19848
rect 38252 19836 38258 19848
rect 38841 19839 38899 19845
rect 38841 19836 38853 19839
rect 38252 19808 38853 19836
rect 38252 19796 38258 19808
rect 38841 19805 38853 19808
rect 38887 19836 38899 19839
rect 39850 19836 39856 19848
rect 38887 19808 39856 19836
rect 38887 19805 38899 19808
rect 38841 19799 38899 19805
rect 39850 19796 39856 19808
rect 39908 19796 39914 19848
rect 40405 19839 40463 19845
rect 40405 19805 40417 19839
rect 40451 19836 40463 19839
rect 41046 19836 41052 19848
rect 40451 19808 41052 19836
rect 40451 19805 40463 19808
rect 40405 19799 40463 19805
rect 41046 19796 41052 19808
rect 41104 19796 41110 19848
rect 46014 19796 46020 19848
rect 46072 19796 46078 19848
rect 46842 19796 46848 19848
rect 46900 19796 46906 19848
rect 47489 19839 47547 19845
rect 47489 19805 47501 19839
rect 47535 19805 47547 19839
rect 47489 19799 47547 19805
rect 32631 19740 33916 19768
rect 32631 19737 32643 19740
rect 32585 19731 32643 19737
rect 34238 19728 34244 19780
rect 34296 19768 34302 19780
rect 36354 19768 36360 19780
rect 34296 19740 36360 19768
rect 34296 19728 34302 19740
rect 36354 19728 36360 19740
rect 36412 19728 36418 19780
rect 36449 19771 36507 19777
rect 36449 19737 36461 19771
rect 36495 19768 36507 19771
rect 40034 19768 40040 19780
rect 36495 19740 40040 19768
rect 36495 19737 36507 19740
rect 36449 19731 36507 19737
rect 40034 19728 40040 19740
rect 40092 19728 40098 19780
rect 33318 19700 33324 19712
rect 32416 19672 33324 19700
rect 33318 19660 33324 19672
rect 33376 19660 33382 19712
rect 33594 19660 33600 19712
rect 33652 19700 33658 19712
rect 34330 19700 34336 19712
rect 33652 19672 34336 19700
rect 33652 19660 33658 19672
rect 34330 19660 34336 19672
rect 34388 19700 34394 19712
rect 34425 19703 34483 19709
rect 34425 19700 34437 19703
rect 34388 19672 34437 19700
rect 34388 19660 34394 19672
rect 34425 19669 34437 19672
rect 34471 19669 34483 19703
rect 34425 19663 34483 19669
rect 35621 19703 35679 19709
rect 35621 19669 35633 19703
rect 35667 19700 35679 19703
rect 35802 19700 35808 19712
rect 35667 19672 35808 19700
rect 35667 19669 35679 19672
rect 35621 19663 35679 19669
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 36078 19660 36084 19712
rect 36136 19660 36142 19712
rect 36538 19660 36544 19712
rect 36596 19660 36602 19712
rect 37185 19703 37243 19709
rect 37185 19669 37197 19703
rect 37231 19700 37243 19703
rect 37369 19703 37427 19709
rect 37369 19700 37381 19703
rect 37231 19672 37381 19700
rect 37231 19669 37243 19672
rect 37185 19663 37243 19669
rect 37369 19669 37381 19672
rect 37415 19700 37427 19703
rect 37550 19700 37556 19712
rect 37415 19672 37556 19700
rect 37415 19669 37427 19672
rect 37369 19663 37427 19669
rect 37550 19660 37556 19672
rect 37608 19660 37614 19712
rect 38378 19660 38384 19712
rect 38436 19700 38442 19712
rect 38565 19703 38623 19709
rect 38565 19700 38577 19703
rect 38436 19672 38577 19700
rect 38436 19660 38442 19672
rect 38565 19669 38577 19672
rect 38611 19669 38623 19703
rect 38565 19663 38623 19669
rect 40773 19703 40831 19709
rect 40773 19669 40785 19703
rect 40819 19700 40831 19703
rect 40862 19700 40868 19712
rect 40819 19672 40868 19700
rect 40819 19669 40831 19672
rect 40773 19663 40831 19669
rect 40862 19660 40868 19672
rect 40920 19660 40926 19712
rect 46658 19660 46664 19712
rect 46716 19700 46722 19712
rect 47504 19700 47532 19799
rect 47578 19796 47584 19848
rect 47636 19836 47642 19848
rect 49329 19839 49387 19845
rect 49329 19836 49341 19839
rect 47636 19808 49341 19836
rect 47636 19796 47642 19808
rect 49329 19805 49341 19808
rect 49375 19836 49387 19839
rect 49418 19836 49424 19848
rect 49375 19808 49424 19836
rect 49375 19805 49387 19808
rect 49329 19799 49387 19805
rect 49418 19796 49424 19808
rect 49476 19796 49482 19848
rect 47670 19728 47676 19780
rect 47728 19768 47734 19780
rect 47949 19771 48007 19777
rect 47949 19768 47961 19771
rect 47728 19740 47961 19768
rect 47728 19728 47734 19740
rect 47949 19737 47961 19740
rect 47995 19737 48007 19771
rect 47949 19731 48007 19737
rect 48133 19771 48191 19777
rect 48133 19737 48145 19771
rect 48179 19768 48191 19771
rect 48685 19771 48743 19777
rect 48685 19768 48697 19771
rect 48179 19740 48697 19768
rect 48179 19737 48191 19740
rect 48133 19731 48191 19737
rect 48685 19737 48697 19740
rect 48731 19737 48743 19771
rect 48685 19731 48743 19737
rect 46716 19672 47532 19700
rect 46716 19660 46722 19672
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 7616 19468 10977 19496
rect 7616 19456 7622 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 13446 19496 13452 19508
rect 12492 19468 13452 19496
rect 12492 19456 12498 19468
rect 13446 19456 13452 19468
rect 13504 19496 13510 19508
rect 13504 19468 14504 19496
rect 13504 19456 13510 19468
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 3476 19400 3617 19428
rect 3476 19388 3482 19400
rect 3605 19397 3617 19400
rect 3651 19397 3663 19431
rect 9214 19428 9220 19440
rect 3605 19391 3663 19397
rect 4540 19400 9220 19428
rect 1762 19320 1768 19372
rect 1820 19320 1826 19372
rect 2961 19363 3019 19369
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 4540 19360 4568 19400
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 10505 19431 10563 19437
rect 10505 19397 10517 19431
rect 10551 19428 10563 19431
rect 12250 19428 12256 19440
rect 10551 19400 12256 19428
rect 10551 19397 10563 19400
rect 10505 19391 10563 19397
rect 12250 19388 12256 19400
rect 12308 19388 12314 19440
rect 13170 19388 13176 19440
rect 13228 19388 13234 19440
rect 14476 19428 14504 19468
rect 15378 19456 15384 19508
rect 15436 19456 15442 19508
rect 15470 19456 15476 19508
rect 15528 19496 15534 19508
rect 16114 19496 16120 19508
rect 15528 19468 16120 19496
rect 15528 19456 15534 19468
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 16850 19456 16856 19508
rect 16908 19456 16914 19508
rect 17310 19456 17316 19508
rect 17368 19496 17374 19508
rect 19886 19496 19892 19508
rect 17368 19468 19892 19496
rect 17368 19456 17374 19468
rect 19886 19456 19892 19468
rect 19944 19456 19950 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 25406 19496 25412 19508
rect 21223 19468 25412 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 16022 19428 16028 19440
rect 14476 19400 16028 19428
rect 3007 19332 4568 19360
rect 4801 19363 4859 19369
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 5445 19363 5503 19369
rect 4847 19332 5396 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 5261 19295 5319 19301
rect 5261 19292 5273 19295
rect 3936 19264 5273 19292
rect 3936 19252 3942 19264
rect 5261 19261 5273 19264
rect 5307 19261 5319 19295
rect 5368 19292 5396 19332
rect 5445 19329 5457 19363
rect 5491 19360 5503 19363
rect 5810 19360 5816 19372
rect 5491 19332 5816 19360
rect 5491 19329 5503 19332
rect 5445 19323 5503 19329
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 11606 19360 11612 19372
rect 11195 19332 11612 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 11747 19332 12173 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 12161 19329 12173 19332
rect 12207 19360 12219 19363
rect 12894 19360 12900 19372
rect 12207 19332 12434 19360
rect 12207 19329 12219 19332
rect 12161 19323 12219 19329
rect 6822 19292 6828 19304
rect 5368 19264 6828 19292
rect 5261 19255 5319 19261
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19292 9919 19295
rect 10410 19292 10416 19304
rect 9907 19264 10416 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 12406 19292 12434 19332
rect 12544 19332 12900 19360
rect 12544 19292 12572 19332
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 14476 19369 14504 19400
rect 16022 19388 16028 19400
rect 16080 19428 16086 19440
rect 16942 19428 16948 19440
rect 16080 19400 16948 19428
rect 16080 19388 16086 19400
rect 16942 19388 16948 19400
rect 17000 19388 17006 19440
rect 18049 19431 18107 19437
rect 18049 19397 18061 19431
rect 18095 19428 18107 19431
rect 18322 19428 18328 19440
rect 18095 19400 18328 19428
rect 18095 19397 18107 19400
rect 18049 19391 18107 19397
rect 18322 19388 18328 19400
rect 18380 19388 18386 19440
rect 19518 19388 19524 19440
rect 19576 19428 19582 19440
rect 20732 19428 20760 19459
rect 25406 19456 25412 19468
rect 25464 19456 25470 19508
rect 25498 19456 25504 19508
rect 25556 19496 25562 19508
rect 28258 19496 28264 19508
rect 25556 19468 28264 19496
rect 25556 19456 25562 19468
rect 28258 19456 28264 19468
rect 28316 19456 28322 19508
rect 28445 19499 28503 19505
rect 28445 19465 28457 19499
rect 28491 19496 28503 19499
rect 28718 19496 28724 19508
rect 28491 19468 28724 19496
rect 28491 19465 28503 19468
rect 28445 19459 28503 19465
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 31386 19456 31392 19508
rect 31444 19496 31450 19508
rect 32677 19499 32735 19505
rect 32677 19496 32689 19499
rect 31444 19468 32689 19496
rect 31444 19456 31450 19468
rect 32677 19465 32689 19468
rect 32723 19465 32735 19499
rect 32677 19459 32735 19465
rect 32858 19456 32864 19508
rect 32916 19496 32922 19508
rect 33045 19499 33103 19505
rect 33045 19496 33057 19499
rect 32916 19468 33057 19496
rect 32916 19456 32922 19468
rect 33045 19465 33057 19468
rect 33091 19465 33103 19499
rect 33045 19459 33103 19465
rect 34238 19456 34244 19508
rect 34296 19456 34302 19508
rect 34882 19456 34888 19508
rect 34940 19496 34946 19508
rect 35069 19499 35127 19505
rect 35069 19496 35081 19499
rect 34940 19468 35081 19496
rect 34940 19456 34946 19468
rect 35069 19465 35081 19468
rect 35115 19465 35127 19499
rect 35069 19459 35127 19465
rect 35437 19499 35495 19505
rect 35437 19465 35449 19499
rect 35483 19496 35495 19499
rect 36538 19496 36544 19508
rect 35483 19468 36544 19496
rect 35483 19465 35495 19468
rect 35437 19459 35495 19465
rect 36538 19456 36544 19468
rect 36596 19456 36602 19508
rect 36906 19456 36912 19508
rect 36964 19496 36970 19508
rect 37277 19499 37335 19505
rect 37277 19496 37289 19499
rect 36964 19468 37289 19496
rect 36964 19456 36970 19468
rect 37277 19465 37289 19468
rect 37323 19496 37335 19499
rect 38470 19496 38476 19508
rect 37323 19468 38476 19496
rect 37323 19465 37335 19468
rect 37277 19459 37335 19465
rect 38470 19456 38476 19468
rect 38528 19456 38534 19508
rect 40034 19456 40040 19508
rect 40092 19496 40098 19508
rect 40129 19499 40187 19505
rect 40129 19496 40141 19499
rect 40092 19468 40141 19496
rect 40092 19456 40098 19468
rect 40129 19465 40141 19468
rect 40175 19465 40187 19499
rect 40129 19459 40187 19465
rect 40497 19499 40555 19505
rect 40497 19465 40509 19499
rect 40543 19496 40555 19499
rect 47029 19499 47087 19505
rect 47029 19496 47041 19499
rect 40543 19468 47041 19496
rect 40543 19465 40555 19468
rect 40497 19459 40555 19465
rect 47029 19465 47041 19468
rect 47075 19465 47087 19499
rect 47029 19459 47087 19465
rect 47673 19499 47731 19505
rect 47673 19465 47685 19499
rect 47719 19496 47731 19499
rect 48406 19496 48412 19508
rect 47719 19468 48412 19496
rect 47719 19465 47731 19468
rect 47673 19459 47731 19465
rect 19576 19400 20760 19428
rect 19576 19388 19582 19400
rect 22094 19388 22100 19440
rect 22152 19388 22158 19440
rect 22646 19388 22652 19440
rect 22704 19428 22710 19440
rect 22925 19431 22983 19437
rect 22925 19428 22937 19431
rect 22704 19400 22937 19428
rect 22704 19388 22710 19400
rect 22925 19397 22937 19400
rect 22971 19397 22983 19431
rect 22925 19391 22983 19397
rect 24486 19388 24492 19440
rect 24544 19388 24550 19440
rect 26142 19388 26148 19440
rect 26200 19428 26206 19440
rect 28626 19428 28632 19440
rect 26200 19400 28632 19428
rect 26200 19388 26206 19400
rect 28626 19388 28632 19400
rect 28684 19388 28690 19440
rect 28966 19400 29132 19428
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 15930 19360 15936 19372
rect 15519 19332 15936 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 16209 19363 16267 19369
rect 16209 19329 16221 19363
rect 16255 19360 16267 19363
rect 16666 19360 16672 19372
rect 16255 19332 16672 19360
rect 16255 19329 16267 19332
rect 16209 19323 16267 19329
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 17184 19332 17233 19360
rect 17184 19320 17190 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 18414 19360 18420 19372
rect 17359 19332 18420 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 21085 19363 21143 19369
rect 18524 19332 18828 19360
rect 11900 19264 12296 19292
rect 12406 19264 12572 19292
rect 7466 19184 7472 19236
rect 7524 19224 7530 19236
rect 11900 19224 11928 19264
rect 7524 19196 11928 19224
rect 7524 19184 7530 19196
rect 11974 19184 11980 19236
rect 12032 19184 12038 19236
rect 12268 19224 12296 19264
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 13722 19292 13728 19304
rect 12676 19264 13728 19292
rect 12676 19252 12682 19264
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 14231 19264 14504 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 14476 19224 14504 19264
rect 14550 19252 14556 19304
rect 14608 19292 14614 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14608 19264 14841 19292
rect 14608 19252 14614 19264
rect 14829 19261 14841 19264
rect 14875 19292 14887 19295
rect 17034 19292 17040 19304
rect 14875 19264 17040 19292
rect 14875 19261 14887 19264
rect 14829 19255 14887 19261
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 12268 19196 13216 19224
rect 14476 19196 15148 19224
rect 5810 19116 5816 19168
rect 5868 19116 5874 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 11882 19156 11888 19168
rect 8352 19128 11888 19156
rect 8352 19116 8358 19128
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12713 19159 12771 19165
rect 12713 19125 12725 19159
rect 12759 19156 12771 19159
rect 12802 19156 12808 19168
rect 12759 19128 12808 19156
rect 12759 19125 12771 19128
rect 12713 19119 12771 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13188 19156 13216 19196
rect 13814 19156 13820 19168
rect 13188 19128 13820 19156
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 15010 19116 15016 19168
rect 15068 19116 15074 19168
rect 15120 19156 15148 19196
rect 15194 19184 15200 19236
rect 15252 19224 15258 19236
rect 16025 19227 16083 19233
rect 16025 19224 16037 19227
rect 15252 19196 16037 19224
rect 15252 19184 15258 19196
rect 16025 19193 16037 19196
rect 16071 19193 16083 19227
rect 16025 19187 16083 19193
rect 16114 19184 16120 19236
rect 16172 19224 16178 19236
rect 17420 19224 17448 19255
rect 16172 19196 17448 19224
rect 16172 19184 16178 19196
rect 15930 19156 15936 19168
rect 15120 19128 15936 19156
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 18524 19156 18552 19332
rect 18800 19292 18828 19332
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 23290 19360 23296 19372
rect 21131 19332 23296 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19360 25283 19363
rect 25682 19360 25688 19372
rect 25271 19332 25688 19360
rect 25271 19329 25283 19332
rect 25225 19323 25283 19329
rect 25682 19320 25688 19332
rect 25740 19320 25746 19372
rect 26237 19363 26295 19369
rect 26237 19329 26249 19363
rect 26283 19360 26295 19363
rect 26418 19360 26424 19372
rect 26283 19332 26424 19360
rect 26283 19329 26295 19332
rect 26237 19323 26295 19329
rect 26418 19320 26424 19332
rect 26476 19320 26482 19372
rect 27617 19363 27675 19369
rect 27617 19329 27629 19363
rect 27663 19360 27675 19363
rect 28350 19360 28356 19372
rect 27663 19332 28356 19360
rect 27663 19329 27675 19332
rect 27617 19323 27675 19329
rect 28350 19320 28356 19332
rect 28408 19320 28414 19372
rect 28813 19363 28871 19369
rect 28813 19329 28825 19363
rect 28859 19360 28871 19363
rect 28966 19360 28994 19400
rect 28859 19332 28994 19360
rect 29104 19360 29132 19400
rect 31478 19388 31484 19440
rect 31536 19388 31542 19440
rect 31754 19388 31760 19440
rect 31812 19428 31818 19440
rect 32585 19431 32643 19437
rect 32585 19428 32597 19431
rect 31812 19400 32597 19428
rect 31812 19388 31818 19400
rect 32585 19397 32597 19400
rect 32631 19397 32643 19431
rect 32585 19391 32643 19397
rect 33778 19388 33784 19440
rect 33836 19428 33842 19440
rect 34606 19428 34612 19440
rect 33836 19400 34612 19428
rect 33836 19388 33842 19400
rect 34606 19388 34612 19400
rect 34664 19388 34670 19440
rect 34974 19388 34980 19440
rect 35032 19428 35038 19440
rect 36173 19431 36231 19437
rect 36173 19428 36185 19431
rect 35032 19400 36185 19428
rect 35032 19388 35038 19400
rect 36173 19397 36185 19400
rect 36219 19397 36231 19431
rect 36173 19391 36231 19397
rect 46385 19431 46443 19437
rect 46385 19397 46397 19431
rect 46431 19428 46443 19431
rect 47578 19428 47584 19440
rect 46431 19400 47584 19428
rect 46431 19397 46443 19400
rect 46385 19391 46443 19397
rect 47578 19388 47584 19400
rect 47636 19388 47642 19440
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 29104 19332 29745 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 30282 19320 30288 19372
rect 30340 19320 30346 19372
rect 30745 19363 30803 19369
rect 30745 19329 30757 19363
rect 30791 19329 30803 19363
rect 30745 19323 30803 19329
rect 19426 19292 19432 19304
rect 18800 19264 19432 19292
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 19794 19252 19800 19304
rect 19852 19252 19858 19304
rect 20073 19295 20131 19301
rect 20073 19261 20085 19295
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 21407 19264 22094 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 17000 19128 18552 19156
rect 17000 19116 17006 19128
rect 19610 19116 19616 19168
rect 19668 19156 19674 19168
rect 20088 19156 20116 19255
rect 19668 19128 20116 19156
rect 20441 19159 20499 19165
rect 19668 19116 19674 19128
rect 20441 19125 20453 19159
rect 20487 19156 20499 19159
rect 20530 19156 20536 19168
rect 20487 19128 20536 19156
rect 20487 19125 20499 19128
rect 20441 19119 20499 19125
rect 20530 19116 20536 19128
rect 20588 19156 20594 19168
rect 20898 19156 20904 19168
rect 20588 19128 20904 19156
rect 20588 19116 20594 19128
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 22066 19156 22094 19264
rect 24946 19252 24952 19304
rect 25004 19292 25010 19304
rect 25590 19292 25596 19304
rect 25004 19264 25596 19292
rect 25004 19252 25010 19264
rect 25590 19252 25596 19264
rect 25648 19252 25654 19304
rect 26326 19252 26332 19304
rect 26384 19292 26390 19304
rect 27522 19292 27528 19304
rect 26384 19264 27528 19292
rect 26384 19252 26390 19264
rect 27522 19252 27528 19264
rect 27580 19252 27586 19304
rect 27706 19252 27712 19304
rect 27764 19252 27770 19304
rect 27801 19295 27859 19301
rect 27801 19261 27813 19295
rect 27847 19292 27859 19295
rect 28166 19292 28172 19304
rect 27847 19264 28172 19292
rect 27847 19261 27859 19264
rect 27801 19255 27859 19261
rect 22278 19184 22284 19236
rect 22336 19224 22342 19236
rect 22336 19196 23980 19224
rect 22336 19184 22342 19196
rect 23477 19159 23535 19165
rect 23477 19156 23489 19159
rect 22066 19128 23489 19156
rect 23477 19125 23489 19128
rect 23523 19156 23535 19159
rect 23842 19156 23848 19168
rect 23523 19128 23848 19156
rect 23523 19125 23535 19128
rect 23477 19119 23535 19125
rect 23842 19116 23848 19128
rect 23900 19116 23906 19168
rect 23952 19156 23980 19196
rect 25222 19184 25228 19236
rect 25280 19224 25286 19236
rect 26602 19224 26608 19236
rect 25280 19196 26608 19224
rect 25280 19184 25286 19196
rect 26602 19184 26608 19196
rect 26660 19184 26666 19236
rect 26786 19184 26792 19236
rect 26844 19224 26850 19236
rect 27816 19224 27844 19255
rect 28166 19252 28172 19264
rect 28224 19252 28230 19304
rect 28626 19252 28632 19304
rect 28684 19292 28690 19304
rect 28905 19295 28963 19301
rect 28905 19292 28917 19295
rect 28684 19264 28917 19292
rect 28684 19252 28690 19264
rect 28905 19261 28917 19264
rect 28951 19261 28963 19295
rect 28905 19255 28963 19261
rect 29089 19295 29147 19301
rect 29089 19261 29101 19295
rect 29135 19292 29147 19295
rect 29362 19292 29368 19304
rect 29135 19264 29368 19292
rect 29135 19261 29147 19264
rect 29089 19255 29147 19261
rect 26844 19196 27844 19224
rect 26844 19184 26850 19196
rect 28258 19184 28264 19236
rect 28316 19224 28322 19236
rect 29104 19224 29132 19255
rect 29362 19252 29368 19264
rect 29420 19252 29426 19304
rect 30300 19292 30328 19320
rect 29472 19264 30328 19292
rect 29472 19236 29500 19264
rect 30374 19252 30380 19304
rect 30432 19292 30438 19304
rect 30760 19292 30788 19323
rect 33870 19320 33876 19372
rect 33928 19320 33934 19372
rect 34790 19320 34796 19372
rect 34848 19360 34854 19372
rect 34848 19332 35020 19360
rect 34848 19320 34854 19332
rect 30432 19264 30788 19292
rect 30432 19252 30438 19264
rect 32306 19252 32312 19304
rect 32364 19292 32370 19304
rect 32401 19295 32459 19301
rect 32401 19292 32413 19295
rect 32364 19264 32413 19292
rect 32364 19252 32370 19264
rect 32401 19261 32413 19264
rect 32447 19261 32459 19295
rect 32401 19255 32459 19261
rect 32674 19252 32680 19304
rect 32732 19292 32738 19304
rect 33594 19292 33600 19304
rect 32732 19264 33600 19292
rect 32732 19252 32738 19264
rect 33594 19252 33600 19264
rect 33652 19252 33658 19304
rect 33689 19295 33747 19301
rect 33689 19261 33701 19295
rect 33735 19292 33747 19295
rect 34422 19292 34428 19304
rect 33735 19264 34428 19292
rect 33735 19261 33747 19264
rect 33689 19255 33747 19261
rect 34422 19252 34428 19264
rect 34480 19252 34486 19304
rect 34992 19301 35020 19332
rect 35894 19320 35900 19372
rect 35952 19360 35958 19372
rect 36265 19363 36323 19369
rect 36265 19360 36277 19363
rect 35952 19332 36277 19360
rect 35952 19320 35958 19332
rect 36265 19329 36277 19332
rect 36311 19329 36323 19363
rect 36265 19323 36323 19329
rect 38286 19320 38292 19372
rect 38344 19320 38350 19372
rect 40586 19320 40592 19372
rect 40644 19360 40650 19372
rect 41325 19363 41383 19369
rect 41325 19360 41337 19363
rect 40644 19332 41337 19360
rect 40644 19320 40650 19332
rect 41325 19329 41337 19332
rect 41371 19360 41383 19363
rect 47026 19360 47032 19372
rect 41371 19332 47032 19360
rect 41371 19329 41383 19332
rect 41325 19323 41383 19329
rect 47026 19320 47032 19332
rect 47084 19320 47090 19372
rect 47213 19363 47271 19369
rect 47213 19329 47225 19363
rect 47259 19360 47271 19363
rect 47688 19360 47716 19459
rect 48406 19456 48412 19468
rect 48464 19456 48470 19508
rect 47259 19332 47716 19360
rect 48133 19363 48191 19369
rect 47259 19329 47271 19332
rect 47213 19323 47271 19329
rect 48133 19329 48145 19363
rect 48179 19360 48191 19363
rect 48685 19363 48743 19369
rect 48685 19360 48697 19363
rect 48179 19332 48697 19360
rect 48179 19329 48191 19332
rect 48133 19323 48191 19329
rect 48685 19329 48697 19332
rect 48731 19329 48743 19363
rect 48685 19323 48743 19329
rect 49326 19320 49332 19372
rect 49384 19320 49390 19372
rect 34885 19295 34943 19301
rect 34885 19261 34897 19295
rect 34931 19261 34943 19295
rect 34885 19255 34943 19261
rect 34977 19295 35035 19301
rect 34977 19261 34989 19295
rect 35023 19261 35035 19295
rect 34977 19255 35035 19261
rect 28316 19196 29132 19224
rect 28316 19184 28322 19196
rect 29454 19184 29460 19236
rect 29512 19184 29518 19236
rect 29638 19184 29644 19236
rect 29696 19184 29702 19236
rect 30193 19227 30251 19233
rect 30193 19193 30205 19227
rect 30239 19193 30251 19227
rect 30193 19187 30251 19193
rect 25240 19156 25268 19184
rect 23952 19128 25268 19156
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 27246 19116 27252 19168
rect 27304 19116 27310 19168
rect 27706 19116 27712 19168
rect 27764 19156 27770 19168
rect 28442 19156 28448 19168
rect 27764 19128 28448 19156
rect 27764 19116 27770 19128
rect 28442 19116 28448 19128
rect 28500 19156 28506 19168
rect 29086 19156 29092 19168
rect 28500 19128 29092 19156
rect 28500 19116 28506 19128
rect 29086 19116 29092 19128
rect 29144 19116 29150 19168
rect 29656 19156 29684 19184
rect 30208 19156 30236 19187
rect 30282 19184 30288 19236
rect 30340 19224 30346 19236
rect 34900 19224 34928 19255
rect 35986 19252 35992 19304
rect 36044 19252 36050 19304
rect 37553 19295 37611 19301
rect 37553 19261 37565 19295
rect 37599 19292 37611 19295
rect 37826 19292 37832 19304
rect 37599 19264 37832 19292
rect 37599 19261 37611 19264
rect 37553 19255 37611 19261
rect 37826 19252 37832 19264
rect 37884 19292 37890 19304
rect 38304 19292 38332 19320
rect 37884 19264 38332 19292
rect 37884 19252 37890 19264
rect 39390 19252 39396 19304
rect 39448 19252 39454 19304
rect 39666 19252 39672 19304
rect 39724 19252 39730 19304
rect 40681 19295 40739 19301
rect 40681 19292 40693 19295
rect 39776 19264 40693 19292
rect 37734 19224 37740 19236
rect 30340 19196 33732 19224
rect 34900 19196 37740 19224
rect 30340 19184 30346 19196
rect 33704 19168 33732 19196
rect 37734 19184 37740 19196
rect 37792 19224 37798 19236
rect 37792 19196 38056 19224
rect 37792 19184 37798 19196
rect 31754 19156 31760 19168
rect 29656 19128 31760 19156
rect 31754 19116 31760 19128
rect 31812 19116 31818 19168
rect 32490 19116 32496 19168
rect 32548 19156 32554 19168
rect 33410 19156 33416 19168
rect 32548 19128 33416 19156
rect 32548 19116 32554 19128
rect 33410 19116 33416 19128
rect 33468 19116 33474 19168
rect 33686 19116 33692 19168
rect 33744 19116 33750 19168
rect 33778 19116 33784 19168
rect 33836 19156 33842 19168
rect 36446 19156 36452 19168
rect 33836 19128 36452 19156
rect 33836 19116 33842 19128
rect 36446 19116 36452 19128
rect 36504 19116 36510 19168
rect 36630 19116 36636 19168
rect 36688 19116 36694 19168
rect 36906 19116 36912 19168
rect 36964 19116 36970 19168
rect 37826 19116 37832 19168
rect 37884 19156 37890 19168
rect 37921 19159 37979 19165
rect 37921 19156 37933 19159
rect 37884 19128 37933 19156
rect 37884 19116 37890 19128
rect 37921 19125 37933 19128
rect 37967 19125 37979 19159
rect 38028 19156 38056 19196
rect 39776 19156 39804 19264
rect 40681 19261 40693 19264
rect 40727 19261 40739 19295
rect 40681 19255 40739 19261
rect 46569 19295 46627 19301
rect 46569 19261 46581 19295
rect 46615 19292 46627 19295
rect 49344 19292 49372 19320
rect 46615 19264 49372 19292
rect 46615 19261 46627 19264
rect 46569 19255 46627 19261
rect 39850 19184 39856 19236
rect 39908 19224 39914 19236
rect 47949 19227 48007 19233
rect 47949 19224 47961 19227
rect 39908 19196 47961 19224
rect 39908 19184 39914 19196
rect 47949 19193 47961 19196
rect 47995 19193 48007 19227
rect 47949 19187 48007 19193
rect 38028 19128 39804 19156
rect 37921 19119 37979 19125
rect 40494 19116 40500 19168
rect 40552 19156 40558 19168
rect 41141 19159 41199 19165
rect 41141 19156 41153 19159
rect 40552 19128 41153 19156
rect 40552 19116 40558 19128
rect 41141 19125 41153 19128
rect 41187 19156 41199 19159
rect 42058 19156 42064 19168
rect 41187 19128 42064 19156
rect 41187 19125 41199 19128
rect 41141 19119 41199 19125
rect 42058 19116 42064 19128
rect 42116 19116 42122 19168
rect 46658 19116 46664 19168
rect 46716 19116 46722 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 6880 18924 9229 18952
rect 6880 18912 6886 18924
rect 9217 18921 9229 18924
rect 9263 18952 9275 18955
rect 11146 18952 11152 18964
rect 9263 18924 11152 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 11514 18912 11520 18964
rect 11572 18952 11578 18964
rect 12529 18955 12587 18961
rect 12529 18952 12541 18955
rect 11572 18924 12541 18952
rect 11572 18912 11578 18924
rect 12529 18921 12541 18924
rect 12575 18921 12587 18955
rect 12529 18915 12587 18921
rect 13630 18912 13636 18964
rect 13688 18912 13694 18964
rect 13814 18912 13820 18964
rect 13872 18912 13878 18964
rect 13924 18924 15884 18952
rect 11238 18884 11244 18896
rect 10888 18856 11244 18884
rect 3786 18776 3792 18828
rect 3844 18816 3850 18828
rect 4157 18819 4215 18825
rect 4157 18816 4169 18819
rect 3844 18788 4169 18816
rect 3844 18776 3850 18788
rect 4157 18785 4169 18788
rect 4203 18785 4215 18819
rect 10888 18816 10916 18856
rect 11238 18844 11244 18856
rect 11296 18844 11302 18896
rect 11882 18844 11888 18896
rect 11940 18844 11946 18896
rect 13354 18844 13360 18896
rect 13412 18884 13418 18896
rect 13924 18884 13952 18924
rect 13412 18856 13952 18884
rect 13412 18844 13418 18856
rect 4157 18779 4215 18785
rect 8312 18788 10916 18816
rect 10965 18819 11023 18825
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18717 3019 18751
rect 2961 18711 3019 18717
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 7742 18748 7748 18760
rect 5399 18720 7748 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 1394 18640 1400 18692
rect 1452 18680 1458 18692
rect 1765 18683 1823 18689
rect 1765 18680 1777 18683
rect 1452 18652 1777 18680
rect 1452 18640 1458 18652
rect 1765 18649 1777 18652
rect 1811 18649 1823 18683
rect 1765 18643 1823 18649
rect 2976 18612 3004 18711
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 8312 18757 8340 18788
rect 10965 18785 10977 18819
rect 11011 18816 11023 18819
rect 12434 18816 12440 18828
rect 11011 18788 12440 18816
rect 11011 18785 11023 18788
rect 10965 18779 11023 18785
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 13078 18776 13084 18828
rect 13136 18776 13142 18828
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18816 14335 18819
rect 14550 18816 14556 18828
rect 14323 18788 14556 18816
rect 14323 18785 14335 18788
rect 14277 18779 14335 18785
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 15010 18776 15016 18828
rect 15068 18816 15074 18828
rect 15068 18788 15608 18816
rect 15068 18776 15074 18788
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 8113 18683 8171 18689
rect 8113 18680 8125 18683
rect 4396 18652 8125 18680
rect 4396 18640 4402 18652
rect 8113 18649 8125 18652
rect 8159 18649 8171 18683
rect 8113 18643 8171 18649
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10284 18652 10640 18680
rect 10284 18640 10290 18652
rect 7374 18612 7380 18624
rect 2976 18584 7380 18612
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 10612 18612 10640 18652
rect 10686 18640 10692 18692
rect 10744 18640 10750 18692
rect 12084 18680 12112 18711
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 15580 18748 15608 18788
rect 15654 18748 15660 18760
rect 12308 18720 12664 18748
rect 15580 18720 15660 18748
rect 12308 18708 12314 18720
rect 12434 18680 12440 18692
rect 12084 18652 12440 18680
rect 12434 18640 12440 18652
rect 12492 18640 12498 18692
rect 12636 18680 12664 18720
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 15856 18748 15884 18924
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 16025 18955 16083 18961
rect 16025 18952 16037 18955
rect 15988 18924 16037 18952
rect 15988 18912 15994 18924
rect 16025 18921 16037 18924
rect 16071 18952 16083 18955
rect 16114 18952 16120 18964
rect 16071 18924 16120 18952
rect 16071 18921 16083 18924
rect 16025 18915 16083 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 18141 18955 18199 18961
rect 18141 18952 18153 18955
rect 16540 18924 18153 18952
rect 16540 18912 16546 18924
rect 18141 18921 18153 18924
rect 18187 18921 18199 18955
rect 18141 18915 18199 18921
rect 19886 18912 19892 18964
rect 19944 18912 19950 18964
rect 20364 18924 22094 18952
rect 16758 18844 16764 18896
rect 16816 18884 16822 18896
rect 16945 18887 17003 18893
rect 16945 18884 16957 18887
rect 16816 18856 16957 18884
rect 16816 18844 16822 18856
rect 16945 18853 16957 18856
rect 16991 18853 17003 18887
rect 16945 18847 17003 18853
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 16632 18788 17509 18816
rect 16632 18776 16638 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 19702 18816 19708 18828
rect 18831 18788 19708 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 20364 18825 20392 18924
rect 20714 18844 20720 18896
rect 20772 18884 20778 18896
rect 21085 18887 21143 18893
rect 21085 18884 21097 18887
rect 20772 18856 21097 18884
rect 20772 18844 20778 18856
rect 21085 18853 21097 18856
rect 21131 18853 21143 18887
rect 21085 18847 21143 18853
rect 20349 18819 20407 18825
rect 20349 18785 20361 18819
rect 20395 18785 20407 18819
rect 20349 18779 20407 18785
rect 20438 18776 20444 18828
rect 20496 18776 20502 18828
rect 21174 18776 21180 18828
rect 21232 18816 21238 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21232 18788 21649 18816
rect 21232 18776 21238 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 22066 18816 22094 18924
rect 22278 18912 22284 18964
rect 22336 18912 22342 18964
rect 22738 18912 22744 18964
rect 22796 18952 22802 18964
rect 27614 18952 27620 18964
rect 22796 18924 27620 18952
rect 22796 18912 22802 18924
rect 27614 18912 27620 18924
rect 27672 18912 27678 18964
rect 27706 18912 27712 18964
rect 27764 18952 27770 18964
rect 28077 18955 28135 18961
rect 28077 18952 28089 18955
rect 27764 18924 28089 18952
rect 27764 18912 27770 18924
rect 28077 18921 28089 18924
rect 28123 18952 28135 18955
rect 30006 18952 30012 18964
rect 28123 18924 30012 18952
rect 28123 18921 28135 18924
rect 28077 18915 28135 18921
rect 30006 18912 30012 18924
rect 30064 18912 30070 18964
rect 30926 18912 30932 18964
rect 30984 18912 30990 18964
rect 32950 18912 32956 18964
rect 33008 18952 33014 18964
rect 33781 18955 33839 18961
rect 33781 18952 33793 18955
rect 33008 18924 33793 18952
rect 33008 18912 33014 18924
rect 33781 18921 33793 18924
rect 33827 18952 33839 18955
rect 34974 18952 34980 18964
rect 33827 18924 34980 18952
rect 33827 18921 33839 18924
rect 33781 18915 33839 18921
rect 34974 18912 34980 18924
rect 35032 18912 35038 18964
rect 37369 18955 37427 18961
rect 35084 18924 36952 18952
rect 25056 18856 25912 18884
rect 25056 18816 25084 18856
rect 22066 18788 25084 18816
rect 21637 18779 21695 18785
rect 25222 18776 25228 18828
rect 25280 18776 25286 18828
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 25740 18788 25789 18816
rect 25740 18776 25746 18788
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 25884 18816 25912 18856
rect 27062 18844 27068 18896
rect 27120 18884 27126 18896
rect 31481 18887 31539 18893
rect 31481 18884 31493 18887
rect 27120 18856 31493 18884
rect 27120 18844 27126 18856
rect 31481 18853 31493 18856
rect 31527 18853 31539 18887
rect 32674 18884 32680 18896
rect 31481 18847 31539 18853
rect 31956 18856 32680 18884
rect 26694 18816 26700 18828
rect 25884 18788 26700 18816
rect 25777 18779 25835 18785
rect 26694 18776 26700 18788
rect 26752 18776 26758 18828
rect 27525 18819 27583 18825
rect 27525 18785 27537 18819
rect 27571 18816 27583 18819
rect 28442 18816 28448 18828
rect 27571 18788 28448 18816
rect 27571 18785 27583 18788
rect 27525 18779 27583 18785
rect 28442 18776 28448 18788
rect 28500 18816 28506 18828
rect 28902 18816 28908 18828
rect 28500 18788 28908 18816
rect 28500 18776 28506 18788
rect 28902 18776 28908 18788
rect 28960 18776 28966 18828
rect 29638 18816 29644 18828
rect 29104 18788 29644 18816
rect 15856 18720 17540 18748
rect 12897 18683 12955 18689
rect 12897 18680 12909 18683
rect 12636 18652 12909 18680
rect 12897 18649 12909 18652
rect 12943 18649 12955 18683
rect 12897 18643 12955 18649
rect 12989 18683 13047 18689
rect 12989 18649 13001 18683
rect 13035 18680 13047 18683
rect 13035 18652 14504 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 10612 18584 11345 18612
rect 11333 18581 11345 18584
rect 11379 18612 11391 18615
rect 11609 18615 11667 18621
rect 11609 18612 11621 18615
rect 11379 18584 11621 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11609 18581 11621 18584
rect 11655 18612 11667 18615
rect 11974 18612 11980 18624
rect 11655 18584 11980 18612
rect 11655 18581 11667 18584
rect 11609 18575 11667 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 14476 18612 14504 18652
rect 14550 18640 14556 18692
rect 14608 18640 14614 18692
rect 16669 18683 16727 18689
rect 16669 18649 16681 18683
rect 16715 18680 16727 18683
rect 17512 18680 17540 18720
rect 18506 18708 18512 18760
rect 18564 18708 18570 18760
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 20898 18748 20904 18760
rect 18647 18720 20904 18748
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 22278 18708 22284 18760
rect 22336 18748 22342 18760
rect 24029 18751 24087 18757
rect 22336 18720 22678 18748
rect 22336 18708 22342 18720
rect 24029 18717 24041 18751
rect 24075 18748 24087 18751
rect 24118 18748 24124 18760
rect 24075 18720 24124 18748
rect 24075 18717 24087 18720
rect 24029 18711 24087 18717
rect 24118 18708 24124 18720
rect 24176 18748 24182 18760
rect 25700 18748 25728 18776
rect 24176 18720 25728 18748
rect 24176 18708 24182 18720
rect 27430 18708 27436 18760
rect 27488 18748 27494 18760
rect 27801 18751 27859 18757
rect 27801 18748 27813 18751
rect 27488 18720 27813 18748
rect 27488 18708 27494 18720
rect 27801 18717 27813 18720
rect 27847 18717 27859 18751
rect 27801 18711 27859 18717
rect 28166 18708 28172 18760
rect 28224 18748 28230 18760
rect 29104 18748 29132 18788
rect 29638 18776 29644 18788
rect 29696 18776 29702 18828
rect 29914 18776 29920 18828
rect 29972 18776 29978 18828
rect 31956 18825 31984 18856
rect 32674 18844 32680 18856
rect 32732 18844 32738 18896
rect 33226 18884 33232 18896
rect 32876 18856 33232 18884
rect 32876 18825 32904 18856
rect 33226 18844 33232 18856
rect 33284 18844 33290 18896
rect 33686 18844 33692 18896
rect 33744 18884 33750 18896
rect 35084 18884 35112 18924
rect 33744 18856 35112 18884
rect 36924 18884 36952 18924
rect 37369 18921 37381 18955
rect 37415 18952 37427 18955
rect 39390 18952 39396 18964
rect 37415 18924 39396 18952
rect 37415 18921 37427 18924
rect 37369 18915 37427 18921
rect 39390 18912 39396 18924
rect 39448 18912 39454 18964
rect 41506 18952 41512 18964
rect 39500 18924 41512 18952
rect 39500 18884 39528 18924
rect 41506 18912 41512 18924
rect 41564 18912 41570 18964
rect 42058 18912 42064 18964
rect 42116 18912 42122 18964
rect 46845 18955 46903 18961
rect 46845 18921 46857 18955
rect 46891 18952 46903 18955
rect 47486 18952 47492 18964
rect 46891 18924 47492 18952
rect 46891 18921 46903 18924
rect 46845 18915 46903 18921
rect 47486 18912 47492 18924
rect 47544 18912 47550 18964
rect 36924 18856 39528 18884
rect 33744 18844 33750 18856
rect 41874 18844 41880 18896
rect 41932 18884 41938 18896
rect 48041 18887 48099 18893
rect 48041 18884 48053 18887
rect 41932 18856 48053 18884
rect 41932 18844 41938 18856
rect 48041 18853 48053 18856
rect 48087 18853 48099 18887
rect 48041 18847 48099 18853
rect 31941 18819 31999 18825
rect 31941 18785 31953 18819
rect 31987 18785 31999 18819
rect 31941 18779 31999 18785
rect 32125 18819 32183 18825
rect 32125 18785 32137 18819
rect 32171 18785 32183 18819
rect 32125 18779 32183 18785
rect 32861 18819 32919 18825
rect 32861 18785 32873 18819
rect 32907 18785 32919 18819
rect 32861 18779 32919 18785
rect 32953 18819 33011 18825
rect 32953 18785 32965 18819
rect 32999 18816 33011 18819
rect 34146 18816 34152 18828
rect 32999 18788 34152 18816
rect 32999 18785 33011 18788
rect 32953 18779 33011 18785
rect 28224 18720 29132 18748
rect 29181 18751 29239 18757
rect 28224 18708 28230 18720
rect 29181 18717 29193 18751
rect 29227 18748 29239 18751
rect 29227 18720 32076 18748
rect 29227 18717 29239 18720
rect 29181 18711 29239 18717
rect 19334 18680 19340 18692
rect 16715 18652 17448 18680
rect 17512 18652 19340 18680
rect 16715 18649 16727 18652
rect 16669 18643 16727 18649
rect 17420 18624 17448 18652
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 19429 18683 19487 18689
rect 19429 18649 19441 18683
rect 19475 18680 19487 18683
rect 19610 18680 19616 18692
rect 19475 18652 19616 18680
rect 19475 18649 19487 18652
rect 19429 18643 19487 18649
rect 19610 18640 19616 18652
rect 19668 18640 19674 18692
rect 20257 18683 20315 18689
rect 20257 18649 20269 18683
rect 20303 18680 20315 18683
rect 20303 18652 22508 18680
rect 20303 18649 20315 18652
rect 20257 18643 20315 18649
rect 15562 18612 15568 18624
rect 14476 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15838 18572 15844 18624
rect 15896 18612 15902 18624
rect 16393 18615 16451 18621
rect 16393 18612 16405 18615
rect 15896 18584 16405 18612
rect 15896 18572 15902 18584
rect 16393 18581 16405 18584
rect 16439 18612 16451 18615
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 16439 18584 17325 18612
rect 16439 18581 16451 18584
rect 16393 18575 16451 18581
rect 17313 18581 17325 18584
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 17402 18572 17408 18624
rect 17460 18572 17466 18624
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 19521 18615 19579 18621
rect 19521 18612 19533 18615
rect 17552 18584 19533 18612
rect 17552 18572 17558 18584
rect 19521 18581 19533 18584
rect 19567 18612 19579 18615
rect 21358 18612 21364 18624
rect 19567 18584 21364 18612
rect 19567 18581 19579 18584
rect 19521 18575 19579 18581
rect 21358 18572 21364 18584
rect 21416 18612 21422 18624
rect 21453 18615 21511 18621
rect 21453 18612 21465 18615
rect 21416 18584 21465 18612
rect 21416 18572 21422 18584
rect 21453 18581 21465 18584
rect 21499 18581 21511 18615
rect 21453 18575 21511 18581
rect 21545 18615 21603 18621
rect 21545 18581 21557 18615
rect 21591 18612 21603 18615
rect 21634 18612 21640 18624
rect 21591 18584 21640 18612
rect 21591 18581 21603 18584
rect 21545 18575 21603 18581
rect 21634 18572 21640 18584
rect 21692 18572 21698 18624
rect 22480 18612 22508 18652
rect 23474 18640 23480 18692
rect 23532 18680 23538 18692
rect 23753 18683 23811 18689
rect 23753 18680 23765 18683
rect 23532 18652 23765 18680
rect 23532 18640 23538 18652
rect 23753 18649 23765 18652
rect 23799 18649 23811 18683
rect 23753 18643 23811 18649
rect 23842 18640 23848 18692
rect 23900 18680 23906 18692
rect 26053 18683 26111 18689
rect 26053 18680 26065 18683
rect 23900 18652 26065 18680
rect 23900 18640 23906 18652
rect 26053 18649 26065 18652
rect 26099 18649 26111 18683
rect 26053 18643 26111 18649
rect 26142 18640 26148 18692
rect 26200 18680 26206 18692
rect 29362 18680 29368 18692
rect 26200 18652 26542 18680
rect 27724 18652 29368 18680
rect 26200 18640 26206 18652
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 22480 18584 24593 18612
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 24762 18572 24768 18624
rect 24820 18612 24826 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24820 18584 24961 18612
rect 24820 18572 24826 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 25038 18572 25044 18624
rect 25096 18572 25102 18624
rect 25130 18572 25136 18624
rect 25188 18612 25194 18624
rect 27724 18612 27752 18652
rect 29362 18640 29368 18652
rect 29420 18640 29426 18692
rect 29822 18640 29828 18692
rect 29880 18680 29886 18692
rect 30101 18683 30159 18689
rect 30101 18680 30113 18683
rect 29880 18652 30113 18680
rect 29880 18640 29886 18652
rect 30101 18649 30113 18652
rect 30147 18649 30159 18683
rect 30742 18680 30748 18692
rect 30101 18643 30159 18649
rect 30208 18652 30748 18680
rect 25188 18584 27752 18612
rect 25188 18572 25194 18584
rect 28350 18572 28356 18624
rect 28408 18572 28414 18624
rect 28626 18572 28632 18624
rect 28684 18572 28690 18624
rect 28997 18615 29055 18621
rect 28997 18581 29009 18615
rect 29043 18612 29055 18615
rect 29178 18612 29184 18624
rect 29043 18584 29184 18612
rect 29043 18581 29055 18584
rect 28997 18575 29055 18581
rect 29178 18572 29184 18584
rect 29236 18572 29242 18624
rect 29638 18572 29644 18624
rect 29696 18612 29702 18624
rect 30009 18615 30067 18621
rect 30009 18612 30021 18615
rect 29696 18584 30021 18612
rect 29696 18572 29702 18584
rect 30009 18581 30021 18584
rect 30055 18612 30067 18615
rect 30208 18612 30236 18652
rect 30742 18640 30748 18652
rect 30800 18640 30806 18692
rect 30055 18584 30236 18612
rect 30055 18581 30067 18584
rect 30009 18575 30067 18581
rect 30466 18572 30472 18624
rect 30524 18572 30530 18624
rect 31018 18572 31024 18624
rect 31076 18612 31082 18624
rect 31113 18615 31171 18621
rect 31113 18612 31125 18615
rect 31076 18584 31125 18612
rect 31076 18572 31082 18584
rect 31113 18581 31125 18584
rect 31159 18612 31171 18615
rect 31294 18612 31300 18624
rect 31159 18584 31300 18612
rect 31159 18581 31171 18584
rect 31113 18575 31171 18581
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 31846 18572 31852 18624
rect 31904 18572 31910 18624
rect 32048 18612 32076 18720
rect 32140 18680 32168 18779
rect 32674 18708 32680 18760
rect 32732 18748 32738 18760
rect 32968 18748 32996 18779
rect 34146 18776 34152 18788
rect 34204 18776 34210 18828
rect 34514 18776 34520 18828
rect 34572 18816 34578 18828
rect 35621 18819 35679 18825
rect 35621 18816 35633 18819
rect 34572 18788 35633 18816
rect 34572 18776 34578 18788
rect 35621 18785 35633 18788
rect 35667 18785 35679 18819
rect 35621 18779 35679 18785
rect 37274 18776 37280 18828
rect 37332 18816 37338 18828
rect 37332 18788 38516 18816
rect 37332 18776 37338 18788
rect 32732 18720 32996 18748
rect 32732 18708 32738 18720
rect 33502 18708 33508 18760
rect 33560 18748 33566 18760
rect 33870 18748 33876 18760
rect 33560 18720 33876 18748
rect 33560 18708 33566 18720
rect 33870 18708 33876 18720
rect 33928 18748 33934 18760
rect 34241 18751 34299 18757
rect 34241 18748 34253 18751
rect 33928 18720 34253 18748
rect 33928 18708 33934 18720
rect 34241 18717 34253 18720
rect 34287 18717 34299 18751
rect 34241 18711 34299 18717
rect 34425 18751 34483 18757
rect 34425 18717 34437 18751
rect 34471 18748 34483 18751
rect 34606 18748 34612 18760
rect 34471 18720 34612 18748
rect 34471 18717 34483 18720
rect 34425 18711 34483 18717
rect 34606 18708 34612 18720
rect 34664 18708 34670 18760
rect 35161 18751 35219 18757
rect 35161 18717 35173 18751
rect 35207 18748 35219 18751
rect 35526 18748 35532 18760
rect 35207 18720 35532 18748
rect 35207 18717 35219 18720
rect 35161 18711 35219 18717
rect 35526 18708 35532 18720
rect 35584 18708 35590 18760
rect 38381 18751 38439 18757
rect 38381 18748 38393 18751
rect 37200 18720 38393 18748
rect 35342 18680 35348 18692
rect 32140 18652 35348 18680
rect 35342 18640 35348 18652
rect 35400 18680 35406 18692
rect 35897 18683 35955 18689
rect 35897 18680 35909 18683
rect 35400 18652 35909 18680
rect 35400 18640 35406 18652
rect 35897 18649 35909 18652
rect 35943 18649 35955 18683
rect 35897 18643 35955 18649
rect 36096 18652 36386 18680
rect 36096 18624 36124 18652
rect 32766 18612 32772 18624
rect 32048 18584 32772 18612
rect 32766 18572 32772 18584
rect 32824 18572 32830 18624
rect 32950 18572 32956 18624
rect 33008 18612 33014 18624
rect 33045 18615 33103 18621
rect 33045 18612 33057 18615
rect 33008 18584 33057 18612
rect 33008 18572 33014 18584
rect 33045 18581 33057 18584
rect 33091 18581 33103 18615
rect 33045 18575 33103 18581
rect 33413 18615 33471 18621
rect 33413 18581 33425 18615
rect 33459 18612 33471 18615
rect 33778 18612 33784 18624
rect 33459 18584 33784 18612
rect 33459 18581 33471 18584
rect 33413 18575 33471 18581
rect 33778 18572 33784 18584
rect 33836 18572 33842 18624
rect 33870 18572 33876 18624
rect 33928 18572 33934 18624
rect 36078 18572 36084 18624
rect 36136 18572 36142 18624
rect 36814 18572 36820 18624
rect 36872 18612 36878 18624
rect 37200 18612 37228 18720
rect 38381 18717 38393 18720
rect 38427 18717 38439 18751
rect 38488 18748 38516 18788
rect 38562 18776 38568 18828
rect 38620 18776 38626 18828
rect 39666 18776 39672 18828
rect 39724 18816 39730 18828
rect 41785 18819 41843 18825
rect 41785 18816 41797 18819
rect 39724 18788 41797 18816
rect 39724 18776 39730 18788
rect 41785 18785 41797 18788
rect 41831 18785 41843 18819
rect 48406 18816 48412 18828
rect 41785 18779 41843 18785
rect 47504 18788 48412 18816
rect 47504 18757 47532 18788
rect 48406 18776 48412 18788
rect 48464 18776 48470 18828
rect 47489 18751 47547 18757
rect 38488 18720 40264 18748
rect 38381 18711 38439 18717
rect 39577 18683 39635 18689
rect 39577 18680 39589 18683
rect 37660 18652 39589 18680
rect 36872 18584 37228 18612
rect 36872 18572 36878 18584
rect 37550 18572 37556 18624
rect 37608 18612 37614 18624
rect 37660 18621 37688 18652
rect 39577 18649 39589 18652
rect 39623 18680 39635 18683
rect 39666 18680 39672 18692
rect 39623 18652 39672 18680
rect 39623 18649 39635 18652
rect 39577 18643 39635 18649
rect 39666 18640 39672 18652
rect 39724 18640 39730 18692
rect 37645 18615 37703 18621
rect 37645 18612 37657 18615
rect 37608 18584 37657 18612
rect 37608 18572 37614 18584
rect 37645 18581 37657 18584
rect 37691 18581 37703 18615
rect 37645 18575 37703 18581
rect 38010 18572 38016 18624
rect 38068 18572 38074 18624
rect 38470 18572 38476 18624
rect 38528 18572 38534 18624
rect 40037 18615 40095 18621
rect 40037 18581 40049 18615
rect 40083 18612 40095 18615
rect 40126 18612 40132 18624
rect 40083 18584 40132 18612
rect 40083 18581 40095 18584
rect 40037 18575 40095 18581
rect 40126 18572 40132 18584
rect 40184 18572 40190 18624
rect 40236 18612 40264 18720
rect 47489 18717 47501 18751
rect 47535 18717 47547 18751
rect 47489 18711 47547 18717
rect 48225 18751 48283 18757
rect 48225 18717 48237 18751
rect 48271 18748 48283 18751
rect 48685 18751 48743 18757
rect 48685 18748 48697 18751
rect 48271 18720 48697 18748
rect 48271 18717 48283 18720
rect 48225 18711 48283 18717
rect 48685 18717 48697 18720
rect 48731 18717 48743 18751
rect 48685 18711 48743 18717
rect 49329 18751 49387 18757
rect 49329 18717 49341 18751
rect 49375 18748 49387 18751
rect 49418 18748 49424 18760
rect 49375 18720 49424 18748
rect 49375 18717 49387 18720
rect 49329 18711 49387 18717
rect 40494 18640 40500 18692
rect 40552 18640 40558 18692
rect 41509 18683 41567 18689
rect 41509 18649 41521 18683
rect 41555 18649 41567 18683
rect 41509 18643 41567 18649
rect 47029 18683 47087 18689
rect 47029 18649 47041 18683
rect 47075 18680 47087 18683
rect 49344 18680 49372 18711
rect 49418 18708 49424 18720
rect 49476 18708 49482 18760
rect 47075 18652 49372 18680
rect 47075 18649 47087 18652
rect 47029 18643 47087 18649
rect 41524 18612 41552 18643
rect 40236 18584 41552 18612
rect 47302 18572 47308 18624
rect 47360 18572 47366 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 3602 18368 3608 18420
rect 3660 18368 3666 18420
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 9858 18408 9864 18420
rect 9815 18380 9864 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 10410 18368 10416 18420
rect 10468 18408 10474 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 10468 18380 10793 18408
rect 10468 18368 10474 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 10781 18371 10839 18377
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 17957 18411 18015 18417
rect 17957 18408 17969 18411
rect 12492 18380 17969 18408
rect 12492 18368 12498 18380
rect 17957 18377 17969 18380
rect 18003 18377 18015 18411
rect 17957 18371 18015 18377
rect 18417 18411 18475 18417
rect 18417 18377 18429 18411
rect 18463 18408 18475 18411
rect 22097 18411 22155 18417
rect 22097 18408 22109 18411
rect 18463 18380 22109 18408
rect 18463 18377 18475 18380
rect 18417 18371 18475 18377
rect 22097 18377 22109 18380
rect 22143 18377 22155 18411
rect 22097 18371 22155 18377
rect 22465 18411 22523 18417
rect 22465 18377 22477 18411
rect 22511 18408 22523 18411
rect 25774 18408 25780 18420
rect 22511 18380 25780 18408
rect 22511 18377 22523 18380
rect 22465 18371 22523 18377
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 27246 18408 27252 18420
rect 26283 18380 27252 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27617 18411 27675 18417
rect 27617 18377 27629 18411
rect 27663 18408 27675 18411
rect 27706 18408 27712 18420
rect 27663 18380 27712 18408
rect 27663 18377 27675 18380
rect 27617 18371 27675 18377
rect 27706 18368 27712 18380
rect 27764 18368 27770 18420
rect 28721 18411 28779 18417
rect 28721 18377 28733 18411
rect 28767 18408 28779 18411
rect 30190 18408 30196 18420
rect 28767 18380 30196 18408
rect 28767 18377 28779 18380
rect 28721 18371 28779 18377
rect 30190 18368 30196 18380
rect 30248 18368 30254 18420
rect 30837 18411 30895 18417
rect 30837 18377 30849 18411
rect 30883 18408 30895 18411
rect 31202 18408 31208 18420
rect 30883 18380 31208 18408
rect 30883 18377 30895 18380
rect 30837 18371 30895 18377
rect 31202 18368 31208 18380
rect 31260 18368 31266 18420
rect 32582 18368 32588 18420
rect 32640 18368 32646 18420
rect 32766 18368 32772 18420
rect 32824 18408 32830 18420
rect 32824 18380 35204 18408
rect 32824 18368 32830 18380
rect 4522 18340 4528 18352
rect 3436 18312 4528 18340
rect 3436 18281 3464 18312
rect 4522 18300 4528 18312
rect 4580 18300 4586 18352
rect 7650 18300 7656 18352
rect 7708 18300 7714 18352
rect 11422 18340 11428 18352
rect 9968 18312 11428 18340
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18241 3019 18275
rect 2961 18235 3019 18241
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 1762 18164 1768 18216
rect 1820 18164 1826 18216
rect 2976 18068 3004 18235
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 9968 18281 9996 18312
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 13078 18300 13084 18352
rect 13136 18340 13142 18352
rect 13173 18343 13231 18349
rect 13173 18340 13185 18343
rect 13136 18312 13185 18340
rect 13136 18300 13142 18312
rect 13173 18309 13185 18312
rect 13219 18309 13231 18343
rect 13173 18303 13231 18309
rect 13538 18300 13544 18352
rect 13596 18340 13602 18352
rect 14277 18343 14335 18349
rect 14277 18340 14289 18343
rect 13596 18312 14289 18340
rect 13596 18300 13602 18312
rect 14277 18309 14289 18312
rect 14323 18309 14335 18343
rect 14277 18303 14335 18309
rect 14369 18343 14427 18349
rect 14369 18309 14381 18343
rect 14415 18340 14427 18343
rect 16758 18340 16764 18352
rect 14415 18312 16764 18340
rect 14415 18309 14427 18312
rect 14369 18303 14427 18309
rect 16758 18300 16764 18312
rect 16816 18300 16822 18352
rect 16942 18300 16948 18352
rect 17000 18300 17006 18352
rect 17494 18340 17500 18352
rect 17328 18312 17500 18340
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4120 18244 4445 18272
rect 4120 18232 4126 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18272 10931 18275
rect 11882 18272 11888 18284
rect 10919 18244 11888 18272
rect 10919 18241 10931 18244
rect 10873 18235 10931 18241
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4246 18204 4252 18216
rect 4203 18176 4252 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 7852 18136 7880 18235
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10652 18176 10977 18204
rect 10652 18164 10658 18176
rect 10965 18173 10977 18176
rect 11011 18204 11023 18207
rect 11698 18204 11704 18216
rect 11011 18176 11704 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 11974 18164 11980 18216
rect 12032 18204 12038 18216
rect 12084 18204 12112 18258
rect 13446 18232 13452 18284
rect 13504 18232 13510 18284
rect 15010 18272 15016 18284
rect 13556 18244 15016 18272
rect 13556 18204 13584 18244
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 16298 18232 16304 18284
rect 16356 18232 16362 18284
rect 17034 18232 17040 18284
rect 17092 18272 17098 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 17092 18244 17233 18272
rect 17092 18232 17098 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 12032 18176 13584 18204
rect 12032 18164 12038 18176
rect 14550 18164 14556 18216
rect 14608 18164 14614 18216
rect 14918 18164 14924 18216
rect 14976 18164 14982 18216
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16761 18207 16819 18213
rect 15703 18176 16252 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 7852 18108 11836 18136
rect 9674 18068 9680 18080
rect 2976 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 9824 18040 10425 18068
rect 9824 18028 9830 18040
rect 10413 18037 10425 18040
rect 10459 18037 10471 18071
rect 10413 18031 10471 18037
rect 11698 18028 11704 18080
rect 11756 18028 11762 18080
rect 11808 18068 11836 18108
rect 13722 18096 13728 18148
rect 13780 18136 13786 18148
rect 13909 18139 13967 18145
rect 13909 18136 13921 18139
rect 13780 18108 13921 18136
rect 13780 18096 13786 18108
rect 13909 18105 13921 18108
rect 13955 18105 13967 18139
rect 13909 18099 13967 18105
rect 15930 18096 15936 18148
rect 15988 18136 15994 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15988 18108 16129 18136
rect 15988 18096 15994 18108
rect 16117 18105 16129 18108
rect 16163 18105 16175 18139
rect 16224 18136 16252 18176
rect 16761 18173 16773 18207
rect 16807 18204 16819 18207
rect 17328 18204 17356 18312
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 19150 18340 19156 18352
rect 18616 18312 19156 18340
rect 17405 18275 17463 18281
rect 17405 18241 17417 18275
rect 17451 18241 17463 18275
rect 17405 18235 17463 18241
rect 18325 18275 18383 18281
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 18506 18272 18512 18284
rect 18371 18244 18512 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 16807 18176 17356 18204
rect 16807 18173 16819 18176
rect 16761 18167 16819 18173
rect 16666 18136 16672 18148
rect 16224 18108 16672 18136
rect 16117 18099 16175 18105
rect 16666 18096 16672 18108
rect 16724 18096 16730 18148
rect 17420 18136 17448 18235
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 18616 18213 18644 18312
rect 19150 18300 19156 18312
rect 19208 18340 19214 18352
rect 19889 18343 19947 18349
rect 19889 18340 19901 18343
rect 19208 18312 19901 18340
rect 19208 18300 19214 18312
rect 19889 18309 19901 18312
rect 19935 18309 19947 18343
rect 19889 18303 19947 18309
rect 20622 18300 20628 18352
rect 20680 18300 20686 18352
rect 22646 18300 22652 18352
rect 22704 18340 22710 18352
rect 22704 18312 23336 18340
rect 22704 18300 22710 18312
rect 21266 18232 21272 18284
rect 21324 18272 21330 18284
rect 22557 18275 22615 18281
rect 21324 18244 22094 18272
rect 21324 18232 21330 18244
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 19610 18204 19616 18216
rect 19383 18176 19616 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 22066 18136 22094 18244
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 22738 18272 22744 18284
rect 22603 18244 22744 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 22738 18232 22744 18244
rect 22796 18232 22802 18284
rect 23308 18281 23336 18312
rect 24118 18300 24124 18352
rect 24176 18300 24182 18352
rect 24486 18300 24492 18352
rect 24544 18340 24550 18352
rect 28813 18343 28871 18349
rect 24544 18312 25452 18340
rect 24544 18300 24550 18312
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 23382 18272 23388 18284
rect 23339 18244 23388 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 24670 18232 24676 18284
rect 24728 18272 24734 18284
rect 25041 18275 25099 18281
rect 25041 18272 25053 18275
rect 24728 18244 25053 18272
rect 24728 18232 24734 18244
rect 25041 18241 25053 18244
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 22649 18207 22707 18213
rect 22649 18173 22661 18207
rect 22695 18173 22707 18207
rect 22649 18167 22707 18173
rect 22664 18136 22692 18167
rect 25314 18164 25320 18216
rect 25372 18164 25378 18216
rect 25424 18204 25452 18312
rect 26528 18312 28580 18340
rect 26329 18275 26387 18281
rect 26329 18241 26341 18275
rect 26375 18272 26387 18275
rect 26528 18272 26556 18312
rect 26375 18244 26556 18272
rect 27525 18275 27583 18281
rect 26375 18241 26387 18244
rect 26329 18235 26387 18241
rect 27525 18241 27537 18275
rect 27571 18272 27583 18275
rect 28552 18272 28580 18312
rect 28813 18309 28825 18343
rect 28859 18340 28871 18343
rect 32122 18340 32128 18352
rect 28859 18312 32128 18340
rect 28859 18309 28871 18312
rect 28813 18303 28871 18309
rect 32122 18300 32128 18312
rect 32180 18300 32186 18352
rect 33226 18300 33232 18352
rect 33284 18340 33290 18352
rect 33962 18340 33968 18352
rect 33284 18312 33968 18340
rect 33284 18300 33290 18312
rect 33962 18300 33968 18312
rect 34020 18300 34026 18352
rect 35176 18340 35204 18380
rect 35342 18368 35348 18420
rect 35400 18368 35406 18420
rect 35897 18411 35955 18417
rect 35897 18377 35909 18411
rect 35943 18377 35955 18411
rect 35897 18371 35955 18377
rect 35912 18340 35940 18371
rect 37182 18368 37188 18420
rect 37240 18408 37246 18420
rect 40405 18411 40463 18417
rect 40405 18408 40417 18411
rect 37240 18380 40417 18408
rect 37240 18368 37246 18380
rect 40405 18377 40417 18380
rect 40451 18377 40463 18411
rect 40405 18371 40463 18377
rect 40862 18368 40868 18420
rect 40920 18368 40926 18420
rect 47673 18411 47731 18417
rect 47673 18377 47685 18411
rect 47719 18408 47731 18411
rect 48406 18408 48412 18420
rect 47719 18380 48412 18408
rect 47719 18377 47731 18380
rect 47673 18371 47731 18377
rect 48406 18368 48412 18380
rect 48464 18368 48470 18420
rect 35176 18312 35940 18340
rect 36078 18300 36084 18352
rect 36136 18340 36142 18352
rect 36136 18312 37044 18340
rect 36136 18300 36142 18312
rect 30098 18272 30104 18284
rect 27571 18244 28488 18272
rect 28552 18244 30104 18272
rect 27571 18241 27583 18244
rect 27525 18235 27583 18241
rect 26421 18207 26479 18213
rect 26421 18204 26433 18207
rect 25424 18176 26433 18204
rect 26421 18173 26433 18176
rect 26467 18173 26479 18207
rect 26421 18167 26479 18173
rect 26694 18164 26700 18216
rect 26752 18204 26758 18216
rect 27709 18207 27767 18213
rect 27709 18204 27721 18207
rect 26752 18176 27721 18204
rect 26752 18164 26758 18176
rect 27709 18173 27721 18176
rect 27755 18173 27767 18207
rect 27709 18167 27767 18173
rect 17420 18108 19748 18136
rect 22066 18108 22692 18136
rect 13538 18068 13544 18080
rect 11808 18040 13544 18068
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 15197 18071 15255 18077
rect 15197 18037 15209 18071
rect 15243 18068 15255 18071
rect 15286 18068 15292 18080
rect 15243 18040 15292 18068
rect 15243 18037 15255 18040
rect 15197 18031 15255 18037
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 18969 18071 19027 18077
rect 18969 18068 18981 18071
rect 18656 18040 18981 18068
rect 18656 18028 18662 18040
rect 18969 18037 18981 18040
rect 19015 18037 19027 18071
rect 19720 18068 19748 18108
rect 23658 18096 23664 18148
rect 23716 18136 23722 18148
rect 24673 18139 24731 18145
rect 24673 18136 24685 18139
rect 23716 18108 24685 18136
rect 23716 18096 23722 18108
rect 24673 18105 24685 18108
rect 24719 18105 24731 18139
rect 24673 18099 24731 18105
rect 24780 18108 26004 18136
rect 21174 18068 21180 18080
rect 19720 18040 21180 18068
rect 18969 18031 19027 18037
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21450 18068 21456 18080
rect 21407 18040 21456 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 22462 18028 22468 18080
rect 22520 18068 22526 18080
rect 24780 18068 24808 18108
rect 22520 18040 24808 18068
rect 22520 18028 22526 18040
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25869 18071 25927 18077
rect 25869 18068 25881 18071
rect 25096 18040 25881 18068
rect 25096 18028 25102 18040
rect 25869 18037 25881 18040
rect 25915 18037 25927 18071
rect 25976 18068 26004 18108
rect 26050 18096 26056 18148
rect 26108 18136 26114 18148
rect 28353 18139 28411 18145
rect 28353 18136 28365 18139
rect 26108 18108 28365 18136
rect 26108 18096 26114 18108
rect 28353 18105 28365 18108
rect 28399 18105 28411 18139
rect 28460 18136 28488 18244
rect 30098 18232 30104 18244
rect 30156 18232 30162 18284
rect 30377 18275 30435 18281
rect 30377 18272 30389 18275
rect 30208 18244 30389 18272
rect 28902 18164 28908 18216
rect 28960 18164 28966 18216
rect 30208 18204 30236 18244
rect 30377 18241 30389 18244
rect 30423 18241 30435 18275
rect 30377 18235 30435 18241
rect 30469 18275 30527 18281
rect 30469 18241 30481 18275
rect 30515 18272 30527 18275
rect 31297 18275 31355 18281
rect 31297 18272 31309 18275
rect 30515 18244 31309 18272
rect 30515 18241 30527 18244
rect 30469 18235 30527 18241
rect 31297 18241 31309 18244
rect 31343 18241 31355 18275
rect 31297 18235 31355 18241
rect 32030 18232 32036 18284
rect 32088 18272 32094 18284
rect 32677 18275 32735 18281
rect 32677 18272 32689 18275
rect 32088 18244 32689 18272
rect 32088 18232 32094 18244
rect 32677 18241 32689 18244
rect 32723 18272 32735 18275
rect 33134 18272 33140 18284
rect 32723 18244 33140 18272
rect 32723 18241 32735 18244
rect 32677 18235 32735 18241
rect 33134 18232 33140 18244
rect 33192 18232 33198 18284
rect 35250 18272 35256 18284
rect 35006 18244 35256 18272
rect 35250 18232 35256 18244
rect 35308 18272 35314 18284
rect 36096 18272 36124 18300
rect 35308 18244 36124 18272
rect 35308 18232 35314 18244
rect 36262 18232 36268 18284
rect 36320 18232 36326 18284
rect 36357 18275 36415 18281
rect 36357 18241 36369 18275
rect 36403 18272 36415 18275
rect 36906 18272 36912 18284
rect 36403 18244 36912 18272
rect 36403 18241 36415 18244
rect 36357 18235 36415 18241
rect 36906 18232 36912 18244
rect 36964 18232 36970 18284
rect 37016 18272 37044 18312
rect 37274 18300 37280 18352
rect 37332 18340 37338 18352
rect 38010 18340 38016 18352
rect 37332 18312 38016 18340
rect 37332 18300 37338 18312
rect 38010 18300 38016 18312
rect 38068 18300 38074 18352
rect 40773 18343 40831 18349
rect 40773 18309 40785 18343
rect 40819 18340 40831 18343
rect 47302 18340 47308 18352
rect 40819 18312 47308 18340
rect 40819 18309 40831 18312
rect 40773 18303 40831 18309
rect 47302 18300 47308 18312
rect 47360 18300 47366 18352
rect 37461 18275 37519 18281
rect 37461 18272 37473 18275
rect 37016 18244 37473 18272
rect 37461 18241 37473 18244
rect 37507 18272 37519 18275
rect 38378 18272 38384 18284
rect 37507 18244 38384 18272
rect 37507 18241 37519 18244
rect 37461 18235 37519 18241
rect 38378 18232 38384 18244
rect 38436 18232 38442 18284
rect 39758 18232 39764 18284
rect 39816 18232 39822 18284
rect 48225 18275 48283 18281
rect 48225 18241 48237 18275
rect 48271 18272 48283 18275
rect 48685 18275 48743 18281
rect 48685 18272 48697 18275
rect 48271 18244 48697 18272
rect 48271 18241 48283 18244
rect 48225 18235 48283 18241
rect 48685 18241 48697 18244
rect 48731 18241 48743 18275
rect 48685 18235 48743 18241
rect 49326 18232 49332 18284
rect 49384 18232 49390 18284
rect 29748 18176 30236 18204
rect 28994 18136 29000 18148
rect 28460 18108 29000 18136
rect 28353 18099 28411 18105
rect 28994 18096 29000 18108
rect 29052 18136 29058 18148
rect 29270 18136 29276 18148
rect 29052 18108 29276 18136
rect 29052 18096 29058 18108
rect 29270 18096 29276 18108
rect 29328 18096 29334 18148
rect 26326 18068 26332 18080
rect 25976 18040 26332 18068
rect 25869 18031 25927 18037
rect 26326 18028 26332 18040
rect 26384 18028 26390 18080
rect 27154 18028 27160 18080
rect 27212 18028 27218 18080
rect 28258 18028 28264 18080
rect 28316 18068 28322 18080
rect 28902 18068 28908 18080
rect 28316 18040 28908 18068
rect 28316 18028 28322 18040
rect 28902 18028 28908 18040
rect 28960 18028 28966 18080
rect 29638 18028 29644 18080
rect 29696 18068 29702 18080
rect 29748 18077 29776 18176
rect 30282 18164 30288 18216
rect 30340 18164 30346 18216
rect 32490 18164 32496 18216
rect 32548 18164 32554 18216
rect 33594 18164 33600 18216
rect 33652 18164 33658 18216
rect 33870 18164 33876 18216
rect 33928 18164 33934 18216
rect 36541 18207 36599 18213
rect 36541 18173 36553 18207
rect 36587 18204 36599 18207
rect 37734 18204 37740 18216
rect 36587 18176 37740 18204
rect 36587 18173 36599 18176
rect 36541 18167 36599 18173
rect 37734 18164 37740 18176
rect 37792 18164 37798 18216
rect 37826 18164 37832 18216
rect 37884 18204 37890 18216
rect 39485 18207 39543 18213
rect 39485 18204 39497 18207
rect 37884 18176 39497 18204
rect 37884 18164 37890 18176
rect 39485 18173 39497 18176
rect 39531 18204 39543 18207
rect 40957 18207 41015 18213
rect 40957 18204 40969 18207
rect 39531 18176 40969 18204
rect 39531 18173 39543 18176
rect 39485 18167 39543 18173
rect 40957 18173 40969 18176
rect 41003 18173 41015 18207
rect 40957 18167 41015 18173
rect 47397 18207 47455 18213
rect 47397 18173 47409 18207
rect 47443 18204 47455 18207
rect 49344 18204 49372 18232
rect 47443 18176 49372 18204
rect 47443 18173 47455 18176
rect 47397 18167 47455 18173
rect 30006 18096 30012 18148
rect 30064 18136 30070 18148
rect 33410 18136 33416 18148
rect 30064 18108 33416 18136
rect 30064 18096 30070 18108
rect 33410 18096 33416 18108
rect 33468 18096 33474 18148
rect 36998 18096 37004 18148
rect 37056 18096 37062 18148
rect 37369 18139 37427 18145
rect 37369 18105 37381 18139
rect 37415 18136 37427 18139
rect 37550 18136 37556 18148
rect 37415 18108 37556 18136
rect 37415 18105 37427 18108
rect 37369 18099 37427 18105
rect 37550 18096 37556 18108
rect 37608 18096 37614 18148
rect 38010 18096 38016 18148
rect 38068 18096 38074 18148
rect 29733 18071 29791 18077
rect 29733 18068 29745 18071
rect 29696 18040 29745 18068
rect 29696 18028 29702 18040
rect 29733 18037 29745 18040
rect 29779 18037 29791 18071
rect 29733 18031 29791 18037
rect 30742 18028 30748 18080
rect 30800 18068 30806 18080
rect 32950 18068 32956 18080
rect 30800 18040 32956 18068
rect 30800 18028 30806 18040
rect 32950 18028 32956 18040
rect 33008 18028 33014 18080
rect 33045 18071 33103 18077
rect 33045 18037 33057 18071
rect 33091 18068 33103 18071
rect 35894 18068 35900 18080
rect 33091 18040 35900 18068
rect 33091 18037 33103 18040
rect 33045 18031 33103 18037
rect 35894 18028 35900 18040
rect 35952 18028 35958 18080
rect 36722 18028 36728 18080
rect 36780 18068 36786 18080
rect 37645 18071 37703 18077
rect 37645 18068 37657 18071
rect 36780 18040 37657 18068
rect 36780 18028 36786 18040
rect 37645 18037 37657 18040
rect 37691 18037 37703 18071
rect 37645 18031 37703 18037
rect 40034 18028 40040 18080
rect 40092 18068 40098 18080
rect 40494 18068 40500 18080
rect 40092 18040 40500 18068
rect 40092 18028 40098 18040
rect 40494 18028 40500 18040
rect 40552 18028 40558 18080
rect 48038 18028 48044 18080
rect 48096 18028 48102 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 10137 17867 10195 17873
rect 10137 17833 10149 17867
rect 10183 17864 10195 17867
rect 10226 17864 10232 17876
rect 10183 17836 10232 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 10594 17824 10600 17876
rect 10652 17824 10658 17876
rect 12434 17864 12440 17876
rect 10704 17836 12440 17864
rect 3326 17756 3332 17808
rect 3384 17796 3390 17808
rect 10704 17796 10732 17836
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12584 17836 12909 17864
rect 12584 17824 12590 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 12897 17827 12955 17833
rect 14277 17867 14335 17873
rect 14277 17833 14289 17867
rect 14323 17864 14335 17867
rect 14550 17864 14556 17876
rect 14323 17836 14556 17864
rect 14323 17833 14335 17836
rect 14277 17827 14335 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15102 17824 15108 17876
rect 15160 17864 15166 17876
rect 16574 17864 16580 17876
rect 15160 17836 16580 17864
rect 15160 17824 15166 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17276 17836 17509 17864
rect 17276 17824 17282 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17497 17827 17555 17833
rect 19426 17824 19432 17876
rect 19484 17824 19490 17876
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 21082 17864 21088 17876
rect 19668 17836 21088 17864
rect 19668 17824 19674 17836
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 21174 17824 21180 17876
rect 21232 17864 21238 17876
rect 21232 17836 21956 17864
rect 21232 17824 21238 17836
rect 19518 17796 19524 17808
rect 3384 17768 10732 17796
rect 15948 17768 19524 17796
rect 3384 17756 3390 17768
rect 12345 17731 12403 17737
rect 12345 17697 12357 17731
rect 12391 17728 12403 17731
rect 12526 17728 12532 17740
rect 12391 17700 12532 17728
rect 12391 17697 12403 17700
rect 12345 17691 12403 17697
rect 12526 17688 12532 17700
rect 12584 17728 12590 17740
rect 13446 17728 13452 17740
rect 12584 17700 13452 17728
rect 12584 17688 12590 17700
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 15948 17728 15976 17768
rect 19518 17756 19524 17768
rect 19576 17756 19582 17808
rect 13740 17700 15976 17728
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 10410 17660 10416 17672
rect 3007 17632 10416 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 13740 17669 13768 17700
rect 16022 17688 16028 17740
rect 16080 17728 16086 17740
rect 16390 17728 16396 17740
rect 16080 17700 16396 17728
rect 16080 17688 16086 17700
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 16945 17731 17003 17737
rect 16945 17697 16957 17731
rect 16991 17728 17003 17731
rect 17310 17728 17316 17740
rect 16991 17700 17316 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 19628 17728 19656 17824
rect 21928 17796 21956 17836
rect 23290 17824 23296 17876
rect 23348 17824 23354 17876
rect 23566 17824 23572 17876
rect 23624 17864 23630 17876
rect 25777 17867 25835 17873
rect 25777 17864 25789 17867
rect 23624 17836 25789 17864
rect 23624 17824 23630 17836
rect 25777 17833 25789 17836
rect 25823 17833 25835 17867
rect 29270 17864 29276 17876
rect 25777 17827 25835 17833
rect 25976 17836 29276 17864
rect 24581 17799 24639 17805
rect 24581 17796 24593 17799
rect 21928 17768 24593 17796
rect 24581 17765 24593 17768
rect 24627 17765 24639 17799
rect 24581 17759 24639 17765
rect 21634 17728 21640 17740
rect 18831 17700 19656 17728
rect 20456 17700 21640 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 1026 17552 1032 17604
rect 1084 17592 1090 17604
rect 1765 17595 1823 17601
rect 1765 17592 1777 17595
rect 1084 17564 1777 17592
rect 1084 17552 1090 17564
rect 1765 17561 1777 17564
rect 1811 17561 1823 17595
rect 11638 17564 11744 17592
rect 1765 17555 1823 17561
rect 10318 17484 10324 17536
rect 10376 17484 10382 17536
rect 11716 17524 11744 17564
rect 11790 17552 11796 17604
rect 11848 17592 11854 17604
rect 12066 17592 12072 17604
rect 11848 17564 12072 17592
rect 11848 17552 11854 17564
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 13096 17592 13124 17623
rect 16666 17620 16672 17672
rect 16724 17660 16730 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 16724 17632 17141 17660
rect 16724 17620 16730 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 17770 17620 17776 17672
rect 17828 17660 17834 17672
rect 18414 17660 18420 17672
rect 17828 17632 18420 17660
rect 17828 17620 17834 17632
rect 18414 17620 18420 17632
rect 18472 17660 18478 17672
rect 19613 17663 19671 17669
rect 18472 17632 19380 17660
rect 18472 17620 18478 17632
rect 13998 17592 14004 17604
rect 13096 17564 14004 17592
rect 13998 17552 14004 17564
rect 14056 17552 14062 17604
rect 15010 17552 15016 17604
rect 15068 17552 15074 17604
rect 15749 17595 15807 17601
rect 15749 17561 15761 17595
rect 15795 17592 15807 17595
rect 16022 17592 16028 17604
rect 15795 17564 16028 17592
rect 15795 17561 15807 17564
rect 15749 17555 15807 17561
rect 16022 17552 16028 17564
rect 16080 17552 16086 17604
rect 17037 17595 17095 17601
rect 17037 17561 17049 17595
rect 17083 17592 17095 17595
rect 17494 17592 17500 17604
rect 17083 17564 17500 17592
rect 17083 17561 17095 17564
rect 17037 17555 17095 17561
rect 17494 17552 17500 17564
rect 17552 17552 17558 17604
rect 17957 17595 18015 17601
rect 17957 17561 17969 17595
rect 18003 17592 18015 17595
rect 18598 17592 18604 17604
rect 18003 17564 18604 17592
rect 18003 17561 18015 17564
rect 17957 17555 18015 17561
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 19352 17592 19380 17632
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 20346 17660 20352 17672
rect 19659 17632 20352 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20456 17592 20484 17700
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 21726 17688 21732 17740
rect 21784 17688 21790 17740
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22094 17728 22100 17740
rect 22051 17700 22100 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 23750 17688 23756 17740
rect 23808 17688 23814 17740
rect 23937 17731 23995 17737
rect 23937 17697 23949 17731
rect 23983 17728 23995 17731
rect 24946 17728 24952 17740
rect 23983 17700 24952 17728
rect 23983 17697 23995 17700
rect 23937 17691 23995 17697
rect 24946 17688 24952 17700
rect 25004 17688 25010 17740
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17697 25191 17731
rect 25133 17691 25191 17697
rect 22278 17620 22284 17672
rect 22336 17620 22342 17672
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 25148 17660 25176 17691
rect 25976 17669 26004 17836
rect 29270 17824 29276 17836
rect 29328 17824 29334 17876
rect 29546 17824 29552 17876
rect 29604 17824 29610 17876
rect 33410 17824 33416 17876
rect 33468 17864 33474 17876
rect 34425 17867 34483 17873
rect 34425 17864 34437 17867
rect 33468 17836 34437 17864
rect 33468 17824 33474 17836
rect 34425 17833 34437 17836
rect 34471 17833 34483 17867
rect 34425 17827 34483 17833
rect 35526 17824 35532 17876
rect 35584 17864 35590 17876
rect 36170 17864 36176 17876
rect 35584 17836 36176 17864
rect 35584 17824 35590 17836
rect 36170 17824 36176 17836
rect 36228 17824 36234 17876
rect 37295 17867 37353 17873
rect 37295 17833 37307 17867
rect 37341 17864 37353 17867
rect 37642 17864 37648 17876
rect 37341 17836 37648 17864
rect 37341 17833 37353 17836
rect 37295 17827 37353 17833
rect 37642 17824 37648 17836
rect 37700 17824 37706 17876
rect 38470 17824 38476 17876
rect 38528 17864 38534 17876
rect 40497 17867 40555 17873
rect 40497 17864 40509 17867
rect 38528 17836 40509 17864
rect 38528 17824 38534 17836
rect 40497 17833 40509 17836
rect 40543 17833 40555 17867
rect 40497 17827 40555 17833
rect 28902 17756 28908 17808
rect 28960 17796 28966 17808
rect 29178 17796 29184 17808
rect 28960 17768 29184 17796
rect 28960 17756 28966 17768
rect 29178 17756 29184 17768
rect 29236 17756 29242 17808
rect 32674 17796 32680 17808
rect 31404 17768 32680 17796
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 31404 17728 31432 17768
rect 32674 17756 32680 17768
rect 32732 17756 32738 17808
rect 33965 17799 34023 17805
rect 33965 17796 33977 17799
rect 32968 17768 33977 17796
rect 26200 17700 31432 17728
rect 26200 17688 26206 17700
rect 31478 17688 31484 17740
rect 31536 17688 31542 17740
rect 32968 17737 32996 17768
rect 33965 17765 33977 17768
rect 34011 17796 34023 17799
rect 35066 17796 35072 17808
rect 34011 17768 35072 17796
rect 34011 17765 34023 17768
rect 33965 17759 34023 17765
rect 35066 17756 35072 17768
rect 35124 17796 35130 17808
rect 35250 17796 35256 17808
rect 35124 17768 35256 17796
rect 35124 17756 35130 17768
rect 35250 17756 35256 17768
rect 35308 17756 35314 17808
rect 37476 17768 38654 17796
rect 32953 17731 33011 17737
rect 32953 17697 32965 17731
rect 32999 17697 33011 17731
rect 32953 17691 33011 17697
rect 33045 17731 33103 17737
rect 33045 17697 33057 17731
rect 33091 17728 33103 17731
rect 33318 17728 33324 17740
rect 33091 17700 33324 17728
rect 33091 17697 33103 17700
rect 33045 17691 33103 17697
rect 33318 17688 33324 17700
rect 33376 17688 33382 17740
rect 33873 17731 33931 17737
rect 33873 17697 33885 17731
rect 33919 17728 33931 17731
rect 37476 17728 37504 17768
rect 33919 17700 37504 17728
rect 33919 17697 33931 17700
rect 33873 17691 33931 17697
rect 23532 17632 25176 17660
rect 25961 17663 26019 17669
rect 23532 17620 23538 17632
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 26234 17620 26240 17672
rect 26292 17620 26298 17672
rect 27430 17620 27436 17672
rect 27488 17620 27494 17672
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17660 28871 17663
rect 28902 17660 28908 17672
rect 28859 17632 28908 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 28902 17620 28908 17632
rect 28960 17660 28966 17672
rect 30653 17663 30711 17669
rect 30653 17660 30665 17663
rect 28960 17632 30665 17660
rect 28960 17628 28994 17632
rect 30653 17629 30665 17632
rect 30699 17660 30711 17663
rect 31386 17660 31392 17672
rect 30699 17632 31392 17660
rect 30699 17629 30711 17632
rect 28960 17620 28966 17628
rect 30653 17623 30711 17629
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 31573 17663 31631 17669
rect 31573 17629 31585 17663
rect 31619 17660 31631 17663
rect 31754 17660 31760 17672
rect 31619 17632 31760 17660
rect 31619 17629 31631 17632
rect 31573 17623 31631 17629
rect 31754 17620 31760 17632
rect 31812 17660 31818 17672
rect 33888 17660 33916 17691
rect 37642 17688 37648 17740
rect 37700 17728 37706 17740
rect 38105 17731 38163 17737
rect 38105 17728 38117 17731
rect 37700 17700 38117 17728
rect 37700 17688 37706 17700
rect 38105 17697 38117 17700
rect 38151 17697 38163 17731
rect 38105 17691 38163 17697
rect 31812 17632 33916 17660
rect 31812 17620 31818 17632
rect 36170 17620 36176 17672
rect 36228 17620 36234 17672
rect 37550 17620 37556 17672
rect 37608 17620 37614 17672
rect 38626 17660 38654 17768
rect 46934 17756 46940 17808
rect 46992 17796 46998 17808
rect 48041 17799 48099 17805
rect 48041 17796 48053 17799
rect 46992 17768 48053 17796
rect 46992 17756 46998 17768
rect 48041 17765 48053 17768
rect 48087 17765 48099 17799
rect 48041 17759 48099 17765
rect 40678 17688 40684 17740
rect 40736 17728 40742 17740
rect 40957 17731 41015 17737
rect 40957 17728 40969 17731
rect 40736 17700 40969 17728
rect 40736 17688 40742 17700
rect 40957 17697 40969 17700
rect 41003 17697 41015 17731
rect 40957 17691 41015 17697
rect 41049 17731 41107 17737
rect 41049 17697 41061 17731
rect 41095 17697 41107 17731
rect 41049 17691 41107 17697
rect 38626 17632 40724 17660
rect 19352 17564 20484 17592
rect 20714 17552 20720 17604
rect 20772 17552 20778 17604
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 22833 17595 22891 17601
rect 21692 17564 22784 17592
rect 21692 17552 21698 17564
rect 11974 17524 11980 17536
rect 11716 17496 11980 17524
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 13538 17484 13544 17536
rect 13596 17484 13602 17536
rect 16482 17484 16488 17536
rect 16540 17484 16546 17536
rect 18782 17484 18788 17536
rect 18840 17524 18846 17536
rect 20257 17527 20315 17533
rect 20257 17524 20269 17527
rect 18840 17496 20269 17524
rect 18840 17484 18846 17496
rect 20257 17493 20269 17496
rect 20303 17524 20315 17527
rect 22554 17524 22560 17536
rect 20303 17496 22560 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 22756 17524 22784 17564
rect 22833 17561 22845 17595
rect 22879 17592 22891 17595
rect 23661 17595 23719 17601
rect 23661 17592 23673 17595
rect 22879 17564 23673 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 23661 17561 23673 17564
rect 23707 17561 23719 17595
rect 25130 17592 25136 17604
rect 23661 17555 23719 17561
rect 23768 17564 25136 17592
rect 23768 17524 23796 17564
rect 25130 17552 25136 17564
rect 25188 17552 25194 17604
rect 25222 17552 25228 17604
rect 25280 17592 25286 17604
rect 25280 17564 27108 17592
rect 25280 17552 25286 17564
rect 27080 17536 27108 17564
rect 28442 17552 28448 17604
rect 28500 17592 28506 17604
rect 28537 17595 28595 17601
rect 28537 17592 28549 17595
rect 28500 17564 28549 17592
rect 28500 17552 28506 17564
rect 28537 17561 28549 17564
rect 28583 17561 28595 17595
rect 28537 17555 28595 17561
rect 29178 17552 29184 17604
rect 29236 17592 29242 17604
rect 29365 17595 29423 17601
rect 29365 17592 29377 17595
rect 29236 17564 29377 17592
rect 29236 17552 29242 17564
rect 29365 17561 29377 17564
rect 29411 17592 29423 17595
rect 29917 17595 29975 17601
rect 29917 17592 29929 17595
rect 29411 17564 29929 17592
rect 29411 17561 29423 17564
rect 29365 17555 29423 17561
rect 29917 17561 29929 17564
rect 29963 17592 29975 17595
rect 30098 17592 30104 17604
rect 29963 17564 30104 17592
rect 29963 17561 29975 17564
rect 29917 17555 29975 17561
rect 30098 17552 30104 17564
rect 30156 17592 30162 17604
rect 30374 17592 30380 17604
rect 30156 17564 30380 17592
rect 30156 17552 30162 17564
rect 30374 17552 30380 17564
rect 30432 17552 30438 17604
rect 31662 17552 31668 17604
rect 31720 17552 31726 17604
rect 32398 17592 32404 17604
rect 32048 17564 32404 17592
rect 22756 17496 23796 17524
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24728 17496 24961 17524
rect 24728 17484 24734 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 25038 17484 25044 17536
rect 25096 17524 25102 17536
rect 26421 17527 26479 17533
rect 26421 17524 26433 17527
rect 25096 17496 26433 17524
rect 25096 17484 25102 17496
rect 26421 17493 26433 17496
rect 26467 17524 26479 17527
rect 26602 17524 26608 17536
rect 26467 17496 26608 17524
rect 26467 17493 26479 17496
rect 26421 17487 26479 17493
rect 26602 17484 26608 17496
rect 26660 17484 26666 17536
rect 27062 17484 27068 17536
rect 27120 17524 27126 17536
rect 28258 17524 28264 17536
rect 27120 17496 28264 17524
rect 27120 17484 27126 17496
rect 28258 17484 28264 17496
rect 28316 17484 28322 17536
rect 29086 17484 29092 17536
rect 29144 17484 29150 17536
rect 32048 17533 32076 17564
rect 32398 17552 32404 17564
rect 32456 17552 32462 17604
rect 40586 17592 40592 17604
rect 38764 17564 40592 17592
rect 32033 17527 32091 17533
rect 32033 17493 32045 17527
rect 32079 17493 32091 17527
rect 32033 17487 32091 17493
rect 32122 17484 32128 17536
rect 32180 17524 32186 17536
rect 32309 17527 32367 17533
rect 32309 17524 32321 17527
rect 32180 17496 32321 17524
rect 32180 17484 32186 17496
rect 32309 17493 32321 17496
rect 32355 17493 32367 17527
rect 32309 17487 32367 17493
rect 33137 17527 33195 17533
rect 33137 17493 33149 17527
rect 33183 17524 33195 17527
rect 33410 17524 33416 17536
rect 33183 17496 33416 17524
rect 33183 17493 33195 17496
rect 33137 17487 33195 17493
rect 33410 17484 33416 17496
rect 33468 17484 33474 17536
rect 33505 17527 33563 17533
rect 33505 17493 33517 17527
rect 33551 17524 33563 17527
rect 33686 17524 33692 17536
rect 33551 17496 33692 17524
rect 33551 17493 33563 17496
rect 33505 17487 33563 17493
rect 33686 17484 33692 17496
rect 33744 17484 33750 17536
rect 34333 17527 34391 17533
rect 34333 17493 34345 17527
rect 34379 17524 34391 17527
rect 34422 17524 34428 17536
rect 34379 17496 34428 17524
rect 34379 17493 34391 17496
rect 34333 17487 34391 17493
rect 34422 17484 34428 17496
rect 34480 17484 34486 17536
rect 35066 17484 35072 17536
rect 35124 17484 35130 17536
rect 35434 17484 35440 17536
rect 35492 17484 35498 17536
rect 35526 17484 35532 17536
rect 35584 17524 35590 17536
rect 35805 17527 35863 17533
rect 35805 17524 35817 17527
rect 35584 17496 35817 17524
rect 35584 17484 35590 17496
rect 35805 17493 35817 17496
rect 35851 17493 35863 17527
rect 35805 17487 35863 17493
rect 36630 17484 36636 17536
rect 36688 17524 36694 17536
rect 38289 17527 38347 17533
rect 38289 17524 38301 17527
rect 36688 17496 38301 17524
rect 36688 17484 36694 17496
rect 38289 17493 38301 17496
rect 38335 17493 38347 17527
rect 38289 17487 38347 17493
rect 38378 17484 38384 17536
rect 38436 17484 38442 17536
rect 38764 17533 38792 17564
rect 40586 17552 40592 17564
rect 40644 17552 40650 17604
rect 38749 17527 38807 17533
rect 38749 17493 38761 17527
rect 38795 17493 38807 17527
rect 38749 17487 38807 17493
rect 38930 17484 38936 17536
rect 38988 17524 38994 17536
rect 39025 17527 39083 17533
rect 39025 17524 39037 17527
rect 38988 17496 39037 17524
rect 38988 17484 38994 17496
rect 39025 17493 39037 17496
rect 39071 17493 39083 17527
rect 39025 17487 39083 17493
rect 39114 17484 39120 17536
rect 39172 17524 39178 17536
rect 39209 17527 39267 17533
rect 39209 17524 39221 17527
rect 39172 17496 39221 17524
rect 39172 17484 39178 17496
rect 39209 17493 39221 17496
rect 39255 17524 39267 17527
rect 40034 17524 40040 17536
rect 39255 17496 40040 17524
rect 39255 17493 39267 17496
rect 39209 17487 39267 17493
rect 40034 17484 40040 17496
rect 40092 17484 40098 17536
rect 40696 17524 40724 17632
rect 40770 17620 40776 17672
rect 40828 17660 40834 17672
rect 41064 17660 41092 17691
rect 40828 17632 41092 17660
rect 48225 17663 48283 17669
rect 40828 17620 40834 17632
rect 48225 17629 48237 17663
rect 48271 17660 48283 17663
rect 48685 17663 48743 17669
rect 48685 17660 48697 17663
rect 48271 17632 48697 17660
rect 48271 17629 48283 17632
rect 48225 17623 48283 17629
rect 48685 17629 48697 17632
rect 48731 17629 48743 17663
rect 48685 17623 48743 17629
rect 49326 17620 49332 17672
rect 49384 17620 49390 17672
rect 40865 17595 40923 17601
rect 40865 17561 40877 17595
rect 40911 17592 40923 17595
rect 47026 17592 47032 17604
rect 40911 17564 47032 17592
rect 40911 17561 40923 17564
rect 40865 17555 40923 17561
rect 47026 17552 47032 17564
rect 47084 17552 47090 17604
rect 47489 17595 47547 17601
rect 47489 17561 47501 17595
rect 47535 17592 47547 17595
rect 49344 17592 49372 17620
rect 47535 17564 49372 17592
rect 47535 17561 47547 17564
rect 47489 17555 47547 17561
rect 43438 17524 43444 17536
rect 40696 17496 43444 17524
rect 43438 17484 43444 17496
rect 43496 17484 43502 17536
rect 47670 17484 47676 17536
rect 47728 17484 47734 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 11793 17323 11851 17329
rect 11793 17320 11805 17323
rect 7432 17292 11805 17320
rect 7432 17280 7438 17292
rect 11793 17289 11805 17292
rect 11839 17289 11851 17323
rect 11793 17283 11851 17289
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 12492 17292 14197 17320
rect 12492 17280 12498 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 17092 17292 17417 17320
rect 17092 17280 17098 17292
rect 17405 17289 17417 17292
rect 17451 17289 17463 17323
rect 17405 17283 17463 17289
rect 19150 17280 19156 17332
rect 19208 17280 19214 17332
rect 22554 17320 22560 17332
rect 19306 17292 22560 17320
rect 10318 17212 10324 17264
rect 10376 17252 10382 17264
rect 11885 17255 11943 17261
rect 11885 17252 11897 17255
rect 10376 17224 11897 17252
rect 10376 17212 10382 17224
rect 11885 17221 11897 17224
rect 11931 17221 11943 17255
rect 11885 17215 11943 17221
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 4338 17184 4344 17196
rect 3007 17156 4344 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 5810 17144 5816 17196
rect 5868 17184 5874 17196
rect 9858 17184 9864 17196
rect 5868 17156 9864 17184
rect 5868 17144 5874 17156
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10008 17156 10793 17184
rect 10008 17144 10014 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 11900 17184 11928 17215
rect 11974 17212 11980 17264
rect 12032 17252 12038 17264
rect 12989 17255 13047 17261
rect 12989 17252 13001 17255
rect 12032 17224 13001 17252
rect 12032 17212 12038 17224
rect 12989 17221 13001 17224
rect 13035 17221 13047 17255
rect 12989 17215 13047 17221
rect 13081 17255 13139 17261
rect 13081 17221 13093 17255
rect 13127 17252 13139 17255
rect 13630 17252 13636 17264
rect 13127 17224 13636 17252
rect 13127 17221 13139 17224
rect 13081 17215 13139 17221
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 14274 17212 14280 17264
rect 14332 17212 14338 17264
rect 16390 17212 16396 17264
rect 16448 17252 16454 17264
rect 17957 17255 18015 17261
rect 17957 17252 17969 17255
rect 16448 17224 17969 17252
rect 16448 17212 16454 17224
rect 17957 17221 17969 17224
rect 18003 17252 18015 17255
rect 18874 17252 18880 17264
rect 18003 17224 18880 17252
rect 18003 17221 18015 17224
rect 17957 17215 18015 17221
rect 18874 17212 18880 17224
rect 18932 17212 18938 17264
rect 18966 17212 18972 17264
rect 19024 17252 19030 17264
rect 19306 17252 19334 17292
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 22649 17323 22707 17329
rect 22649 17289 22661 17323
rect 22695 17320 22707 17323
rect 23474 17320 23480 17332
rect 22695 17292 23480 17320
rect 22695 17289 22707 17292
rect 22649 17283 22707 17289
rect 23474 17280 23480 17292
rect 23532 17280 23538 17332
rect 24854 17280 24860 17332
rect 24912 17280 24918 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 27341 17323 27399 17329
rect 27341 17320 27353 17323
rect 25363 17292 27353 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 27341 17289 27353 17292
rect 27387 17289 27399 17323
rect 27341 17283 27399 17289
rect 27798 17280 27804 17332
rect 27856 17320 27862 17332
rect 28997 17323 29055 17329
rect 28997 17320 29009 17323
rect 27856 17292 29009 17320
rect 27856 17280 27862 17292
rect 28997 17289 29009 17292
rect 29043 17289 29055 17323
rect 30650 17320 30656 17332
rect 28997 17283 29055 17289
rect 30116 17292 30656 17320
rect 20530 17252 20536 17264
rect 19024 17224 19334 17252
rect 20194 17224 20536 17252
rect 19024 17212 19030 17224
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 20625 17255 20683 17261
rect 20625 17221 20637 17255
rect 20671 17252 20683 17255
rect 21266 17252 21272 17264
rect 20671 17224 21272 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 21266 17212 21272 17224
rect 21324 17212 21330 17264
rect 21542 17212 21548 17264
rect 21600 17252 21606 17264
rect 21726 17252 21732 17264
rect 21600 17224 21732 17252
rect 21600 17212 21606 17224
rect 21726 17212 21732 17224
rect 21784 17252 21790 17264
rect 21913 17255 21971 17261
rect 21913 17252 21925 17255
rect 21784 17224 21925 17252
rect 21784 17212 21790 17224
rect 21913 17221 21925 17224
rect 21959 17221 21971 17255
rect 22094 17252 22100 17264
rect 21913 17215 21971 17221
rect 22066 17212 22100 17252
rect 22152 17252 22158 17264
rect 22738 17252 22744 17264
rect 22152 17224 22744 17252
rect 22152 17212 22158 17224
rect 22738 17212 22744 17224
rect 22796 17212 22802 17264
rect 24118 17212 24124 17264
rect 24176 17252 24182 17264
rect 24176 17224 24440 17252
rect 24176 17212 24182 17224
rect 14182 17184 14188 17196
rect 11900 17156 14188 17184
rect 10781 17147 10839 17153
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 934 17076 940 17128
rect 992 17116 998 17128
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 992 17088 1777 17116
rect 992 17076 998 17088
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 9490 17076 9496 17128
rect 9548 17076 9554 17128
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 5442 17008 5448 17060
rect 5500 17048 5506 17060
rect 9769 17051 9827 17057
rect 5500 17020 9628 17048
rect 5500 17008 5506 17020
rect 9600 16980 9628 17020
rect 9769 17017 9781 17051
rect 9815 17048 9827 17051
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 9815 17020 10057 17048
rect 9815 17017 9827 17020
rect 9769 17011 9827 17017
rect 10045 17017 10057 17020
rect 10091 17048 10103 17051
rect 10520 17048 10548 17079
rect 10594 17076 10600 17128
rect 10652 17116 10658 17128
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 10652 17088 10701 17116
rect 10652 17076 10658 17088
rect 10689 17085 10701 17088
rect 10735 17085 10747 17119
rect 12342 17116 12348 17128
rect 10689 17079 10747 17085
rect 11072 17088 12348 17116
rect 11072 17048 11100 17088
rect 12342 17076 12348 17088
rect 12400 17116 12406 17128
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 12400 17088 12817 17116
rect 12400 17076 12406 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 14292 17116 14320 17212
rect 15102 17144 15108 17196
rect 15160 17144 15166 17196
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15436 17156 15945 17184
rect 15436 17144 15442 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 12805 17079 12863 17085
rect 13832 17088 14320 17116
rect 16025 17119 16083 17125
rect 10091 17020 11100 17048
rect 11149 17051 11207 17057
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 11790 17048 11796 17060
rect 11195 17020 11796 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 11790 17008 11796 17020
rect 11848 17008 11854 17060
rect 12437 17051 12495 17057
rect 12437 17017 12449 17051
rect 12483 17048 12495 17051
rect 13832 17048 13860 17088
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 12483 17020 13860 17048
rect 12483 17017 12495 17020
rect 12437 17011 12495 17017
rect 13906 17008 13912 17060
rect 13964 17048 13970 17060
rect 14921 17051 14979 17057
rect 14921 17048 14933 17051
rect 13964 17020 14933 17048
rect 13964 17008 13970 17020
rect 14921 17017 14933 17020
rect 14967 17017 14979 17051
rect 14921 17011 14979 17017
rect 15562 17008 15568 17060
rect 15620 17008 15626 17060
rect 16040 17048 16068 17079
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 17050 17116 17078 17147
rect 18598 17144 18604 17196
rect 18656 17184 18662 17196
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 18656 17156 18705 17184
rect 18656 17144 18662 17156
rect 18693 17153 18705 17156
rect 18739 17184 18751 17187
rect 19058 17184 19064 17196
rect 18739 17156 19064 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 22066 17184 22094 17212
rect 24412 17193 24440 17224
rect 25958 17212 25964 17264
rect 26016 17212 26022 17264
rect 26878 17212 26884 17264
rect 26936 17252 26942 17264
rect 28905 17255 28963 17261
rect 26936 17224 28120 17252
rect 26936 17212 26942 17224
rect 20947 17156 22094 17184
rect 24397 17187 24455 17193
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 19886 17116 19892 17128
rect 17050 17088 19892 17116
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 16482 17048 16488 17060
rect 16040 17020 16488 17048
rect 16482 17008 16488 17020
rect 16540 17048 16546 17060
rect 21269 17051 21327 17057
rect 16540 17020 17080 17048
rect 16540 17008 16546 17020
rect 12250 16980 12256 16992
rect 9600 16952 12256 16980
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 13354 16940 13360 16992
rect 13412 16980 13418 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 13412 16952 13461 16980
rect 13412 16940 13418 16952
rect 13449 16949 13461 16952
rect 13495 16949 13507 16983
rect 13449 16943 13507 16949
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 15838 16980 15844 16992
rect 13780 16952 15844 16980
rect 13780 16940 13786 16952
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 15988 16952 16957 16980
rect 15988 16940 15994 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 17052 16980 17080 17020
rect 21269 17017 21281 17051
rect 21315 17048 21327 17051
rect 21634 17048 21640 17060
rect 21315 17020 21640 17048
rect 21315 17017 21327 17020
rect 21269 17011 21327 17017
rect 21634 17008 21640 17020
rect 21692 17048 21698 17060
rect 22278 17048 22284 17060
rect 21692 17020 22284 17048
rect 21692 17008 21698 17020
rect 22278 17008 22284 17020
rect 22336 17048 22342 17060
rect 23032 17048 23060 17170
rect 24397 17153 24409 17187
rect 24443 17153 24455 17187
rect 24397 17147 24455 17153
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17184 25283 17187
rect 25590 17184 25596 17196
rect 25271 17156 25596 17184
rect 25271 17153 25283 17156
rect 25225 17147 25283 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 27614 17144 27620 17196
rect 27672 17184 27678 17196
rect 27709 17187 27767 17193
rect 27709 17184 27721 17187
rect 27672 17156 27721 17184
rect 27672 17144 27678 17156
rect 27709 17153 27721 17156
rect 27755 17153 27767 17187
rect 27982 17184 27988 17196
rect 27709 17147 27767 17153
rect 27816 17156 27988 17184
rect 24121 17119 24179 17125
rect 24121 17085 24133 17119
rect 24167 17116 24179 17119
rect 24486 17116 24492 17128
rect 24167 17088 24492 17116
rect 24167 17085 24179 17088
rect 24121 17079 24179 17085
rect 24486 17076 24492 17088
rect 24544 17076 24550 17128
rect 25498 17076 25504 17128
rect 25556 17076 25562 17128
rect 26970 17076 26976 17128
rect 27028 17116 27034 17128
rect 27816 17125 27844 17156
rect 27982 17144 27988 17156
rect 28040 17144 28046 17196
rect 28092 17184 28120 17224
rect 28905 17221 28917 17255
rect 28951 17252 28963 17255
rect 29546 17252 29552 17264
rect 28951 17224 29552 17252
rect 28951 17221 28963 17224
rect 28905 17215 28963 17221
rect 29546 17212 29552 17224
rect 29604 17212 29610 17264
rect 30116 17184 30144 17292
rect 30650 17280 30656 17292
rect 30708 17280 30714 17332
rect 31386 17280 31392 17332
rect 31444 17320 31450 17332
rect 33594 17320 33600 17332
rect 31444 17292 33600 17320
rect 31444 17280 31450 17292
rect 30193 17255 30251 17261
rect 30193 17221 30205 17255
rect 30239 17252 30251 17255
rect 32030 17252 32036 17264
rect 30239 17224 32036 17252
rect 30239 17221 30251 17224
rect 30193 17215 30251 17221
rect 32030 17212 32036 17224
rect 32088 17212 32094 17264
rect 28092 17156 28948 17184
rect 27801 17119 27859 17125
rect 27801 17116 27813 17119
rect 27028 17088 27813 17116
rect 27028 17076 27034 17088
rect 27801 17085 27813 17088
rect 27847 17085 27859 17119
rect 27801 17079 27859 17085
rect 27890 17076 27896 17128
rect 27948 17076 27954 17128
rect 28721 17119 28779 17125
rect 28721 17085 28733 17119
rect 28767 17085 28779 17119
rect 28721 17079 28779 17085
rect 22336 17020 23060 17048
rect 22336 17008 22342 17020
rect 27246 17008 27252 17060
rect 27304 17048 27310 17060
rect 28736 17048 28764 17079
rect 27304 17020 28764 17048
rect 27304 17008 27310 17020
rect 22370 16980 22376 16992
rect 17052 16952 22376 16980
rect 16945 16943 17003 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 28920 16980 28948 17156
rect 30024 17156 30144 17184
rect 29730 17076 29736 17128
rect 29788 17116 29794 17128
rect 30024 17125 30052 17156
rect 30558 17144 30564 17196
rect 30616 17184 30622 17196
rect 31297 17187 31355 17193
rect 31297 17184 31309 17187
rect 30616 17156 31309 17184
rect 30616 17144 30622 17156
rect 31297 17153 31309 17156
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 31389 17187 31447 17193
rect 31389 17153 31401 17187
rect 31435 17153 31447 17187
rect 31389 17147 31447 17153
rect 30009 17119 30067 17125
rect 30009 17116 30021 17119
rect 29788 17088 30021 17116
rect 29788 17076 29794 17088
rect 30009 17085 30021 17088
rect 30055 17085 30067 17119
rect 30009 17079 30067 17085
rect 30098 17076 30104 17128
rect 30156 17076 30162 17128
rect 30374 17076 30380 17128
rect 30432 17116 30438 17128
rect 30432 17088 30604 17116
rect 30432 17076 30438 17088
rect 29365 17051 29423 17057
rect 29365 17017 29377 17051
rect 29411 17048 29423 17051
rect 30282 17048 30288 17060
rect 29411 17020 30288 17048
rect 29411 17017 29423 17020
rect 29365 17011 29423 17017
rect 30282 17008 30288 17020
rect 30340 17008 30346 17060
rect 30576 17057 30604 17088
rect 30742 17076 30748 17128
rect 30800 17116 30806 17128
rect 31113 17119 31171 17125
rect 31113 17116 31125 17119
rect 30800 17088 31125 17116
rect 30800 17076 30806 17088
rect 31113 17085 31125 17088
rect 31159 17085 31171 17119
rect 31113 17079 31171 17085
rect 30561 17051 30619 17057
rect 30561 17017 30573 17051
rect 30607 17017 30619 17051
rect 31404 17048 31432 17147
rect 32214 17144 32220 17196
rect 32272 17184 32278 17196
rect 32324 17193 32352 17292
rect 33594 17280 33600 17292
rect 33652 17280 33658 17332
rect 35066 17280 35072 17332
rect 35124 17320 35130 17332
rect 37829 17323 37887 17329
rect 37829 17320 37841 17323
rect 35124 17292 37841 17320
rect 35124 17280 35130 17292
rect 37829 17289 37841 17292
rect 37875 17289 37887 17323
rect 37829 17283 37887 17289
rect 38470 17280 38476 17332
rect 38528 17320 38534 17332
rect 38654 17320 38660 17332
rect 38528 17292 38660 17320
rect 38528 17280 38534 17292
rect 38654 17280 38660 17292
rect 38712 17280 38718 17332
rect 40034 17280 40040 17332
rect 40092 17320 40098 17332
rect 40957 17323 41015 17329
rect 40957 17320 40969 17323
rect 40092 17292 40969 17320
rect 40092 17280 40098 17292
rect 40957 17289 40969 17292
rect 41003 17320 41015 17323
rect 41046 17320 41052 17332
rect 41003 17292 41052 17320
rect 41003 17289 41015 17292
rect 40957 17283 41015 17289
rect 41046 17280 41052 17292
rect 41104 17280 41110 17332
rect 47026 17280 47032 17332
rect 47084 17280 47090 17332
rect 34422 17252 34428 17264
rect 33810 17224 34428 17252
rect 34422 17212 34428 17224
rect 34480 17212 34486 17264
rect 35434 17212 35440 17264
rect 35492 17252 35498 17264
rect 35529 17255 35587 17261
rect 35529 17252 35541 17255
rect 35492 17224 35541 17252
rect 35492 17212 35498 17224
rect 35529 17221 35541 17224
rect 35575 17252 35587 17255
rect 37001 17255 37059 17261
rect 37001 17252 37013 17255
rect 35575 17224 37013 17252
rect 35575 17221 35587 17224
rect 35529 17215 35587 17221
rect 37001 17221 37013 17224
rect 37047 17221 37059 17255
rect 38672 17252 38700 17280
rect 39114 17252 39120 17264
rect 38672 17224 39120 17252
rect 37001 17215 37059 17221
rect 39114 17212 39120 17224
rect 39172 17252 39178 17264
rect 39172 17224 39238 17252
rect 39172 17212 39178 17224
rect 40126 17212 40132 17264
rect 40184 17252 40190 17264
rect 40405 17255 40463 17261
rect 40405 17252 40417 17255
rect 40184 17224 40417 17252
rect 40184 17212 40190 17224
rect 40405 17221 40417 17224
rect 40451 17221 40463 17255
rect 40405 17215 40463 17221
rect 47670 17212 47676 17264
rect 47728 17252 47734 17264
rect 48222 17252 48228 17264
rect 47728 17224 48228 17252
rect 47728 17212 47734 17224
rect 48222 17212 48228 17224
rect 48280 17252 48286 17264
rect 48280 17224 49372 17252
rect 48280 17212 48286 17224
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 32272 17156 32321 17184
rect 32272 17144 32278 17156
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 35158 17144 35164 17196
rect 35216 17184 35222 17196
rect 36265 17187 36323 17193
rect 36265 17184 36277 17187
rect 35216 17156 36277 17184
rect 35216 17144 35222 17156
rect 36265 17153 36277 17156
rect 36311 17153 36323 17187
rect 36265 17147 36323 17153
rect 36354 17144 36360 17196
rect 36412 17144 36418 17196
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17184 37979 17187
rect 38930 17184 38936 17196
rect 37967 17156 38936 17184
rect 37967 17153 37979 17156
rect 37921 17147 37979 17153
rect 38930 17144 38936 17156
rect 38988 17144 38994 17196
rect 49344 17193 49372 17224
rect 47213 17187 47271 17193
rect 47213 17153 47225 17187
rect 47259 17184 47271 17187
rect 48133 17187 48191 17193
rect 47259 17156 47716 17184
rect 47259 17153 47271 17156
rect 47213 17147 47271 17153
rect 32582 17076 32588 17128
rect 32640 17076 32646 17128
rect 32674 17076 32680 17128
rect 32732 17116 32738 17128
rect 34057 17119 34115 17125
rect 34057 17116 34069 17119
rect 32732 17088 34069 17116
rect 32732 17076 32738 17088
rect 34057 17085 34069 17088
rect 34103 17085 34115 17119
rect 34057 17079 34115 17085
rect 34790 17076 34796 17128
rect 34848 17076 34854 17128
rect 36081 17119 36139 17125
rect 36081 17085 36093 17119
rect 36127 17116 36139 17119
rect 36538 17116 36544 17128
rect 36127 17088 36544 17116
rect 36127 17085 36139 17088
rect 36081 17079 36139 17085
rect 36538 17076 36544 17088
rect 36596 17076 36602 17128
rect 37826 17076 37832 17128
rect 37884 17116 37890 17128
rect 38013 17119 38071 17125
rect 38013 17116 38025 17119
rect 37884 17088 38025 17116
rect 37884 17076 37890 17088
rect 38013 17085 38025 17088
rect 38059 17085 38071 17119
rect 38013 17079 38071 17085
rect 38626 17088 40632 17116
rect 31570 17048 31576 17060
rect 31404 17020 31576 17048
rect 30561 17011 30619 17017
rect 31570 17008 31576 17020
rect 31628 17008 31634 17060
rect 33870 17008 33876 17060
rect 33928 17048 33934 17060
rect 38626 17048 38654 17088
rect 33928 17020 38654 17048
rect 40604 17048 40632 17088
rect 40678 17076 40684 17128
rect 40736 17076 40742 17128
rect 40604 17020 41414 17048
rect 33928 17008 33934 17020
rect 30190 16980 30196 16992
rect 28920 16952 30196 16980
rect 30190 16940 30196 16952
rect 30248 16940 30254 16992
rect 31754 16940 31760 16992
rect 31812 16940 31818 16992
rect 35342 16940 35348 16992
rect 35400 16980 35406 16992
rect 36630 16980 36636 16992
rect 35400 16952 36636 16980
rect 35400 16940 35406 16952
rect 36630 16940 36636 16952
rect 36688 16940 36694 16992
rect 36725 16983 36783 16989
rect 36725 16949 36737 16983
rect 36771 16980 36783 16983
rect 37274 16980 37280 16992
rect 36771 16952 37280 16980
rect 36771 16949 36783 16952
rect 36725 16943 36783 16949
rect 37274 16940 37280 16952
rect 37332 16940 37338 16992
rect 37458 16940 37464 16992
rect 37516 16940 37522 16992
rect 38838 16940 38844 16992
rect 38896 16980 38902 16992
rect 38933 16983 38991 16989
rect 38933 16980 38945 16983
rect 38896 16952 38945 16980
rect 38896 16940 38902 16952
rect 38933 16949 38945 16952
rect 38979 16980 38991 16983
rect 40770 16980 40776 16992
rect 38979 16952 40776 16980
rect 38979 16949 38991 16952
rect 38933 16943 38991 16949
rect 40770 16940 40776 16952
rect 40828 16940 40834 16992
rect 41386 16980 41414 17020
rect 41690 16980 41696 16992
rect 41386 16952 41696 16980
rect 41690 16940 41696 16952
rect 41748 16940 41754 16992
rect 47688 16989 47716 17156
rect 48133 17153 48145 17187
rect 48179 17184 48191 17187
rect 48685 17187 48743 17193
rect 48685 17184 48697 17187
rect 48179 17156 48697 17184
rect 48179 17153 48191 17156
rect 48133 17147 48191 17153
rect 48685 17153 48697 17156
rect 48731 17153 48743 17187
rect 48685 17147 48743 17153
rect 49329 17187 49387 17193
rect 49329 17153 49341 17187
rect 49375 17153 49387 17187
rect 49329 17147 49387 17153
rect 47946 17076 47952 17128
rect 48004 17076 48010 17128
rect 47673 16983 47731 16989
rect 47673 16949 47685 16983
rect 47719 16980 47731 16983
rect 48314 16980 48320 16992
rect 47719 16952 48320 16980
rect 47719 16949 47731 16952
rect 47673 16943 47731 16949
rect 48314 16940 48320 16952
rect 48372 16940 48378 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 10410 16736 10416 16788
rect 10468 16736 10474 16788
rect 11974 16776 11980 16788
rect 10520 16748 11980 16776
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 10520 16708 10548 16748
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 13722 16776 13728 16788
rect 12308 16748 13728 16776
rect 12308 16736 12314 16748
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 13906 16736 13912 16788
rect 13964 16776 13970 16788
rect 14918 16776 14924 16788
rect 13964 16748 14924 16776
rect 13964 16736 13970 16748
rect 14918 16736 14924 16748
rect 14976 16736 14982 16788
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16264 16748 16681 16776
rect 16264 16736 16270 16748
rect 16669 16745 16681 16748
rect 16715 16776 16727 16779
rect 18966 16776 18972 16788
rect 16715 16748 18972 16776
rect 16715 16745 16727 16748
rect 16669 16739 16727 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19058 16736 19064 16788
rect 19116 16776 19122 16788
rect 23382 16776 23388 16788
rect 19116 16748 23388 16776
rect 19116 16736 19122 16748
rect 23382 16736 23388 16748
rect 23440 16776 23446 16788
rect 24673 16779 24731 16785
rect 24673 16776 24685 16779
rect 23440 16748 24685 16776
rect 23440 16736 23446 16748
rect 24673 16745 24685 16748
rect 24719 16776 24731 16779
rect 26326 16776 26332 16788
rect 24719 16748 26332 16776
rect 24719 16745 24731 16748
rect 24673 16739 24731 16745
rect 26326 16736 26332 16748
rect 26384 16776 26390 16788
rect 27614 16776 27620 16788
rect 26384 16748 27620 16776
rect 26384 16736 26390 16748
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 28261 16779 28319 16785
rect 28261 16745 28273 16779
rect 28307 16776 28319 16779
rect 28534 16776 28540 16788
rect 28307 16748 28540 16776
rect 28307 16745 28319 16748
rect 28261 16739 28319 16745
rect 28534 16736 28540 16748
rect 28592 16776 28598 16788
rect 28718 16776 28724 16788
rect 28592 16748 28724 16776
rect 28592 16736 28598 16748
rect 28718 16736 28724 16748
rect 28776 16736 28782 16788
rect 29362 16736 29368 16788
rect 29420 16776 29426 16788
rect 30098 16776 30104 16788
rect 29420 16748 30104 16776
rect 29420 16736 29426 16748
rect 30098 16736 30104 16748
rect 30156 16736 30162 16788
rect 33870 16776 33876 16788
rect 30300 16748 33876 16776
rect 9916 16680 10548 16708
rect 9916 16668 9922 16680
rect 10594 16668 10600 16720
rect 10652 16708 10658 16720
rect 14734 16708 14740 16720
rect 10652 16680 13124 16708
rect 10652 16668 10658 16680
rect 4430 16600 4436 16652
rect 4488 16640 4494 16652
rect 7929 16643 7987 16649
rect 4488 16612 7512 16640
rect 4488 16600 4494 16612
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3326 16572 3332 16584
rect 3007 16544 3332 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 1026 16464 1032 16516
rect 1084 16504 1090 16516
rect 1765 16507 1823 16513
rect 1765 16504 1777 16507
rect 1084 16476 1777 16504
rect 1084 16464 1090 16476
rect 1765 16473 1777 16476
rect 1811 16473 1823 16507
rect 7484 16504 7512 16612
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 9030 16640 9036 16652
rect 7975 16612 9036 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9490 16600 9496 16652
rect 9548 16640 9554 16652
rect 10502 16640 10508 16652
rect 9548 16612 10508 16640
rect 9548 16600 9554 16612
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 11146 16600 11152 16652
rect 11204 16600 11210 16652
rect 11790 16600 11796 16652
rect 11848 16640 11854 16652
rect 12618 16640 12624 16652
rect 11848 16612 12624 16640
rect 11848 16600 11854 16612
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 7558 16532 7564 16584
rect 7616 16572 7622 16584
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 7616 16544 8125 16572
rect 7616 16532 7622 16544
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12158 16572 12164 16584
rect 12032 16544 12164 16572
rect 12032 16532 12038 16544
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12308 16544 12357 16572
rect 12308 16532 12314 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 13096 16572 13124 16680
rect 13188 16680 14740 16708
rect 13188 16649 13216 16680
rect 14734 16668 14740 16680
rect 14792 16708 14798 16720
rect 14792 16680 16252 16708
rect 14792 16668 14798 16680
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13906 16640 13912 16652
rect 13311 16612 13912 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13280 16572 13308 16603
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14182 16600 14188 16652
rect 14240 16600 14246 16652
rect 14645 16643 14703 16649
rect 14645 16609 14657 16643
rect 14691 16640 14703 16643
rect 14691 16612 15792 16640
rect 14691 16609 14703 16612
rect 14645 16603 14703 16609
rect 15764 16584 15792 16612
rect 15838 16600 15844 16652
rect 15896 16640 15902 16652
rect 16224 16649 16252 16680
rect 16942 16668 16948 16720
rect 17000 16708 17006 16720
rect 17494 16708 17500 16720
rect 17000 16680 17500 16708
rect 17000 16668 17006 16680
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 20990 16668 20996 16720
rect 21048 16708 21054 16720
rect 21266 16708 21272 16720
rect 21048 16680 21272 16708
rect 21048 16668 21054 16680
rect 21266 16668 21272 16680
rect 21324 16668 21330 16720
rect 26050 16708 26056 16720
rect 23768 16680 26056 16708
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15896 16612 16129 16640
rect 15896 16600 15902 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16609 16267 16643
rect 18230 16640 18236 16652
rect 16209 16603 16267 16609
rect 17420 16612 18236 16640
rect 13096 16544 13308 16572
rect 13357 16575 13415 16581
rect 12345 16535 12403 16541
rect 13357 16541 13369 16575
rect 13403 16572 13415 16575
rect 13814 16572 13820 16584
rect 13403 16544 13820 16572
rect 13403 16541 13415 16544
rect 13357 16535 13415 16541
rect 13814 16532 13820 16544
rect 13872 16572 13878 16584
rect 14829 16575 14887 16581
rect 14829 16572 14841 16575
rect 13872 16544 14841 16572
rect 13872 16532 13878 16544
rect 14829 16541 14841 16544
rect 14875 16541 14887 16575
rect 14829 16535 14887 16541
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 17420 16572 17448 16612
rect 18230 16600 18236 16612
rect 18288 16600 18294 16652
rect 18598 16600 18604 16652
rect 18656 16600 18662 16652
rect 18874 16600 18880 16652
rect 18932 16600 18938 16652
rect 22462 16600 22468 16652
rect 22520 16600 22526 16652
rect 22738 16600 22744 16652
rect 22796 16600 22802 16652
rect 23768 16649 23796 16680
rect 26050 16668 26056 16680
rect 26108 16668 26114 16720
rect 27982 16668 27988 16720
rect 28040 16708 28046 16720
rect 28813 16711 28871 16717
rect 28813 16708 28825 16711
rect 28040 16680 28825 16708
rect 28040 16668 28046 16680
rect 28813 16677 28825 16680
rect 28859 16677 28871 16711
rect 28813 16671 28871 16677
rect 29181 16711 29239 16717
rect 29181 16677 29193 16711
rect 29227 16708 29239 16711
rect 29227 16680 29960 16708
rect 29227 16677 29239 16680
rect 29181 16671 29239 16677
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23937 16643 23995 16649
rect 23937 16609 23949 16643
rect 23983 16640 23995 16643
rect 25593 16643 25651 16649
rect 25593 16640 25605 16643
rect 23983 16612 25605 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 25593 16609 25605 16612
rect 25639 16640 25651 16643
rect 25866 16640 25872 16652
rect 25639 16612 25872 16640
rect 25639 16609 25651 16612
rect 25593 16603 25651 16609
rect 25866 16600 25872 16612
rect 25924 16600 25930 16652
rect 27062 16600 27068 16652
rect 27120 16600 27126 16652
rect 27430 16600 27436 16652
rect 27488 16640 27494 16652
rect 27617 16643 27675 16649
rect 27617 16640 27629 16643
rect 27488 16612 27629 16640
rect 27488 16600 27494 16612
rect 27617 16609 27629 16612
rect 27663 16609 27675 16643
rect 27617 16603 27675 16609
rect 29454 16600 29460 16652
rect 29512 16640 29518 16652
rect 29825 16643 29883 16649
rect 29825 16640 29837 16643
rect 29512 16612 29837 16640
rect 29512 16600 29518 16612
rect 29825 16609 29837 16612
rect 29871 16609 29883 16643
rect 29932 16640 29960 16680
rect 30006 16640 30012 16652
rect 29932 16612 30012 16640
rect 29825 16603 29883 16609
rect 30006 16600 30012 16612
rect 30064 16600 30070 16652
rect 15804 16544 17448 16572
rect 15804 16532 15810 16544
rect 17494 16532 17500 16584
rect 17552 16532 17558 16584
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 8021 16507 8079 16513
rect 8021 16504 8033 16507
rect 7484 16476 8033 16504
rect 1765 16467 1823 16473
rect 8021 16473 8033 16476
rect 8067 16473 8079 16507
rect 9674 16504 9680 16516
rect 8021 16467 8079 16473
rect 8496 16476 9680 16504
rect 8496 16445 8524 16476
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 10045 16507 10103 16513
rect 10045 16473 10057 16507
rect 10091 16504 10103 16507
rect 10502 16504 10508 16516
rect 10091 16476 10508 16504
rect 10091 16473 10103 16476
rect 10045 16467 10103 16473
rect 10502 16464 10508 16476
rect 10560 16464 10566 16516
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 12802 16504 12808 16516
rect 11471 16476 12808 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 14642 16464 14648 16516
rect 14700 16504 14706 16516
rect 20272 16504 20300 16535
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20772 16544 21390 16572
rect 20772 16532 20778 16544
rect 24578 16532 24584 16584
rect 24636 16572 24642 16584
rect 27341 16575 27399 16581
rect 24636 16544 25912 16572
rect 24636 16532 24642 16544
rect 14700 16476 17356 16504
rect 14700 16464 14706 16476
rect 8481 16439 8539 16445
rect 8481 16405 8493 16439
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 9030 16396 9036 16448
rect 9088 16396 9094 16448
rect 11330 16396 11336 16448
rect 11388 16396 11394 16448
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16436 11851 16439
rect 12158 16436 12164 16448
rect 11839 16408 12164 16436
rect 11839 16405 11851 16408
rect 11793 16399 11851 16405
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 12529 16439 12587 16445
rect 12529 16405 12541 16439
rect 12575 16436 12587 16439
rect 12710 16436 12716 16448
rect 12575 16408 12716 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 13504 16408 13737 16436
rect 13504 16396 13510 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 14737 16439 14795 16445
rect 14737 16405 14749 16439
rect 14783 16436 14795 16439
rect 14918 16436 14924 16448
rect 14783 16408 14924 16436
rect 14783 16405 14795 16408
rect 14737 16399 14795 16405
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16436 15255 16439
rect 15470 16436 15476 16448
rect 15243 16408 15476 16436
rect 15243 16405 15255 16408
rect 15197 16399 15255 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15654 16396 15660 16448
rect 15712 16396 15718 16448
rect 16025 16439 16083 16445
rect 16025 16405 16037 16439
rect 16071 16436 16083 16439
rect 16206 16436 16212 16448
rect 16071 16408 16212 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 17126 16396 17132 16448
rect 17184 16396 17190 16448
rect 17328 16436 17356 16476
rect 18248 16476 20116 16504
rect 20272 16476 21220 16504
rect 25884 16490 25912 16544
rect 27341 16541 27353 16575
rect 27387 16572 27399 16575
rect 28902 16572 28908 16584
rect 27387 16544 28908 16572
rect 27387 16541 27399 16544
rect 27341 16535 27399 16541
rect 28902 16532 28908 16544
rect 28960 16532 28966 16584
rect 28994 16532 29000 16584
rect 29052 16572 29058 16584
rect 30101 16575 30159 16581
rect 30101 16572 30113 16575
rect 29052 16544 30113 16572
rect 29052 16532 29058 16544
rect 30101 16541 30113 16544
rect 30147 16541 30159 16575
rect 30101 16535 30159 16541
rect 18248 16436 18276 16476
rect 17328 16408 18276 16436
rect 18322 16396 18328 16448
rect 18380 16436 18386 16448
rect 18966 16436 18972 16448
rect 18380 16408 18972 16436
rect 18380 16396 18386 16408
rect 18966 16396 18972 16408
rect 19024 16396 19030 16448
rect 19426 16396 19432 16448
rect 19484 16396 19490 16448
rect 20088 16445 20116 16476
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16405 20131 16439
rect 20073 16399 20131 16405
rect 20625 16439 20683 16445
rect 20625 16405 20637 16439
rect 20671 16436 20683 16439
rect 20714 16436 20720 16448
rect 20671 16408 20720 16436
rect 20671 16405 20683 16408
rect 20625 16399 20683 16405
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 21192 16436 21220 16476
rect 28442 16464 28448 16516
rect 28500 16504 28506 16516
rect 30300 16504 30328 16748
rect 33870 16736 33876 16748
rect 33928 16736 33934 16788
rect 34422 16736 34428 16788
rect 34480 16776 34486 16788
rect 34517 16779 34575 16785
rect 34517 16776 34529 16779
rect 34480 16748 34529 16776
rect 34480 16736 34486 16748
rect 34517 16745 34529 16748
rect 34563 16776 34575 16779
rect 36170 16776 36176 16788
rect 34563 16748 36176 16776
rect 34563 16745 34575 16748
rect 34517 16739 34575 16745
rect 36170 16736 36176 16748
rect 36228 16736 36234 16788
rect 36265 16779 36323 16785
rect 36265 16745 36277 16779
rect 36311 16776 36323 16779
rect 36354 16776 36360 16788
rect 36311 16748 36360 16776
rect 36311 16745 36323 16748
rect 36265 16739 36323 16745
rect 36354 16736 36360 16748
rect 36412 16736 36418 16788
rect 36630 16736 36636 16788
rect 36688 16776 36694 16788
rect 36688 16748 38240 16776
rect 36688 16736 36694 16748
rect 30558 16668 30564 16720
rect 30616 16708 30622 16720
rect 37550 16708 37556 16720
rect 30616 16680 32352 16708
rect 30616 16668 30622 16680
rect 31110 16600 31116 16652
rect 31168 16600 31174 16652
rect 31205 16643 31263 16649
rect 31205 16609 31217 16643
rect 31251 16640 31263 16643
rect 31251 16612 31754 16640
rect 31251 16609 31263 16612
rect 31205 16603 31263 16609
rect 31018 16572 31024 16584
rect 28500 16476 30328 16504
rect 30392 16544 31024 16572
rect 28500 16464 28506 16476
rect 22830 16436 22836 16448
rect 21192 16408 22836 16436
rect 22830 16396 22836 16408
rect 22888 16396 22894 16448
rect 23290 16396 23296 16448
rect 23348 16396 23354 16448
rect 23658 16396 23664 16448
rect 23716 16396 23722 16448
rect 27522 16396 27528 16448
rect 27580 16436 27586 16448
rect 27985 16439 28043 16445
rect 27985 16436 27997 16439
rect 27580 16408 27997 16436
rect 27580 16396 27586 16408
rect 27985 16405 27997 16408
rect 28031 16405 28043 16439
rect 27985 16399 28043 16405
rect 28166 16396 28172 16448
rect 28224 16436 28230 16448
rect 28537 16439 28595 16445
rect 28537 16436 28549 16439
rect 28224 16408 28549 16436
rect 28224 16396 28230 16408
rect 28537 16405 28549 16408
rect 28583 16405 28595 16439
rect 28537 16399 28595 16405
rect 29362 16396 29368 16448
rect 29420 16436 29426 16448
rect 30392 16436 30420 16544
rect 31018 16532 31024 16544
rect 31076 16532 31082 16584
rect 31726 16572 31754 16612
rect 32214 16600 32220 16652
rect 32272 16600 32278 16652
rect 32324 16640 32352 16680
rect 35084 16680 37556 16708
rect 32490 16640 32496 16652
rect 32324 16612 32496 16640
rect 32490 16600 32496 16612
rect 32548 16600 32554 16652
rect 35084 16649 35112 16680
rect 37550 16668 37556 16680
rect 37608 16668 37614 16720
rect 35069 16643 35127 16649
rect 35069 16609 35081 16643
rect 35115 16609 35127 16643
rect 35069 16603 35127 16609
rect 36909 16643 36967 16649
rect 36909 16609 36921 16643
rect 36955 16640 36967 16643
rect 37090 16640 37096 16652
rect 36955 16612 37096 16640
rect 36955 16609 36967 16612
rect 36909 16603 36967 16609
rect 37090 16600 37096 16612
rect 37148 16600 37154 16652
rect 38212 16640 38240 16748
rect 40218 16736 40224 16788
rect 40276 16736 40282 16788
rect 41046 16736 41052 16788
rect 41104 16736 41110 16788
rect 41230 16736 41236 16788
rect 41288 16736 41294 16788
rect 40236 16708 40264 16736
rect 41509 16711 41567 16717
rect 41509 16708 41521 16711
rect 40236 16680 41521 16708
rect 41509 16677 41521 16680
rect 41555 16708 41567 16711
rect 48774 16708 48780 16720
rect 41555 16680 48780 16708
rect 41555 16677 41567 16680
rect 41509 16671 41567 16677
rect 48774 16668 48780 16680
rect 48832 16668 48838 16720
rect 38838 16640 38844 16652
rect 38212 16612 38844 16640
rect 38838 16600 38844 16612
rect 38896 16640 38902 16652
rect 39209 16643 39267 16649
rect 39209 16640 39221 16643
rect 38896 16612 39221 16640
rect 38896 16600 38902 16612
rect 39209 16609 39221 16612
rect 39255 16609 39267 16643
rect 39209 16603 39267 16609
rect 40221 16643 40279 16649
rect 40221 16609 40233 16643
rect 40267 16640 40279 16643
rect 40310 16640 40316 16652
rect 40267 16612 40316 16640
rect 40267 16609 40279 16612
rect 40221 16603 40279 16609
rect 40310 16600 40316 16612
rect 40368 16600 40374 16652
rect 41046 16600 41052 16652
rect 41104 16640 41110 16652
rect 47673 16643 47731 16649
rect 41104 16612 41414 16640
rect 41104 16600 41110 16612
rect 31938 16572 31944 16584
rect 31726 16544 31944 16572
rect 31938 16532 31944 16544
rect 31996 16532 32002 16584
rect 34422 16572 34428 16584
rect 33626 16544 34428 16572
rect 34422 16532 34428 16544
rect 34480 16532 34486 16584
rect 35434 16532 35440 16584
rect 35492 16572 35498 16584
rect 35805 16575 35863 16581
rect 35805 16572 35817 16575
rect 35492 16544 35817 16572
rect 35492 16532 35498 16544
rect 35805 16541 35817 16544
rect 35851 16541 35863 16575
rect 35805 16535 35863 16541
rect 36630 16532 36636 16584
rect 36688 16572 36694 16584
rect 36725 16575 36783 16581
rect 36725 16572 36737 16575
rect 36688 16544 36737 16572
rect 36688 16532 36694 16544
rect 36725 16541 36737 16544
rect 36771 16572 36783 16575
rect 37277 16575 37335 16581
rect 37277 16572 37289 16575
rect 36771 16544 37289 16572
rect 36771 16541 36783 16544
rect 36725 16535 36783 16541
rect 37277 16541 37289 16544
rect 37323 16541 37335 16575
rect 37277 16535 37335 16541
rect 39482 16532 39488 16584
rect 39540 16572 39546 16584
rect 40678 16572 40684 16584
rect 39540 16544 40684 16572
rect 39540 16532 39546 16544
rect 40678 16532 40684 16544
rect 40736 16532 40742 16584
rect 32122 16504 32128 16516
rect 30484 16476 32128 16504
rect 30484 16445 30512 16476
rect 32122 16464 32128 16476
rect 32180 16464 32186 16516
rect 35894 16504 35900 16516
rect 33980 16476 35900 16504
rect 33980 16448 34008 16476
rect 35894 16464 35900 16476
rect 35952 16464 35958 16516
rect 38654 16464 38660 16516
rect 38712 16464 38718 16516
rect 40218 16464 40224 16516
rect 40276 16504 40282 16516
rect 40313 16507 40371 16513
rect 40313 16504 40325 16507
rect 40276 16476 40325 16504
rect 40276 16464 40282 16476
rect 40313 16473 40325 16476
rect 40359 16473 40371 16507
rect 40313 16467 40371 16473
rect 40405 16507 40463 16513
rect 40405 16473 40417 16507
rect 40451 16504 40463 16507
rect 41230 16504 41236 16516
rect 40451 16476 41236 16504
rect 40451 16473 40463 16476
rect 40405 16467 40463 16473
rect 41230 16464 41236 16476
rect 41288 16464 41294 16516
rect 29420 16408 30420 16436
rect 30469 16439 30527 16445
rect 29420 16396 29426 16408
rect 30469 16405 30481 16439
rect 30515 16405 30527 16439
rect 30469 16399 30527 16405
rect 31294 16396 31300 16448
rect 31352 16396 31358 16448
rect 31665 16439 31723 16445
rect 31665 16405 31677 16439
rect 31711 16436 31723 16439
rect 31846 16436 31852 16448
rect 31711 16408 31852 16436
rect 31711 16405 31723 16408
rect 31665 16399 31723 16405
rect 31846 16396 31852 16408
rect 31904 16396 31910 16448
rect 33962 16396 33968 16448
rect 34020 16396 34026 16448
rect 34330 16396 34336 16448
rect 34388 16436 34394 16448
rect 35526 16436 35532 16448
rect 34388 16408 35532 16436
rect 34388 16396 34394 16408
rect 35526 16396 35532 16408
rect 35584 16396 35590 16448
rect 36633 16439 36691 16445
rect 36633 16405 36645 16439
rect 36679 16436 36691 16439
rect 36722 16436 36728 16448
rect 36679 16408 36728 16436
rect 36679 16405 36691 16408
rect 36633 16399 36691 16405
rect 36722 16396 36728 16408
rect 36780 16396 36786 16448
rect 37737 16439 37795 16445
rect 37737 16405 37749 16439
rect 37783 16436 37795 16439
rect 38562 16436 38568 16448
rect 37783 16408 38568 16436
rect 37783 16405 37795 16408
rect 37737 16399 37795 16405
rect 38562 16396 38568 16408
rect 38620 16396 38626 16448
rect 40773 16439 40831 16445
rect 40773 16405 40785 16439
rect 40819 16436 40831 16439
rect 40954 16436 40960 16448
rect 40819 16408 40960 16436
rect 40819 16405 40831 16408
rect 40773 16399 40831 16405
rect 40954 16396 40960 16408
rect 41012 16396 41018 16448
rect 41386 16436 41414 16612
rect 47673 16609 47685 16643
rect 47719 16640 47731 16643
rect 47719 16612 49372 16640
rect 47719 16609 47731 16612
rect 47673 16603 47731 16609
rect 49344 16584 49372 16612
rect 48225 16575 48283 16581
rect 48225 16541 48237 16575
rect 48271 16572 48283 16575
rect 48685 16575 48743 16581
rect 48685 16572 48697 16575
rect 48271 16544 48697 16572
rect 48271 16541 48283 16544
rect 48225 16535 48283 16541
rect 48685 16541 48697 16544
rect 48731 16541 48743 16575
rect 49326 16572 49332 16584
rect 49287 16544 49332 16572
rect 48685 16535 48743 16541
rect 49326 16532 49332 16544
rect 49384 16532 49390 16584
rect 41598 16436 41604 16448
rect 41386 16408 41604 16436
rect 41598 16396 41604 16408
rect 41656 16396 41662 16448
rect 47854 16396 47860 16448
rect 47912 16436 47918 16448
rect 48041 16439 48099 16445
rect 48041 16436 48053 16439
rect 47912 16408 48053 16436
rect 47912 16396 47918 16408
rect 48041 16405 48053 16408
rect 48087 16405 48099 16439
rect 48041 16399 48099 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 8294 16192 8300 16244
rect 8352 16192 8358 16244
rect 9214 16192 9220 16244
rect 9272 16192 9278 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 9824 16204 10977 16232
rect 9824 16192 9830 16204
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 11054 16192 11060 16244
rect 11112 16192 11118 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11977 16235 12035 16241
rect 11977 16232 11989 16235
rect 11388 16204 11989 16232
rect 11388 16192 11394 16204
rect 11977 16201 11989 16204
rect 12023 16201 12035 16235
rect 11977 16195 12035 16201
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 13173 16235 13231 16241
rect 13173 16232 13185 16235
rect 12483 16204 13185 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 13173 16201 13185 16204
rect 13219 16201 13231 16235
rect 14737 16235 14795 16241
rect 14737 16232 14749 16235
rect 13173 16195 13231 16201
rect 13464 16204 14749 16232
rect 10870 16164 10876 16176
rect 2976 16136 10876 16164
rect 2976 16105 3004 16136
rect 10870 16124 10876 16136
rect 10928 16124 10934 16176
rect 11072 16164 11100 16192
rect 13464 16164 13492 16204
rect 14737 16201 14749 16204
rect 14783 16232 14795 16235
rect 15930 16232 15936 16244
rect 14783 16204 15936 16232
rect 14783 16201 14795 16204
rect 14737 16195 14795 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 17402 16192 17408 16244
rect 17460 16192 17466 16244
rect 17773 16235 17831 16241
rect 17773 16201 17785 16235
rect 17819 16232 17831 16235
rect 18322 16232 18328 16244
rect 17819 16204 18328 16232
rect 17819 16201 17831 16204
rect 17773 16195 17831 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18598 16192 18604 16244
rect 18656 16232 18662 16244
rect 23290 16232 23296 16244
rect 18656 16204 23296 16232
rect 18656 16192 18662 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 23400 16204 30328 16232
rect 11072 16136 13492 16164
rect 13541 16167 13599 16173
rect 13541 16133 13553 16167
rect 13587 16164 13599 16167
rect 13587 16136 14044 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 4304 16068 8217 16096
rect 4304 16056 4310 16068
rect 8205 16065 8217 16068
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 11054 16096 11060 16108
rect 10459 16068 11060 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 1026 15988 1032 16040
rect 1084 16028 1090 16040
rect 1765 16031 1823 16037
rect 1765 16028 1777 16031
rect 1084 16000 1777 16028
rect 1084 15988 1090 16000
rect 1765 15997 1777 16000
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 9030 16028 9036 16040
rect 8159 16000 9036 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 9324 16028 9352 16059
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16096 12403 16099
rect 13906 16096 13912 16108
rect 12391 16068 13912 16096
rect 12391 16065 12403 16068
rect 12345 16059 12403 16065
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 9324 16000 10732 16028
rect 8665 15963 8723 15969
rect 8665 15929 8677 15963
rect 8711 15960 8723 15963
rect 9766 15960 9772 15972
rect 8711 15932 9772 15960
rect 8711 15929 8723 15932
rect 8665 15923 8723 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 9916 15864 10517 15892
rect 9916 15852 9922 15864
rect 10505 15861 10517 15864
rect 10551 15892 10563 15895
rect 10594 15892 10600 15904
rect 10551 15864 10600 15892
rect 10551 15861 10563 15864
rect 10505 15855 10563 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 10704 15892 10732 16000
rect 11348 16000 11836 16028
rect 10778 15920 10784 15972
rect 10836 15960 10842 15972
rect 11348 15960 11376 16000
rect 11808 15960 11836 16000
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12621 16031 12679 16037
rect 12621 16028 12633 16031
rect 12492 16000 12633 16028
rect 12492 15988 12498 16000
rect 12621 15997 12633 16000
rect 12667 16028 12679 16031
rect 13446 16028 13452 16040
rect 12667 16000 13452 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 13538 15988 13544 16040
rect 13596 16028 13602 16040
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 13596 16000 13645 16028
rect 13596 15988 13602 16000
rect 13633 15997 13645 16000
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 13722 15988 13728 16040
rect 13780 15988 13786 16040
rect 14016 16028 14044 16136
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 17184 16136 19441 16164
rect 17184 16124 17190 16136
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14792 16068 14964 16096
rect 14792 16056 14798 16068
rect 14016 16000 14412 16028
rect 14274 15960 14280 15972
rect 10836 15932 11376 15960
rect 11440 15932 11744 15960
rect 11808 15932 14280 15960
rect 10836 15920 10842 15932
rect 11440 15892 11468 15932
rect 10704 15864 11468 15892
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11572 15864 11621 15892
rect 11572 15852 11578 15864
rect 11609 15861 11621 15864
rect 11655 15861 11667 15895
rect 11716 15892 11744 15932
rect 14274 15920 14280 15932
rect 14332 15920 14338 15972
rect 14384 15969 14412 16000
rect 14642 15988 14648 16040
rect 14700 16028 14706 16040
rect 14936 16037 14964 16068
rect 15838 16056 15844 16108
rect 15896 16056 15902 16108
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 14829 16031 14887 16037
rect 14829 16028 14841 16031
rect 14700 16000 14841 16028
rect 14700 15988 14706 16000
rect 14829 15997 14841 16000
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15746 15988 15752 16040
rect 15804 15988 15810 16040
rect 14369 15963 14427 15969
rect 14369 15929 14381 15963
rect 14415 15929 14427 15963
rect 14369 15923 14427 15929
rect 14458 15920 14464 15972
rect 14516 15960 14522 15972
rect 15948 15960 15976 16059
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16908 16068 17049 16096
rect 16908 16056 16914 16068
rect 17037 16065 17049 16068
rect 17083 16096 17095 16099
rect 17402 16096 17408 16108
rect 17083 16068 17408 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17402 16056 17408 16068
rect 17460 16056 17466 16108
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17218 16028 17224 16040
rect 16991 16000 17224 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 17972 16037 18000 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 20714 16164 20720 16176
rect 20654 16136 20720 16164
rect 19429 16127 19487 16133
rect 20714 16124 20720 16136
rect 20772 16164 20778 16176
rect 21634 16164 21640 16176
rect 20772 16136 21640 16164
rect 20772 16124 20778 16136
rect 21634 16124 21640 16136
rect 21692 16124 21698 16176
rect 18874 16056 18880 16108
rect 18932 16096 18938 16108
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 18932 16068 19165 16096
rect 18932 16056 18938 16068
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 23400 16096 23428 16204
rect 24578 16124 24584 16176
rect 24636 16164 24642 16176
rect 27798 16164 27804 16176
rect 24636 16136 24886 16164
rect 26344 16136 27804 16164
rect 24636 16124 24642 16136
rect 19153 16059 19211 16065
rect 20640 16068 23428 16096
rect 23477 16099 23535 16105
rect 17865 16031 17923 16037
rect 17865 15997 17877 16031
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 15997 18015 16031
rect 19978 16028 19984 16040
rect 17957 15991 18015 15997
rect 18064 16000 19984 16028
rect 14516 15932 15976 15960
rect 16301 15963 16359 15969
rect 14516 15920 14522 15932
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 17586 15960 17592 15972
rect 16347 15932 17592 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 17586 15920 17592 15932
rect 17644 15920 17650 15972
rect 17880 15960 17908 15991
rect 18064 15960 18092 16000
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 18877 15963 18935 15969
rect 18877 15960 18889 15963
rect 17880 15932 18092 15960
rect 18340 15932 18889 15960
rect 16482 15892 16488 15904
rect 11716 15864 16488 15892
rect 11609 15855 11667 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 16761 15895 16819 15901
rect 16761 15861 16773 15895
rect 16807 15892 16819 15895
rect 16942 15892 16948 15904
rect 16807 15864 16948 15892
rect 16807 15861 16819 15864
rect 16761 15855 16819 15861
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 18340 15892 18368 15932
rect 18877 15929 18889 15932
rect 18923 15960 18935 15963
rect 19058 15960 19064 15972
rect 18923 15932 19064 15960
rect 18923 15929 18935 15932
rect 18877 15923 18935 15929
rect 19058 15920 19064 15932
rect 19116 15920 19122 15972
rect 17368 15864 18368 15892
rect 17368 15852 17374 15864
rect 18414 15852 18420 15904
rect 18472 15892 18478 15904
rect 18782 15892 18788 15904
rect 18472 15864 18788 15892
rect 18472 15852 18478 15864
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 20640 15892 20668 16068
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23566 16096 23572 16108
rect 23523 16068 23572 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23566 16056 23572 16068
rect 23624 16056 23630 16108
rect 26344 16105 26372 16136
rect 27798 16124 27804 16136
rect 27856 16164 27862 16176
rect 28902 16164 28908 16176
rect 27856 16136 28908 16164
rect 27856 16124 27862 16136
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 26602 16056 26608 16108
rect 26660 16096 26666 16108
rect 27522 16096 27528 16108
rect 26660 16068 27528 16096
rect 26660 16056 26666 16068
rect 27522 16056 27528 16068
rect 27580 16056 27586 16108
rect 27617 16099 27675 16105
rect 27617 16065 27629 16099
rect 27663 16096 27675 16099
rect 28258 16096 28264 16108
rect 27663 16068 28264 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 28258 16056 28264 16068
rect 28316 16056 28322 16108
rect 28368 16105 28396 16136
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 29086 16124 29092 16176
rect 29144 16124 29150 16176
rect 30300 16164 30328 16204
rect 30374 16192 30380 16244
rect 30432 16232 30438 16244
rect 30929 16235 30987 16241
rect 30929 16232 30941 16235
rect 30432 16204 30941 16232
rect 30432 16192 30438 16204
rect 30929 16201 30941 16204
rect 30975 16201 30987 16235
rect 30929 16195 30987 16201
rect 31754 16192 31760 16244
rect 31812 16232 31818 16244
rect 33781 16235 33839 16241
rect 33781 16232 33793 16235
rect 31812 16204 33793 16232
rect 31812 16192 31818 16204
rect 33781 16201 33793 16204
rect 33827 16201 33839 16235
rect 33781 16195 33839 16201
rect 34790 16192 34796 16244
rect 34848 16232 34854 16244
rect 34848 16204 36952 16232
rect 34848 16192 34854 16204
rect 30650 16164 30656 16176
rect 30300 16136 30656 16164
rect 30650 16124 30656 16136
rect 30708 16124 30714 16176
rect 30834 16124 30840 16176
rect 30892 16124 30898 16176
rect 32585 16167 32643 16173
rect 32585 16133 32597 16167
rect 32631 16164 32643 16167
rect 34517 16167 34575 16173
rect 34517 16164 34529 16167
rect 32631 16136 34529 16164
rect 32631 16133 32643 16136
rect 32585 16127 32643 16133
rect 34517 16133 34529 16136
rect 34563 16133 34575 16167
rect 34517 16127 34575 16133
rect 28353 16099 28411 16105
rect 28353 16065 28365 16099
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 20806 15988 20812 16040
rect 20864 16028 20870 16040
rect 20901 16031 20959 16037
rect 20901 16028 20913 16031
rect 20864 16000 20913 16028
rect 20864 15988 20870 16000
rect 20901 15997 20913 16000
rect 20947 16028 20959 16031
rect 21910 16028 21916 16040
rect 20947 16000 21916 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 23293 16031 23351 16037
rect 23293 15997 23305 16031
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 16028 23443 16031
rect 24486 16028 24492 16040
rect 23431 16000 23520 16028
rect 23431 15997 23443 16000
rect 23385 15991 23443 15997
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 22186 15960 22192 15972
rect 20772 15932 22192 15960
rect 20772 15920 20778 15932
rect 22186 15920 22192 15932
rect 22244 15920 22250 15972
rect 19208 15864 20668 15892
rect 19208 15852 19214 15864
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 21545 15895 21603 15901
rect 21545 15861 21557 15895
rect 21591 15892 21603 15895
rect 21634 15892 21640 15904
rect 21591 15864 21640 15892
rect 21591 15861 21603 15864
rect 21545 15855 21603 15861
rect 21634 15852 21640 15864
rect 21692 15892 21698 15904
rect 22741 15895 22799 15901
rect 22741 15892 22753 15895
rect 21692 15864 22753 15892
rect 21692 15852 21698 15864
rect 22741 15861 22753 15864
rect 22787 15861 22799 15895
rect 23308 15892 23336 15991
rect 23492 15972 23520 16000
rect 23584 16000 24492 16028
rect 23474 15920 23480 15972
rect 23532 15920 23538 15972
rect 23584 15892 23612 16000
rect 24486 15988 24492 16000
rect 24544 16028 24550 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24544 16000 24593 16028
rect 24544 15988 24550 16000
rect 24581 15997 24593 16000
rect 24627 15997 24639 16031
rect 24581 15991 24639 15997
rect 26053 16031 26111 16037
rect 26053 15997 26065 16031
rect 26099 16028 26111 16031
rect 26786 16028 26792 16040
rect 26099 16000 26792 16028
rect 26099 15997 26111 16000
rect 26053 15991 26111 15997
rect 26786 15988 26792 16000
rect 26844 15988 26850 16040
rect 27430 16028 27436 16040
rect 26896 16000 27436 16028
rect 23845 15963 23903 15969
rect 23845 15929 23857 15963
rect 23891 15960 23903 15963
rect 24670 15960 24676 15972
rect 23891 15932 24676 15960
rect 23891 15929 23903 15932
rect 23845 15923 23903 15929
rect 24670 15920 24676 15932
rect 24728 15920 24734 15972
rect 26697 15963 26755 15969
rect 26697 15929 26709 15963
rect 26743 15960 26755 15963
rect 26896 15960 26924 16000
rect 27430 15988 27436 16000
rect 27488 15988 27494 16040
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 26743 15932 26924 15960
rect 26743 15929 26755 15932
rect 26697 15923 26755 15929
rect 26970 15920 26976 15972
rect 27028 15960 27034 15972
rect 27724 15960 27752 15991
rect 28626 15988 28632 16040
rect 28684 15988 28690 16040
rect 29822 15988 29828 16040
rect 29880 16028 29886 16040
rect 30653 16031 30711 16037
rect 30653 16028 30665 16031
rect 29880 16000 30665 16028
rect 29880 15988 29886 16000
rect 30653 15997 30665 16000
rect 30699 15997 30711 16031
rect 30653 15991 30711 15997
rect 31849 16031 31907 16037
rect 31849 15997 31861 16031
rect 31895 16028 31907 16031
rect 31938 16028 31944 16040
rect 31895 16000 31944 16028
rect 31895 15997 31907 16000
rect 31849 15991 31907 15997
rect 31938 15988 31944 16000
rect 31996 15988 32002 16040
rect 32214 15988 32220 16040
rect 32272 16028 32278 16040
rect 32401 16031 32459 16037
rect 32401 16028 32413 16031
rect 32272 16000 32413 16028
rect 32272 15988 32278 16000
rect 32401 15997 32413 16000
rect 32447 15997 32459 16031
rect 32401 15991 32459 15997
rect 32600 15960 32628 16127
rect 36170 16124 36176 16176
rect 36228 16124 36234 16176
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16065 32735 16099
rect 32677 16059 32735 16065
rect 27028 15932 27752 15960
rect 29656 15932 32628 15960
rect 32692 15960 32720 16059
rect 33318 16056 33324 16108
rect 33376 16096 33382 16108
rect 36924 16105 36952 16204
rect 36998 16192 37004 16244
rect 37056 16232 37062 16244
rect 40497 16235 40555 16241
rect 40497 16232 40509 16235
rect 37056 16204 40509 16232
rect 37056 16192 37062 16204
rect 40497 16201 40509 16204
rect 40543 16201 40555 16235
rect 40497 16195 40555 16201
rect 40954 16192 40960 16244
rect 41012 16192 41018 16244
rect 38473 16167 38531 16173
rect 38473 16133 38485 16167
rect 38519 16164 38531 16167
rect 38562 16164 38568 16176
rect 38519 16136 38568 16164
rect 38519 16133 38531 16136
rect 38473 16127 38531 16133
rect 38562 16124 38568 16136
rect 38620 16124 38626 16176
rect 38746 16124 38752 16176
rect 38804 16164 38810 16176
rect 38804 16136 38962 16164
rect 38804 16124 38810 16136
rect 33873 16099 33931 16105
rect 33873 16096 33885 16099
rect 33376 16068 33885 16096
rect 33376 16056 33382 16068
rect 33873 16065 33885 16068
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 36909 16099 36967 16105
rect 36909 16065 36921 16099
rect 36955 16096 36967 16099
rect 37366 16096 37372 16108
rect 36955 16068 37372 16096
rect 36955 16065 36967 16068
rect 36909 16059 36967 16065
rect 37366 16056 37372 16068
rect 37424 16096 37430 16108
rect 38197 16099 38255 16105
rect 38197 16096 38209 16099
rect 37424 16068 38209 16096
rect 37424 16056 37430 16068
rect 38197 16065 38209 16068
rect 38243 16065 38255 16099
rect 38197 16059 38255 16065
rect 40865 16099 40923 16105
rect 40865 16065 40877 16099
rect 40911 16096 40923 16099
rect 48314 16096 48320 16108
rect 40911 16068 48320 16096
rect 40911 16065 40923 16068
rect 40865 16059 40923 16065
rect 48314 16056 48320 16068
rect 48372 16056 48378 16108
rect 48409 16099 48467 16105
rect 48409 16065 48421 16099
rect 48455 16096 48467 16099
rect 48682 16096 48688 16108
rect 48455 16068 48688 16096
rect 48455 16065 48467 16068
rect 48409 16059 48467 16065
rect 48682 16056 48688 16068
rect 48740 16056 48746 16108
rect 32766 15988 32772 16040
rect 32824 16028 32830 16040
rect 33597 16031 33655 16037
rect 33597 16028 33609 16031
rect 32824 16000 33609 16028
rect 32824 15988 32830 16000
rect 33597 15997 33609 16000
rect 33643 15997 33655 16031
rect 33597 15991 33655 15997
rect 36633 16031 36691 16037
rect 36633 15997 36645 16031
rect 36679 16028 36691 16031
rect 36679 16000 37136 16028
rect 36679 15997 36691 16000
rect 36633 15991 36691 15997
rect 33410 15960 33416 15972
rect 32692 15932 33416 15960
rect 27028 15920 27034 15932
rect 23308 15864 23612 15892
rect 22741 15855 22799 15861
rect 26878 15852 26884 15904
rect 26936 15892 26942 15904
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 26936 15864 27169 15892
rect 26936 15852 26942 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27157 15855 27215 15861
rect 27338 15852 27344 15904
rect 27396 15892 27402 15904
rect 29656 15892 29684 15932
rect 33410 15920 33416 15932
rect 33468 15960 33474 15972
rect 34241 15963 34299 15969
rect 33468 15932 34192 15960
rect 33468 15920 33474 15932
rect 34164 15904 34192 15932
rect 34241 15929 34253 15963
rect 34287 15960 34299 15963
rect 37108 15960 37136 16000
rect 37458 15988 37464 16040
rect 37516 15988 37522 16040
rect 38562 15988 38568 16040
rect 38620 16028 38626 16040
rect 41049 16031 41107 16037
rect 41049 16028 41061 16031
rect 38620 16000 41061 16028
rect 38620 15988 38626 16000
rect 41049 15997 41061 16000
rect 41095 16028 41107 16031
rect 41782 16028 41788 16040
rect 41095 16000 41788 16028
rect 41095 15997 41107 16000
rect 41049 15991 41107 15997
rect 41782 15988 41788 16000
rect 41840 15988 41846 16040
rect 37642 15960 37648 15972
rect 34287 15932 35664 15960
rect 37108 15932 37648 15960
rect 34287 15929 34299 15932
rect 34241 15923 34299 15929
rect 27396 15864 29684 15892
rect 30101 15895 30159 15901
rect 27396 15852 27402 15864
rect 30101 15861 30113 15895
rect 30147 15892 30159 15895
rect 30742 15892 30748 15904
rect 30147 15864 30748 15892
rect 30147 15861 30159 15864
rect 30101 15855 30159 15861
rect 30742 15852 30748 15864
rect 30800 15852 30806 15904
rect 31297 15895 31355 15901
rect 31297 15861 31309 15895
rect 31343 15892 31355 15895
rect 31386 15892 31392 15904
rect 31343 15864 31392 15892
rect 31343 15861 31355 15864
rect 31297 15855 31355 15861
rect 31386 15852 31392 15864
rect 31444 15852 31450 15904
rect 31665 15895 31723 15901
rect 31665 15861 31677 15895
rect 31711 15892 31723 15895
rect 31754 15892 31760 15904
rect 31711 15864 31760 15892
rect 31711 15861 31723 15864
rect 31665 15855 31723 15861
rect 31754 15852 31760 15864
rect 31812 15852 31818 15904
rect 33045 15895 33103 15901
rect 33045 15861 33057 15895
rect 33091 15892 33103 15895
rect 33686 15892 33692 15904
rect 33091 15864 33692 15892
rect 33091 15861 33103 15864
rect 33045 15855 33103 15861
rect 33686 15852 33692 15864
rect 33744 15852 33750 15904
rect 34146 15852 34152 15904
rect 34204 15892 34210 15904
rect 34701 15895 34759 15901
rect 34701 15892 34713 15895
rect 34204 15864 34713 15892
rect 34204 15852 34210 15864
rect 34701 15861 34713 15864
rect 34747 15861 34759 15895
rect 34701 15855 34759 15861
rect 35158 15852 35164 15904
rect 35216 15852 35222 15904
rect 35636 15892 35664 15932
rect 37642 15920 37648 15932
rect 37700 15920 37706 15972
rect 37182 15892 37188 15904
rect 35636 15864 37188 15892
rect 37182 15852 37188 15864
rect 37240 15852 37246 15904
rect 39945 15895 40003 15901
rect 39945 15861 39957 15895
rect 39991 15892 40003 15895
rect 40310 15892 40316 15904
rect 39991 15864 40316 15892
rect 39991 15861 40003 15864
rect 39945 15855 40003 15861
rect 40310 15852 40316 15864
rect 40368 15852 40374 15904
rect 41598 15852 41604 15904
rect 41656 15852 41662 15904
rect 49326 15852 49332 15904
rect 49384 15852 49390 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10744 15660 10793 15688
rect 10744 15648 10750 15660
rect 10781 15657 10793 15660
rect 10827 15688 10839 15691
rect 12434 15688 12440 15700
rect 10827 15660 12440 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 12986 15648 12992 15700
rect 13044 15688 13050 15700
rect 14366 15688 14372 15700
rect 13044 15660 14372 15688
rect 13044 15648 13050 15660
rect 14366 15648 14372 15660
rect 14424 15688 14430 15700
rect 14918 15688 14924 15700
rect 14424 15660 14924 15688
rect 14424 15648 14430 15660
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 16758 15648 16764 15700
rect 16816 15648 16822 15700
rect 17862 15648 17868 15700
rect 17920 15648 17926 15700
rect 18049 15691 18107 15697
rect 18049 15657 18061 15691
rect 18095 15688 18107 15691
rect 18690 15688 18696 15700
rect 18095 15660 18696 15688
rect 18095 15657 18107 15660
rect 18049 15651 18107 15657
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 18969 15691 19027 15697
rect 18969 15688 18981 15691
rect 18840 15660 18981 15688
rect 18840 15648 18846 15660
rect 18969 15657 18981 15660
rect 19015 15657 19027 15691
rect 18969 15651 19027 15657
rect 19058 15648 19064 15700
rect 19116 15688 19122 15700
rect 19334 15688 19340 15700
rect 19116 15660 19340 15688
rect 19116 15648 19122 15660
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 19886 15648 19892 15700
rect 19944 15648 19950 15700
rect 20898 15648 20904 15700
rect 20956 15688 20962 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20956 15660 21189 15688
rect 20956 15648 20962 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 21177 15651 21235 15657
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 25130 15688 25136 15700
rect 22612 15660 25136 15688
rect 22612 15648 22618 15660
rect 25130 15648 25136 15660
rect 25188 15688 25194 15700
rect 26142 15688 26148 15700
rect 25188 15660 26148 15688
rect 25188 15648 25194 15660
rect 26142 15648 26148 15660
rect 26200 15648 26206 15700
rect 26234 15648 26240 15700
rect 26292 15688 26298 15700
rect 26973 15691 27031 15697
rect 26973 15688 26985 15691
rect 26292 15660 26985 15688
rect 26292 15648 26298 15660
rect 26973 15657 26985 15660
rect 27019 15688 27031 15691
rect 27062 15688 27068 15700
rect 27019 15660 27068 15688
rect 27019 15657 27031 15660
rect 26973 15651 27031 15657
rect 27062 15648 27068 15660
rect 27120 15648 27126 15700
rect 28537 15691 28595 15697
rect 28537 15657 28549 15691
rect 28583 15688 28595 15691
rect 28810 15688 28816 15700
rect 28583 15660 28816 15688
rect 28583 15657 28595 15660
rect 28537 15651 28595 15657
rect 28810 15648 28816 15660
rect 28868 15648 28874 15700
rect 29086 15648 29092 15700
rect 29144 15688 29150 15700
rect 29273 15691 29331 15697
rect 29273 15688 29285 15691
rect 29144 15660 29285 15688
rect 29144 15648 29150 15660
rect 29273 15657 29285 15660
rect 29319 15657 29331 15691
rect 29273 15651 29331 15657
rect 29546 15648 29552 15700
rect 29604 15688 29610 15700
rect 29604 15660 32996 15688
rect 29604 15648 29610 15660
rect 13722 15620 13728 15632
rect 12452 15592 13728 15620
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15552 10563 15555
rect 11054 15552 11060 15564
rect 10551 15524 11060 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12452 15552 12480 15592
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 13906 15580 13912 15632
rect 13964 15620 13970 15632
rect 15010 15620 15016 15632
rect 13964 15592 15016 15620
rect 13964 15580 13970 15592
rect 15010 15580 15016 15592
rect 15068 15580 15074 15632
rect 16482 15580 16488 15632
rect 16540 15620 16546 15632
rect 18417 15623 18475 15629
rect 18417 15620 18429 15623
rect 16540 15592 18429 15620
rect 16540 15580 16546 15592
rect 18417 15589 18429 15592
rect 18463 15589 18475 15623
rect 22281 15623 22339 15629
rect 22281 15620 22293 15623
rect 18417 15583 18475 15589
rect 20456 15592 22293 15620
rect 12299 15524 12480 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12526 15512 12532 15564
rect 12584 15512 12590 15564
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15552 13231 15555
rect 14458 15552 14464 15564
rect 13219 15524 14464 15552
rect 13219 15521 13231 15524
rect 13173 15515 13231 15521
rect 14458 15512 14464 15524
rect 14516 15512 14522 15564
rect 14826 15512 14832 15564
rect 14884 15512 14890 15564
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 15804 15524 16129 15552
rect 15804 15512 15810 15524
rect 16117 15521 16129 15524
rect 16163 15521 16175 15555
rect 16117 15515 16175 15521
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 10226 15484 10232 15496
rect 3007 15456 10232 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 12544 15484 12572 15512
rect 15102 15484 15108 15496
rect 12544 15456 15108 15484
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15930 15444 15936 15496
rect 15988 15444 15994 15496
rect 16022 15444 16028 15496
rect 16080 15484 16086 15496
rect 17328 15484 17356 15515
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 20456 15552 20484 15592
rect 17460 15524 20484 15552
rect 20533 15555 20591 15561
rect 17460 15512 17466 15524
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 21358 15552 21364 15564
rect 20579 15524 21364 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 21729 15555 21787 15561
rect 21729 15552 21741 15555
rect 21508 15524 21741 15552
rect 21508 15512 21514 15524
rect 21729 15521 21741 15524
rect 21775 15521 21787 15555
rect 21729 15515 21787 15521
rect 16080 15456 17356 15484
rect 16080 15444 16086 15456
rect 18414 15444 18420 15496
rect 18472 15444 18478 15496
rect 18598 15444 18604 15496
rect 18656 15444 18662 15496
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 21542 15484 21548 15496
rect 19024 15456 21548 15484
rect 19024 15444 19030 15456
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 21836 15484 21864 15592
rect 22281 15589 22293 15592
rect 22327 15620 22339 15623
rect 24854 15620 24860 15632
rect 22327 15592 24860 15620
rect 22327 15589 22339 15592
rect 22281 15583 22339 15589
rect 24854 15580 24860 15592
rect 24912 15580 24918 15632
rect 26694 15620 26700 15632
rect 25240 15592 26700 15620
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 23661 15555 23719 15561
rect 23661 15552 23673 15555
rect 22152 15524 23673 15552
rect 22152 15512 22158 15524
rect 23661 15521 23673 15524
rect 23707 15521 23719 15555
rect 23661 15515 23719 15521
rect 24302 15512 24308 15564
rect 24360 15552 24366 15564
rect 25240 15561 25268 15592
rect 26694 15580 26700 15592
rect 26752 15580 26758 15632
rect 32217 15623 32275 15629
rect 32217 15589 32229 15623
rect 32263 15620 32275 15623
rect 32582 15620 32588 15632
rect 32263 15592 32588 15620
rect 32263 15589 32275 15592
rect 32217 15583 32275 15589
rect 32582 15580 32588 15592
rect 32640 15580 32646 15632
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 24360 15524 25237 15552
rect 24360 15512 24366 15524
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25225 15515 25283 15521
rect 25314 15512 25320 15564
rect 25372 15552 25378 15564
rect 26421 15555 26479 15561
rect 26421 15552 26433 15555
rect 25372 15524 26433 15552
rect 25372 15512 25378 15524
rect 26421 15521 26433 15524
rect 26467 15521 26479 15555
rect 26421 15515 26479 15521
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 26660 15524 27997 15552
rect 26660 15512 26666 15524
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 30469 15555 30527 15561
rect 30469 15521 30481 15555
rect 30515 15552 30527 15555
rect 31110 15552 31116 15564
rect 30515 15524 31116 15552
rect 30515 15521 30527 15524
rect 30469 15515 30527 15521
rect 31110 15512 31116 15524
rect 31168 15512 31174 15564
rect 32968 15561 32996 15660
rect 34422 15648 34428 15700
rect 34480 15648 34486 15700
rect 36633 15691 36691 15697
rect 36633 15657 36645 15691
rect 36679 15688 36691 15691
rect 37642 15688 37648 15700
rect 36679 15660 37648 15688
rect 36679 15657 36691 15660
rect 36633 15651 36691 15657
rect 37642 15648 37648 15660
rect 37700 15648 37706 15700
rect 37734 15648 37740 15700
rect 37792 15648 37798 15700
rect 41598 15648 41604 15700
rect 41656 15688 41662 15700
rect 42061 15691 42119 15697
rect 42061 15688 42073 15691
rect 41656 15660 42073 15688
rect 41656 15648 41662 15660
rect 42061 15657 42073 15660
rect 42107 15657 42119 15691
rect 42061 15651 42119 15657
rect 48314 15648 48320 15700
rect 48372 15688 48378 15700
rect 48409 15691 48467 15697
rect 48409 15688 48421 15691
rect 48372 15660 48421 15688
rect 48372 15648 48378 15660
rect 48409 15657 48421 15660
rect 48455 15657 48467 15691
rect 48409 15651 48467 15657
rect 49142 15648 49148 15700
rect 49200 15648 49206 15700
rect 41782 15580 41788 15632
rect 41840 15580 41846 15632
rect 32861 15555 32919 15561
rect 32861 15521 32873 15555
rect 32907 15521 32919 15555
rect 32861 15515 32919 15521
rect 32953 15555 33011 15561
rect 32953 15521 32965 15555
rect 32999 15521 33011 15555
rect 32953 15515 33011 15521
rect 21683 15456 21864 15484
rect 23569 15487 23627 15493
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 27154 15484 27160 15496
rect 23615 15456 27160 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27893 15487 27951 15493
rect 27893 15453 27905 15487
rect 27939 15484 27951 15487
rect 28166 15484 28172 15496
rect 27939 15456 28172 15484
rect 27939 15453 27951 15456
rect 27893 15447 27951 15453
rect 28166 15444 28172 15456
rect 28224 15484 28230 15496
rect 28629 15487 28687 15493
rect 28629 15484 28641 15487
rect 28224 15456 28641 15484
rect 28224 15444 28230 15456
rect 28629 15453 28641 15456
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15484 29239 15487
rect 30098 15484 30104 15496
rect 29227 15456 30104 15484
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 30098 15444 30104 15456
rect 30156 15444 30162 15496
rect 32876 15484 32904 15515
rect 34790 15512 34796 15564
rect 34848 15552 34854 15564
rect 34885 15555 34943 15561
rect 34885 15552 34897 15555
rect 34848 15524 34897 15552
rect 34848 15512 34854 15524
rect 34885 15521 34897 15524
rect 34931 15521 34943 15555
rect 34885 15515 34943 15521
rect 35161 15555 35219 15561
rect 35161 15521 35173 15555
rect 35207 15552 35219 15555
rect 35894 15552 35900 15564
rect 35207 15524 35900 15552
rect 35207 15521 35219 15524
rect 35161 15515 35219 15521
rect 35894 15512 35900 15524
rect 35952 15512 35958 15564
rect 36170 15512 36176 15564
rect 36228 15552 36234 15564
rect 36446 15552 36452 15564
rect 36228 15524 36452 15552
rect 36228 15512 36234 15524
rect 34330 15484 34336 15496
rect 32876 15456 34336 15484
rect 34330 15444 34336 15456
rect 34388 15444 34394 15496
rect 36280 15470 36308 15524
rect 36446 15512 36452 15524
rect 36504 15512 36510 15564
rect 37366 15512 37372 15564
rect 37424 15552 37430 15564
rect 39482 15552 39488 15564
rect 37424 15524 39488 15552
rect 37424 15512 37430 15524
rect 39482 15512 39488 15524
rect 39540 15552 39546 15564
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 39540 15524 40049 15552
rect 39540 15512 39546 15524
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 40310 15512 40316 15564
rect 40368 15512 40374 15564
rect 48133 15487 48191 15493
rect 48133 15453 48145 15487
rect 48179 15484 48191 15487
rect 48590 15484 48596 15496
rect 48179 15456 48596 15484
rect 48179 15453 48191 15456
rect 48133 15447 48191 15453
rect 48590 15444 48596 15456
rect 48648 15444 48654 15496
rect 49326 15444 49332 15496
rect 49384 15444 49390 15496
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 1765 15419 1823 15425
rect 1765 15416 1777 15419
rect 992 15388 1777 15416
rect 992 15376 998 15388
rect 1765 15385 1777 15388
rect 1811 15385 1823 15419
rect 1765 15379 1823 15385
rect 4154 15376 4160 15428
rect 4212 15416 4218 15428
rect 6365 15419 6423 15425
rect 6365 15416 6377 15419
rect 4212 15388 6377 15416
rect 4212 15376 4218 15388
rect 6365 15385 6377 15388
rect 6411 15385 6423 15419
rect 6365 15379 6423 15385
rect 6549 15419 6607 15425
rect 6549 15385 6561 15419
rect 6595 15416 6607 15419
rect 6595 15388 10364 15416
rect 11822 15388 12572 15416
rect 6595 15385 6607 15388
rect 6549 15379 6607 15385
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 10336 15348 10364 15388
rect 11238 15348 11244 15360
rect 10336 15320 11244 15348
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 12544 15348 12572 15388
rect 12618 15376 12624 15428
rect 12676 15416 12682 15428
rect 13265 15419 13323 15425
rect 13265 15416 13277 15419
rect 12676 15388 13277 15416
rect 12676 15376 12682 15388
rect 13265 15385 13277 15388
rect 13311 15385 13323 15419
rect 13265 15379 13323 15385
rect 13354 15376 13360 15428
rect 13412 15376 13418 15428
rect 14737 15419 14795 15425
rect 14737 15385 14749 15419
rect 14783 15416 14795 15419
rect 18432 15416 18460 15444
rect 14783 15388 18460 15416
rect 20349 15419 20407 15425
rect 14783 15385 14795 15388
rect 14737 15379 14795 15385
rect 20349 15385 20361 15419
rect 20395 15416 20407 15419
rect 23477 15419 23535 15425
rect 20395 15388 23152 15416
rect 20395 15385 20407 15388
rect 20349 15379 20407 15385
rect 12986 15348 12992 15360
rect 12544 15320 12992 15348
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 13538 15308 13544 15360
rect 13596 15348 13602 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13596 15320 13737 15348
rect 13596 15308 13602 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 13872 15320 14289 15348
rect 13872 15308 13878 15320
rect 14277 15317 14289 15320
rect 14323 15317 14335 15351
rect 14277 15311 14335 15317
rect 14550 15308 14556 15360
rect 14608 15348 14614 15360
rect 14645 15351 14703 15357
rect 14645 15348 14657 15351
rect 14608 15320 14657 15348
rect 14608 15308 14614 15320
rect 14645 15317 14657 15320
rect 14691 15317 14703 15351
rect 14645 15311 14703 15317
rect 15562 15308 15568 15360
rect 15620 15308 15626 15360
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 16025 15351 16083 15357
rect 16025 15348 16037 15351
rect 15804 15320 16037 15348
rect 15804 15308 15810 15320
rect 16025 15317 16037 15320
rect 16071 15317 16083 15351
rect 16025 15311 16083 15317
rect 17126 15308 17132 15360
rect 17184 15308 17190 15360
rect 17221 15351 17279 15357
rect 17221 15317 17233 15351
rect 17267 15348 17279 15351
rect 17862 15348 17868 15360
rect 17267 15320 17868 15348
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 19702 15348 19708 15360
rect 19567 15320 19708 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 20254 15308 20260 15360
rect 20312 15308 20318 15360
rect 21266 15308 21272 15360
rect 21324 15348 21330 15360
rect 21450 15348 21456 15360
rect 21324 15320 21456 15348
rect 21324 15308 21330 15320
rect 21450 15308 21456 15320
rect 21508 15348 21514 15360
rect 23124 15357 23152 15388
rect 23477 15385 23489 15419
rect 23523 15416 23535 15419
rect 23523 15388 24716 15416
rect 23523 15385 23535 15388
rect 23477 15379 23535 15385
rect 21545 15351 21603 15357
rect 21545 15348 21557 15351
rect 21508 15320 21557 15348
rect 21508 15308 21514 15320
rect 21545 15317 21557 15320
rect 21591 15317 21603 15351
rect 21545 15311 21603 15317
rect 23109 15351 23167 15357
rect 23109 15317 23121 15351
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 24118 15308 24124 15360
rect 24176 15308 24182 15360
rect 24688 15357 24716 15388
rect 25038 15376 25044 15428
rect 25096 15416 25102 15428
rect 25682 15416 25688 15428
rect 25096 15388 25688 15416
rect 25096 15376 25102 15388
rect 25682 15376 25688 15388
rect 25740 15376 25746 15428
rect 26234 15376 26240 15428
rect 26292 15376 26298 15428
rect 26326 15376 26332 15428
rect 26384 15416 26390 15428
rect 27801 15419 27859 15425
rect 26384 15388 27200 15416
rect 26384 15376 26390 15388
rect 27172 15360 27200 15388
rect 27801 15385 27813 15419
rect 27847 15416 27859 15419
rect 28810 15416 28816 15428
rect 27847 15388 28816 15416
rect 27847 15385 27859 15388
rect 27801 15379 27859 15385
rect 28810 15376 28816 15388
rect 28868 15376 28874 15428
rect 28997 15419 29055 15425
rect 28997 15385 29009 15419
rect 29043 15416 29055 15419
rect 30466 15416 30472 15428
rect 29043 15388 30472 15416
rect 29043 15385 29055 15388
rect 28997 15379 29055 15385
rect 30466 15376 30472 15388
rect 30524 15376 30530 15428
rect 30742 15376 30748 15428
rect 30800 15376 30806 15428
rect 31754 15376 31760 15428
rect 31812 15376 31818 15428
rect 34882 15416 34888 15428
rect 33428 15388 34888 15416
rect 24673 15351 24731 15357
rect 24673 15317 24685 15351
rect 24719 15317 24731 15351
rect 24673 15311 24731 15317
rect 25130 15308 25136 15360
rect 25188 15308 25194 15360
rect 25866 15308 25872 15360
rect 25924 15308 25930 15360
rect 26786 15308 26792 15360
rect 26844 15348 26850 15360
rect 27065 15351 27123 15357
rect 27065 15348 27077 15351
rect 26844 15320 27077 15348
rect 26844 15308 26850 15320
rect 27065 15317 27077 15320
rect 27111 15317 27123 15351
rect 27065 15311 27123 15317
rect 27154 15308 27160 15360
rect 27212 15308 27218 15360
rect 27430 15308 27436 15360
rect 27488 15308 27494 15360
rect 30006 15308 30012 15360
rect 30064 15308 30070 15360
rect 30282 15308 30288 15360
rect 30340 15348 30346 15360
rect 31662 15348 31668 15360
rect 30340 15320 31668 15348
rect 30340 15308 30346 15320
rect 31662 15308 31668 15320
rect 31720 15308 31726 15360
rect 32030 15308 32036 15360
rect 32088 15348 32094 15360
rect 33042 15348 33048 15360
rect 32088 15320 33048 15348
rect 32088 15308 32094 15320
rect 33042 15308 33048 15320
rect 33100 15308 33106 15360
rect 33428 15357 33456 15388
rect 34882 15376 34888 15388
rect 34940 15376 34946 15428
rect 38746 15376 38752 15428
rect 38804 15376 38810 15428
rect 39209 15419 39267 15425
rect 39209 15385 39221 15419
rect 39255 15385 39267 15419
rect 39209 15379 39267 15385
rect 33413 15351 33471 15357
rect 33413 15317 33425 15351
rect 33459 15317 33471 15351
rect 33413 15311 33471 15317
rect 33870 15308 33876 15360
rect 33928 15308 33934 15360
rect 35894 15308 35900 15360
rect 35952 15348 35958 15360
rect 37093 15351 37151 15357
rect 37093 15348 37105 15351
rect 35952 15320 37105 15348
rect 35952 15308 35958 15320
rect 37093 15317 37105 15320
rect 37139 15317 37151 15351
rect 37093 15311 37151 15317
rect 37826 15308 37832 15360
rect 37884 15348 37890 15360
rect 38562 15348 38568 15360
rect 37884 15320 38568 15348
rect 37884 15308 37890 15320
rect 38562 15308 38568 15320
rect 38620 15348 38626 15360
rect 39224 15348 39252 15379
rect 41046 15376 41052 15428
rect 41104 15376 41110 15428
rect 38620 15320 39252 15348
rect 38620 15308 38626 15320
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 9674 15104 9680 15156
rect 9732 15104 9738 15156
rect 9766 15104 9772 15156
rect 9824 15104 9830 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11790 15144 11796 15156
rect 11296 15116 11796 15144
rect 11296 15104 11302 15116
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 11882 15104 11888 15156
rect 11940 15104 11946 15156
rect 12986 15104 12992 15156
rect 13044 15104 13050 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 13906 15144 13912 15156
rect 13403 15116 13912 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 13906 15104 13912 15116
rect 13964 15144 13970 15156
rect 13964 15116 14504 15144
rect 13964 15104 13970 15116
rect 10870 15036 10876 15088
rect 10928 15036 10934 15088
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 11112 15048 12848 15076
rect 11112 15036 11118 15048
rect 934 14968 940 15020
rect 992 15008 998 15020
rect 1765 15011 1823 15017
rect 1765 15008 1777 15011
rect 992 14980 1777 15008
rect 992 14968 998 14980
rect 1765 14977 1777 14980
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 4154 15008 4160 15020
rect 3007 14980 4160 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 10744 14980 12265 15008
rect 10744 14968 10750 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 12342 14968 12348 15020
rect 12400 14968 12406 15020
rect 12820 15008 12848 15048
rect 14366 15036 14372 15088
rect 14424 15036 14430 15088
rect 14476 15076 14504 15116
rect 15010 15104 15016 15156
rect 15068 15144 15074 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15068 15116 15577 15144
rect 15068 15104 15074 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 15933 15147 15991 15153
rect 15933 15113 15945 15147
rect 15979 15144 15991 15147
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 15979 15116 18337 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 18782 15104 18788 15156
rect 18840 15104 18846 15156
rect 19242 15104 19248 15156
rect 19300 15144 19306 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 19300 15116 19533 15144
rect 19300 15104 19306 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 19521 15107 19579 15113
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22888 15116 22937 15144
rect 22888 15104 22894 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 22925 15107 22983 15113
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23808 15116 24133 15144
rect 23808 15104 23814 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 24121 15107 24179 15113
rect 25130 15104 25136 15156
rect 25188 15144 25194 15156
rect 25317 15147 25375 15153
rect 25317 15144 25329 15147
rect 25188 15116 25329 15144
rect 25188 15104 25194 15116
rect 25317 15113 25329 15116
rect 25363 15113 25375 15147
rect 25317 15107 25375 15113
rect 25593 15147 25651 15153
rect 25593 15113 25605 15147
rect 25639 15144 25651 15147
rect 25682 15144 25688 15156
rect 25639 15116 25688 15144
rect 25639 15113 25651 15116
rect 25593 15107 25651 15113
rect 25682 15104 25688 15116
rect 25740 15104 25746 15156
rect 26329 15147 26387 15153
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 27433 15147 27491 15153
rect 27433 15144 27445 15147
rect 26375 15116 27445 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 27433 15113 27445 15116
rect 27479 15144 27491 15147
rect 29733 15147 29791 15153
rect 27479 15116 29592 15144
rect 27479 15113 27491 15116
rect 27433 15107 27491 15113
rect 14476 15048 15240 15076
rect 12820 14980 13492 15008
rect 9585 14943 9643 14949
rect 9585 14909 9597 14943
rect 9631 14940 9643 14943
rect 9766 14940 9772 14952
rect 9631 14912 9772 14940
rect 9631 14909 9643 14912
rect 9585 14903 9643 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12360 14940 12388 14968
rect 11655 14912 12388 14940
rect 12437 14943 12495 14949
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 10137 14875 10195 14881
rect 10137 14841 10149 14875
rect 10183 14872 10195 14875
rect 11974 14872 11980 14884
rect 10183 14844 11980 14872
rect 10183 14841 10195 14844
rect 10137 14835 10195 14841
rect 11974 14832 11980 14844
rect 12032 14832 12038 14884
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 12452 14872 12480 14903
rect 12124 14844 12480 14872
rect 12124 14832 12130 14844
rect 10597 14807 10655 14813
rect 10597 14773 10609 14807
rect 10643 14804 10655 14807
rect 10686 14804 10692 14816
rect 10643 14776 10692 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 13464 14804 13492 14980
rect 15102 14968 15108 15020
rect 15160 14968 15166 15020
rect 15212 14952 15240 15048
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 16025 15079 16083 15085
rect 16025 15076 16037 15079
rect 15712 15048 16037 15076
rect 15712 15036 15718 15048
rect 16025 15045 16037 15048
rect 16071 15045 16083 15079
rect 18598 15076 18604 15088
rect 16025 15039 16083 15045
rect 17236 15048 18604 15076
rect 17236 15017 17264 15048
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20714 15076 20720 15088
rect 19935 15048 20720 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 21085 15079 21143 15085
rect 21085 15045 21097 15079
rect 21131 15076 21143 15079
rect 21818 15076 21824 15088
rect 21131 15048 21824 15076
rect 21131 15045 21143 15048
rect 21085 15039 21143 15045
rect 21818 15036 21824 15048
rect 21876 15036 21882 15088
rect 23385 15079 23443 15085
rect 23385 15045 23397 15079
rect 23431 15076 23443 15079
rect 25866 15076 25872 15088
rect 23431 15048 25872 15076
rect 23431 15045 23443 15048
rect 23385 15039 23443 15045
rect 25866 15036 25872 15048
rect 25924 15036 25930 15088
rect 27062 15036 27068 15088
rect 27120 15036 27126 15088
rect 28994 15036 29000 15088
rect 29052 15036 29058 15088
rect 29564 15076 29592 15116
rect 29733 15113 29745 15147
rect 29779 15144 29791 15147
rect 29822 15144 29828 15156
rect 29779 15116 29828 15144
rect 29779 15113 29791 15116
rect 29733 15107 29791 15113
rect 29822 15104 29828 15116
rect 29880 15104 29886 15156
rect 30466 15104 30472 15156
rect 30524 15144 30530 15156
rect 30561 15147 30619 15153
rect 30561 15144 30573 15147
rect 30524 15116 30573 15144
rect 30524 15104 30530 15116
rect 30561 15113 30573 15116
rect 30607 15113 30619 15147
rect 30561 15107 30619 15113
rect 31294 15104 31300 15156
rect 31352 15144 31358 15156
rect 31389 15147 31447 15153
rect 31389 15144 31401 15147
rect 31352 15116 31401 15144
rect 31352 15104 31358 15116
rect 31389 15113 31401 15116
rect 31435 15113 31447 15147
rect 31389 15107 31447 15113
rect 31496 15116 33088 15144
rect 31496 15076 31524 15116
rect 31849 15079 31907 15085
rect 31849 15076 31861 15079
rect 29564 15048 31524 15076
rect 31726 15048 31861 15076
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 14977 17279 15011
rect 17221 14971 17279 14977
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 15008 18751 15011
rect 19058 15008 19064 15020
rect 18739 14980 19064 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20898 15008 20904 15020
rect 20027 14980 20904 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21100 14980 22017 15008
rect 21100 14952 21128 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 23290 14968 23296 15020
rect 23348 14968 23354 15020
rect 24118 14968 24124 15020
rect 24176 15008 24182 15020
rect 24489 15011 24547 15017
rect 24489 15008 24501 15011
rect 24176 14980 24501 15008
rect 24176 14968 24182 14980
rect 24489 14977 24501 14980
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 24578 14968 24584 15020
rect 24636 15008 24642 15020
rect 25225 15011 25283 15017
rect 25225 15008 25237 15011
rect 24636 14980 25237 15008
rect 24636 14968 24642 14980
rect 25225 14977 25237 14980
rect 25271 15008 25283 15011
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 25271 14980 26249 15008
rect 25271 14977 25283 14980
rect 25225 14971 25283 14977
rect 26237 14977 26249 14980
rect 26283 15008 26295 15011
rect 27249 15011 27307 15017
rect 27249 15008 27261 15011
rect 26283 14980 27261 15008
rect 26283 14977 26295 14980
rect 26237 14971 26295 14977
rect 27249 14977 27261 14980
rect 27295 15008 27307 15011
rect 27338 15008 27344 15020
rect 27295 14980 27344 15008
rect 27295 14977 27307 14980
rect 27249 14971 27307 14977
rect 27338 14968 27344 14980
rect 27396 14968 27402 15020
rect 27798 14968 27804 15020
rect 27856 15008 27862 15020
rect 27985 15011 28043 15017
rect 27985 15008 27997 15011
rect 27856 14980 27997 15008
rect 27856 14968 27862 14980
rect 27985 14977 27997 14980
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 29546 14968 29552 15020
rect 29604 15008 29610 15020
rect 30653 15011 30711 15017
rect 30653 15008 30665 15011
rect 29604 14980 30665 15008
rect 29604 14968 29610 14980
rect 30653 14977 30665 14980
rect 30699 15008 30711 15011
rect 31726 15008 31754 15048
rect 31849 15045 31861 15048
rect 31895 15045 31907 15079
rect 33060 15076 33088 15116
rect 33870 15104 33876 15156
rect 33928 15104 33934 15156
rect 35069 15147 35127 15153
rect 35069 15113 35081 15147
rect 35115 15144 35127 15147
rect 37458 15144 37464 15156
rect 35115 15116 37464 15144
rect 35115 15113 35127 15116
rect 35069 15107 35127 15113
rect 37458 15104 37464 15116
rect 37516 15104 37522 15156
rect 39669 15147 39727 15153
rect 39669 15144 39681 15147
rect 37568 15116 39681 15144
rect 34054 15076 34060 15088
rect 33060 15048 34060 15076
rect 31849 15039 31907 15045
rect 34054 15036 34060 15048
rect 34112 15036 34118 15088
rect 35802 15036 35808 15088
rect 35860 15076 35866 15088
rect 36173 15079 36231 15085
rect 36173 15076 36185 15079
rect 35860 15048 36185 15076
rect 35860 15036 35866 15048
rect 36173 15045 36185 15048
rect 36219 15045 36231 15079
rect 36173 15039 36231 15045
rect 36265 15079 36323 15085
rect 36265 15045 36277 15079
rect 36311 15076 36323 15079
rect 36354 15076 36360 15088
rect 36311 15048 36360 15076
rect 36311 15045 36323 15048
rect 36265 15039 36323 15045
rect 36354 15036 36360 15048
rect 36412 15036 36418 15088
rect 37568 15076 37596 15116
rect 39669 15113 39681 15116
rect 39715 15113 39727 15147
rect 39669 15107 39727 15113
rect 39942 15104 39948 15156
rect 40000 15144 40006 15156
rect 40129 15147 40187 15153
rect 40129 15144 40141 15147
rect 40000 15116 40141 15144
rect 40000 15104 40006 15116
rect 40129 15113 40141 15116
rect 40175 15113 40187 15147
rect 40129 15107 40187 15113
rect 36556 15048 37596 15076
rect 32677 15011 32735 15017
rect 32677 15008 32689 15011
rect 30699 14980 31754 15008
rect 31864 14980 32689 15008
rect 30699 14977 30711 14980
rect 30653 14971 30711 14977
rect 31864 14952 31892 14980
rect 32677 14977 32689 14980
rect 32723 14977 32735 15011
rect 32677 14971 32735 14977
rect 32769 15011 32827 15017
rect 32769 14977 32781 15011
rect 32815 15008 32827 15011
rect 32815 14980 36216 15008
rect 32815 14977 32827 14980
rect 32769 14971 32827 14977
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 14274 14940 14280 14952
rect 13688 14912 14280 14940
rect 13688 14900 13694 14912
rect 14274 14900 14280 14912
rect 14332 14900 14338 14952
rect 14734 14900 14740 14952
rect 14792 14940 14798 14952
rect 14829 14943 14887 14949
rect 14829 14940 14841 14943
rect 14792 14912 14841 14940
rect 14792 14900 14798 14912
rect 14829 14909 14841 14912
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 15194 14900 15200 14952
rect 15252 14940 15258 14952
rect 16117 14943 16175 14949
rect 16117 14940 16129 14943
rect 15252 14912 16129 14940
rect 15252 14900 15258 14912
rect 16117 14909 16129 14912
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 15028 14844 16988 14872
rect 15028 14804 15056 14844
rect 13464 14776 15056 14804
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 16264 14776 16865 14804
rect 16264 14764 16270 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16960 14804 16988 14844
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 17328 14872 17356 14903
rect 17402 14900 17408 14952
rect 17460 14900 17466 14952
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 20990 14940 20996 14952
rect 20211 14912 20996 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 17276 14844 17356 14872
rect 17276 14832 17282 14844
rect 18046 14832 18052 14884
rect 18104 14832 18110 14884
rect 18892 14872 18920 14903
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 21082 14900 21088 14952
rect 21140 14900 21146 14952
rect 21177 14943 21235 14949
rect 21177 14909 21189 14943
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14940 21419 14943
rect 21542 14940 21548 14952
rect 21407 14912 21548 14940
rect 21407 14909 21419 14912
rect 21361 14903 21419 14909
rect 18966 14872 18972 14884
rect 18892 14844 18972 14872
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 19260 14844 20729 14872
rect 19260 14816 19288 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 21192 14872 21220 14903
rect 21542 14900 21548 14912
rect 21600 14900 21606 14952
rect 23569 14943 23627 14949
rect 23569 14909 23581 14943
rect 23615 14940 23627 14943
rect 24026 14940 24032 14952
rect 23615 14912 24032 14940
rect 23615 14909 23627 14912
rect 23569 14903 23627 14909
rect 24026 14900 24032 14912
rect 24084 14900 24090 14952
rect 24210 14900 24216 14952
rect 24268 14940 24274 14952
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 24268 14912 24685 14940
rect 24268 14900 24274 14912
rect 24673 14909 24685 14912
rect 24719 14909 24731 14943
rect 24673 14903 24731 14909
rect 26421 14943 26479 14949
rect 26421 14909 26433 14943
rect 26467 14909 26479 14943
rect 26421 14903 26479 14909
rect 28261 14943 28319 14949
rect 28261 14909 28273 14943
rect 28307 14940 28319 14943
rect 29730 14940 29736 14952
rect 28307 14912 29736 14940
rect 28307 14909 28319 14912
rect 28261 14903 28319 14909
rect 20717 14835 20775 14841
rect 21100 14844 21220 14872
rect 17770 14804 17776 14816
rect 16960 14776 17776 14804
rect 16853 14767 16911 14773
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 19242 14764 19248 14816
rect 19300 14764 19306 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 21100 14804 21128 14844
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 22796 14844 26004 14872
rect 22796 14832 22802 14844
rect 21726 14804 21732 14816
rect 20588 14776 21732 14804
rect 20588 14764 20594 14776
rect 21726 14764 21732 14776
rect 21784 14764 21790 14816
rect 22186 14764 22192 14816
rect 22244 14804 22250 14816
rect 24118 14804 24124 14816
rect 22244 14776 24124 14804
rect 22244 14764 22250 14776
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 25866 14764 25872 14816
rect 25924 14764 25930 14816
rect 25976 14804 26004 14844
rect 26142 14832 26148 14884
rect 26200 14872 26206 14884
rect 26436 14872 26464 14903
rect 29730 14900 29736 14912
rect 29788 14900 29794 14952
rect 29914 14900 29920 14952
rect 29972 14940 29978 14952
rect 30282 14940 30288 14952
rect 29972 14912 30288 14940
rect 29972 14900 29978 14912
rect 30282 14900 30288 14912
rect 30340 14940 30346 14952
rect 30745 14943 30803 14949
rect 30745 14940 30757 14943
rect 30340 14912 30757 14940
rect 30340 14900 30346 14912
rect 30745 14909 30757 14912
rect 30791 14909 30803 14943
rect 30745 14903 30803 14909
rect 31846 14900 31852 14952
rect 31904 14900 31910 14952
rect 32490 14900 32496 14952
rect 32548 14940 32554 14952
rect 32861 14943 32919 14949
rect 32861 14940 32873 14943
rect 32548 14912 32873 14940
rect 32548 14900 32554 14912
rect 32861 14909 32873 14912
rect 32907 14909 32919 14943
rect 32861 14903 32919 14909
rect 33042 14900 33048 14952
rect 33100 14940 33106 14952
rect 33410 14940 33416 14952
rect 33100 14912 33416 14940
rect 33100 14900 33106 14912
rect 33410 14900 33416 14912
rect 33468 14900 33474 14952
rect 33689 14943 33747 14949
rect 33689 14909 33701 14943
rect 33735 14909 33747 14943
rect 33689 14903 33747 14909
rect 26200 14844 26464 14872
rect 26200 14832 26206 14844
rect 29270 14832 29276 14884
rect 29328 14872 29334 14884
rect 32309 14875 32367 14881
rect 32309 14872 32321 14875
rect 29328 14844 32321 14872
rect 29328 14832 29334 14844
rect 32309 14841 32321 14844
rect 32355 14841 32367 14875
rect 33704 14872 33732 14903
rect 33778 14900 33784 14952
rect 33836 14900 33842 14952
rect 34885 14943 34943 14949
rect 34885 14909 34897 14943
rect 34931 14909 34943 14943
rect 34885 14903 34943 14909
rect 34977 14943 35035 14949
rect 34977 14909 34989 14943
rect 35023 14940 35035 14943
rect 36081 14943 36139 14949
rect 35023 14912 35940 14940
rect 35023 14909 35035 14912
rect 34977 14903 35035 14909
rect 33962 14872 33968 14884
rect 33704 14844 33968 14872
rect 32309 14835 32367 14841
rect 33962 14832 33968 14844
rect 34020 14832 34026 14884
rect 34606 14872 34612 14884
rect 34164 14844 34612 14872
rect 27525 14807 27583 14813
rect 27525 14804 27537 14807
rect 25976 14776 27537 14804
rect 27525 14773 27537 14776
rect 27571 14804 27583 14807
rect 28074 14804 28080 14816
rect 27571 14776 28080 14804
rect 27571 14773 27583 14776
rect 27525 14767 27583 14773
rect 28074 14764 28080 14776
rect 28132 14764 28138 14816
rect 28810 14764 28816 14816
rect 28868 14804 28874 14816
rect 29546 14804 29552 14816
rect 28868 14776 29552 14804
rect 28868 14764 28874 14776
rect 29546 14764 29552 14776
rect 29604 14764 29610 14816
rect 30190 14764 30196 14816
rect 30248 14764 30254 14816
rect 30466 14764 30472 14816
rect 30524 14804 30530 14816
rect 34164 14804 34192 14844
rect 34606 14832 34612 14844
rect 34664 14832 34670 14884
rect 34900 14872 34928 14903
rect 35342 14872 35348 14884
rect 34900 14844 35348 14872
rect 35342 14832 35348 14844
rect 35400 14832 35406 14884
rect 30524 14776 34192 14804
rect 30524 14764 30530 14776
rect 34238 14764 34244 14816
rect 34296 14764 34302 14816
rect 35434 14764 35440 14816
rect 35492 14764 35498 14816
rect 35912 14804 35940 14912
rect 36081 14909 36093 14943
rect 36127 14909 36139 14943
rect 36188 14940 36216 14980
rect 36556 14940 36584 15048
rect 37734 15036 37740 15088
rect 37792 15036 37798 15088
rect 38746 15036 38752 15088
rect 38804 15036 38810 15088
rect 40586 15036 40592 15088
rect 40644 15076 40650 15088
rect 40644 15048 40908 15076
rect 40644 15036 40650 15048
rect 37366 14968 37372 15020
rect 37424 15008 37430 15020
rect 40880 15017 40908 15048
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 37424 14980 37473 15008
rect 37424 14968 37430 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 40037 15011 40095 15017
rect 40037 14977 40049 15011
rect 40083 15008 40095 15011
rect 40865 15011 40923 15017
rect 40083 14980 40724 15008
rect 40083 14977 40095 14980
rect 40037 14971 40095 14977
rect 36188 14912 36584 14940
rect 36081 14903 36139 14909
rect 36096 14872 36124 14903
rect 38470 14900 38476 14952
rect 38528 14940 38534 14952
rect 39209 14943 39267 14949
rect 39209 14940 39221 14943
rect 38528 14912 39221 14940
rect 38528 14900 38534 14912
rect 39209 14909 39221 14912
rect 39255 14909 39267 14943
rect 39209 14903 39267 14909
rect 40218 14900 40224 14952
rect 40276 14900 40282 14952
rect 40696 14940 40724 14980
rect 40865 14977 40877 15011
rect 40911 14977 40923 15011
rect 40865 14971 40923 14977
rect 48225 15011 48283 15017
rect 48225 14977 48237 15011
rect 48271 15008 48283 15011
rect 48685 15011 48743 15017
rect 48685 15008 48697 15011
rect 48271 14980 48697 15008
rect 48271 14977 48283 14980
rect 48225 14971 48283 14977
rect 48685 14977 48697 14980
rect 48731 14977 48743 15011
rect 48685 14971 48743 14977
rect 49326 14968 49332 15020
rect 49384 14968 49390 15020
rect 46934 14940 46940 14952
rect 40696 14912 46940 14940
rect 46934 14900 46940 14912
rect 46992 14900 46998 14952
rect 47673 14943 47731 14949
rect 47673 14909 47685 14943
rect 47719 14940 47731 14943
rect 49344 14940 49372 14968
rect 47719 14912 49372 14940
rect 47719 14909 47731 14912
rect 47673 14903 47731 14909
rect 36538 14872 36544 14884
rect 36096 14844 36544 14872
rect 36538 14832 36544 14844
rect 36596 14832 36602 14884
rect 36633 14875 36691 14881
rect 36633 14841 36645 14875
rect 36679 14872 36691 14875
rect 36679 14844 37596 14872
rect 36679 14841 36691 14844
rect 36633 14835 36691 14841
rect 35986 14804 35992 14816
rect 35912 14776 35992 14804
rect 35986 14764 35992 14776
rect 36044 14804 36050 14816
rect 36909 14807 36967 14813
rect 36909 14804 36921 14807
rect 36044 14776 36921 14804
rect 36044 14764 36050 14776
rect 36909 14773 36921 14776
rect 36955 14773 36967 14807
rect 37568 14804 37596 14844
rect 48038 14832 48044 14884
rect 48096 14832 48102 14884
rect 38746 14804 38752 14816
rect 37568 14776 38752 14804
rect 36909 14767 36967 14773
rect 38746 14764 38752 14776
rect 38804 14764 38810 14816
rect 41049 14807 41107 14813
rect 41049 14773 41061 14807
rect 41095 14804 41107 14807
rect 45646 14804 45652 14816
rect 41095 14776 45652 14804
rect 41095 14773 41107 14776
rect 41049 14767 41107 14773
rect 45646 14764 45652 14776
rect 45704 14764 45710 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11480 14572 11805 14600
rect 11480 14560 11486 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12860 14572 13001 14600
rect 12860 14560 12866 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 14550 14600 14556 14612
rect 14507 14572 14556 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 17494 14560 17500 14612
rect 17552 14600 17558 14612
rect 18141 14603 18199 14609
rect 17552 14572 17632 14600
rect 17552 14560 17558 14572
rect 10226 14492 10232 14544
rect 10284 14492 10290 14544
rect 17604 14532 17632 14572
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18414 14600 18420 14612
rect 18187 14572 18420 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 21542 14560 21548 14612
rect 21600 14600 21606 14612
rect 22462 14600 22468 14612
rect 21600 14572 22468 14600
rect 21600 14560 21606 14572
rect 22462 14560 22468 14572
rect 22520 14600 22526 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 22520 14572 22845 14600
rect 22520 14560 22526 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 22833 14563 22891 14569
rect 25498 14560 25504 14612
rect 25556 14600 25562 14612
rect 25593 14603 25651 14609
rect 25593 14600 25605 14603
rect 25556 14572 25605 14600
rect 25556 14560 25562 14572
rect 25593 14569 25605 14572
rect 25639 14569 25651 14603
rect 25593 14563 25651 14569
rect 26418 14560 26424 14612
rect 26476 14600 26482 14612
rect 30558 14600 30564 14612
rect 26476 14572 30564 14600
rect 26476 14560 26482 14572
rect 30558 14560 30564 14572
rect 30616 14560 30622 14612
rect 31386 14560 31392 14612
rect 31444 14600 31450 14612
rect 33594 14600 33600 14612
rect 31444 14572 33600 14600
rect 31444 14560 31450 14572
rect 33594 14560 33600 14572
rect 33652 14560 33658 14612
rect 34238 14560 34244 14612
rect 34296 14600 34302 14612
rect 34296 14572 36216 14600
rect 34296 14560 34302 14572
rect 19242 14532 19248 14544
rect 14752 14504 17080 14532
rect 17604 14504 19248 14532
rect 934 14424 940 14476
rect 992 14464 998 14476
rect 1765 14467 1823 14473
rect 1765 14464 1777 14467
rect 992 14436 1777 14464
rect 992 14424 998 14436
rect 1765 14433 1777 14436
rect 1811 14433 1823 14467
rect 1765 14427 1823 14433
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 13262 14464 13268 14476
rect 12483 14436 13268 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 13504 14436 13553 14464
rect 13504 14424 13510 14436
rect 13541 14433 13553 14436
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 14185 14467 14243 14473
rect 14185 14433 14197 14467
rect 14231 14464 14243 14467
rect 14752 14464 14780 14504
rect 15120 14473 15148 14504
rect 17052 14476 17080 14504
rect 19242 14492 19248 14504
rect 19300 14492 19306 14544
rect 20162 14492 20168 14544
rect 20220 14532 20226 14544
rect 20717 14535 20775 14541
rect 20717 14532 20729 14535
rect 20220 14504 20729 14532
rect 20220 14492 20226 14504
rect 20717 14501 20729 14504
rect 20763 14501 20775 14535
rect 20717 14495 20775 14501
rect 14231 14436 14780 14464
rect 15105 14467 15163 14473
rect 14231 14433 14243 14436
rect 14185 14427 14243 14433
rect 15105 14433 15117 14467
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 15252 14436 16957 14464
rect 15252 14424 15258 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 17092 14436 17509 14464
rect 17092 14424 17098 14436
rect 17497 14433 17509 14436
rect 17543 14464 17555 14467
rect 18693 14467 18751 14473
rect 18693 14464 18705 14467
rect 17543 14436 18705 14464
rect 17543 14433 17555 14436
rect 17497 14427 17555 14433
rect 18693 14433 18705 14436
rect 18739 14433 18751 14467
rect 18693 14427 18751 14433
rect 20070 14424 20076 14476
rect 20128 14424 20134 14476
rect 20622 14424 20628 14476
rect 20680 14424 20686 14476
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 3007 14368 9505 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14332 14368 14841 14396
rect 14332 14356 14338 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 17460 14368 17601 14396
rect 17460 14356 17466 14368
rect 17589 14365 17601 14368
rect 17635 14365 17647 14399
rect 17589 14359 17647 14365
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 18414 14396 18420 14408
rect 18104 14368 18420 14396
rect 18104 14356 18110 14368
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 18782 14396 18788 14408
rect 18555 14368 18788 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 19889 14399 19947 14405
rect 19889 14396 19901 14399
rect 19668 14368 19901 14396
rect 19668 14356 19674 14368
rect 19889 14365 19901 14368
rect 19935 14396 19947 14399
rect 20640 14396 20668 14424
rect 19935 14368 20668 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14328 9735 14331
rect 9950 14328 9956 14340
rect 9723 14300 9956 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 9950 14288 9956 14300
rect 10008 14288 10014 14340
rect 10410 14288 10416 14340
rect 10468 14288 10474 14340
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12802 14328 12808 14340
rect 12207 14300 12808 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 12802 14288 12808 14300
rect 12860 14288 12866 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 15933 14331 15991 14337
rect 13403 14300 15056 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10560 14232 11161 14260
rect 10560 14220 10566 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 12710 14260 12716 14272
rect 12299 14232 12716 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 13906 14260 13912 14272
rect 13495 14232 13912 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13906 14220 13912 14232
rect 13964 14220 13970 14272
rect 14918 14220 14924 14272
rect 14976 14220 14982 14272
rect 15028 14260 15056 14300
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16761 14331 16819 14337
rect 16761 14328 16773 14331
rect 15979 14300 16773 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16761 14297 16773 14300
rect 16807 14297 16819 14331
rect 16761 14291 16819 14297
rect 16868 14300 18460 14328
rect 16868 14272 16896 14300
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15028 14232 16405 14260
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 16850 14220 16856 14272
rect 16908 14220 16914 14272
rect 17862 14220 17868 14272
rect 17920 14220 17926 14272
rect 18432 14260 18460 14300
rect 19794 14288 19800 14340
rect 19852 14328 19858 14340
rect 20530 14328 20536 14340
rect 19852 14300 20536 14328
rect 19852 14288 19858 14300
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 20732 14328 20760 14495
rect 22554 14492 22560 14544
rect 22612 14532 22618 14544
rect 25038 14532 25044 14544
rect 22612 14504 25044 14532
rect 22612 14492 22618 14504
rect 25038 14492 25044 14504
rect 25096 14492 25102 14544
rect 28534 14532 28540 14544
rect 27908 14504 28540 14532
rect 21082 14424 21088 14476
rect 21140 14424 21146 14476
rect 21358 14424 21364 14476
rect 21416 14424 21422 14476
rect 21726 14424 21732 14476
rect 21784 14464 21790 14476
rect 25774 14464 25780 14476
rect 21784 14436 25780 14464
rect 21784 14424 21790 14436
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 26050 14424 26056 14476
rect 26108 14464 26114 14476
rect 27065 14467 27123 14473
rect 27065 14464 27077 14467
rect 26108 14436 27077 14464
rect 26108 14424 26114 14436
rect 27065 14433 27077 14436
rect 27111 14464 27123 14467
rect 27798 14464 27804 14476
rect 27111 14436 27804 14464
rect 27111 14433 27123 14436
rect 27065 14427 27123 14433
rect 27798 14424 27804 14436
rect 27856 14424 27862 14476
rect 27908 14473 27936 14504
rect 28534 14492 28540 14504
rect 28592 14492 28598 14544
rect 30469 14535 30527 14541
rect 30469 14501 30481 14535
rect 30515 14532 30527 14535
rect 33778 14532 33784 14544
rect 30515 14504 33784 14532
rect 30515 14501 30527 14504
rect 30469 14495 30527 14501
rect 33778 14492 33784 14504
rect 33836 14492 33842 14544
rect 34057 14535 34115 14541
rect 34057 14501 34069 14535
rect 34103 14532 34115 14535
rect 36188 14532 36216 14572
rect 36630 14560 36636 14612
rect 36688 14560 36694 14612
rect 38378 14600 38384 14612
rect 36740 14572 38384 14600
rect 36740 14532 36768 14572
rect 38378 14560 38384 14572
rect 38436 14560 38442 14612
rect 38470 14560 38476 14612
rect 38528 14600 38534 14612
rect 38577 14603 38635 14609
rect 38577 14600 38589 14603
rect 38528 14572 38589 14600
rect 38528 14560 38534 14572
rect 38577 14569 38589 14572
rect 38623 14569 38635 14603
rect 38577 14563 38635 14569
rect 38838 14560 38844 14612
rect 38896 14600 38902 14612
rect 39853 14603 39911 14609
rect 39853 14600 39865 14603
rect 38896 14572 39865 14600
rect 38896 14560 38902 14572
rect 39853 14569 39865 14572
rect 39899 14600 39911 14603
rect 40037 14603 40095 14609
rect 40037 14600 40049 14603
rect 39899 14572 40049 14600
rect 39899 14569 39911 14572
rect 39853 14563 39911 14569
rect 40037 14569 40049 14572
rect 40083 14569 40095 14603
rect 40037 14563 40095 14569
rect 34103 14504 35020 14532
rect 36188 14504 36768 14532
rect 34103 14501 34115 14504
rect 34057 14495 34115 14501
rect 27893 14467 27951 14473
rect 27893 14433 27905 14467
rect 27939 14433 27951 14467
rect 29270 14464 29276 14476
rect 27893 14427 27951 14433
rect 28000 14436 29276 14464
rect 22830 14356 22836 14408
rect 22888 14396 22894 14408
rect 23477 14399 23535 14405
rect 23477 14396 23489 14399
rect 22888 14368 23489 14396
rect 22888 14356 22894 14368
rect 23477 14365 23489 14368
rect 23523 14365 23535 14399
rect 23477 14359 23535 14365
rect 24673 14399 24731 14405
rect 24673 14365 24685 14399
rect 24719 14396 24731 14399
rect 24719 14368 25728 14396
rect 24719 14365 24731 14368
rect 24673 14359 24731 14365
rect 25700 14340 25728 14368
rect 27338 14356 27344 14408
rect 27396 14356 27402 14408
rect 28000 14396 28028 14436
rect 29270 14424 29276 14436
rect 29328 14464 29334 14476
rect 29638 14464 29644 14476
rect 29328 14436 29644 14464
rect 29328 14424 29334 14436
rect 29638 14424 29644 14436
rect 29696 14424 29702 14476
rect 29917 14467 29975 14473
rect 29917 14433 29929 14467
rect 29963 14464 29975 14467
rect 30650 14464 30656 14476
rect 29963 14436 30656 14464
rect 29963 14433 29975 14436
rect 29917 14427 29975 14433
rect 30650 14424 30656 14436
rect 30708 14424 30714 14476
rect 30834 14424 30840 14476
rect 30892 14464 30898 14476
rect 31021 14467 31079 14473
rect 31021 14464 31033 14467
rect 30892 14436 31033 14464
rect 30892 14424 30898 14436
rect 31021 14433 31033 14436
rect 31067 14433 31079 14467
rect 31021 14427 31079 14433
rect 31202 14424 31208 14476
rect 31260 14464 31266 14476
rect 31478 14464 31484 14476
rect 31260 14436 31484 14464
rect 31260 14424 31266 14436
rect 31478 14424 31484 14436
rect 31536 14464 31542 14476
rect 32217 14467 32275 14473
rect 32217 14464 32229 14467
rect 31536 14436 32229 14464
rect 31536 14424 31542 14436
rect 32217 14433 32229 14436
rect 32263 14433 32275 14467
rect 32217 14427 32275 14433
rect 32306 14424 32312 14476
rect 32364 14464 32370 14476
rect 33413 14467 33471 14473
rect 33413 14464 33425 14467
rect 32364 14436 33425 14464
rect 32364 14424 32370 14436
rect 33413 14433 33425 14436
rect 33459 14433 33471 14467
rect 33413 14427 33471 14433
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 34885 14467 34943 14473
rect 34885 14464 34897 14467
rect 34848 14436 34897 14464
rect 34848 14424 34854 14436
rect 34885 14433 34897 14436
rect 34931 14433 34943 14467
rect 34992 14464 35020 14504
rect 37090 14464 37096 14476
rect 34992 14436 37096 14464
rect 34885 14427 34943 14433
rect 37090 14424 37096 14436
rect 37148 14424 37154 14476
rect 37366 14424 37372 14476
rect 37424 14464 37430 14476
rect 38841 14467 38899 14473
rect 38841 14464 38853 14467
rect 37424 14436 38853 14464
rect 37424 14424 37430 14436
rect 38841 14433 38853 14436
rect 38887 14433 38899 14467
rect 38841 14427 38899 14433
rect 47673 14467 47731 14473
rect 47673 14433 47685 14467
rect 47719 14464 47731 14467
rect 47719 14436 49372 14464
rect 47719 14433 47731 14436
rect 47673 14427 47731 14433
rect 49344 14408 49372 14436
rect 27448 14368 28028 14396
rect 21634 14328 21640 14340
rect 20732 14300 21640 14328
rect 21634 14288 21640 14300
rect 21692 14328 21698 14340
rect 21692 14300 21850 14328
rect 22664 14300 25268 14328
rect 21692 14288 21698 14300
rect 18506 14260 18512 14272
rect 18432 14232 18512 14260
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 18598 14220 18604 14272
rect 18656 14220 18662 14272
rect 19518 14220 19524 14272
rect 19576 14220 19582 14272
rect 19702 14220 19708 14272
rect 19760 14260 19766 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19760 14232 19993 14260
rect 19760 14220 19766 14232
rect 19981 14229 19993 14232
rect 20027 14260 20039 14263
rect 22664 14260 22692 14300
rect 20027 14232 22692 14260
rect 20027 14229 20039 14232
rect 19981 14223 20039 14229
rect 23198 14220 23204 14272
rect 23256 14220 23262 14272
rect 23842 14220 23848 14272
rect 23900 14220 23906 14272
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 25130 14220 25136 14272
rect 25188 14220 25194 14272
rect 25240 14260 25268 14300
rect 25682 14288 25688 14340
rect 25740 14328 25746 14340
rect 25740 14300 25898 14328
rect 25740 14288 25746 14300
rect 27448 14260 27476 14368
rect 28074 14356 28080 14408
rect 28132 14396 28138 14408
rect 28626 14396 28632 14408
rect 28132 14368 28632 14396
rect 28132 14356 28138 14368
rect 28626 14356 28632 14368
rect 28684 14356 28690 14408
rect 30006 14356 30012 14408
rect 30064 14396 30070 14408
rect 31297 14399 31355 14405
rect 31297 14396 31309 14399
rect 30064 14368 31309 14396
rect 30064 14356 30070 14368
rect 31297 14365 31309 14368
rect 31343 14365 31355 14399
rect 32401 14399 32459 14405
rect 32401 14396 32413 14399
rect 31297 14359 31355 14365
rect 31404 14368 32413 14396
rect 27706 14288 27712 14340
rect 27764 14328 27770 14340
rect 28169 14331 28227 14337
rect 28169 14328 28181 14331
rect 27764 14300 28181 14328
rect 27764 14288 27770 14300
rect 28169 14297 28181 14300
rect 28215 14297 28227 14331
rect 31205 14331 31263 14337
rect 31205 14328 31217 14331
rect 28169 14291 28227 14297
rect 28552 14300 31217 14328
rect 28552 14269 28580 14300
rect 31205 14297 31217 14300
rect 31251 14297 31263 14331
rect 31205 14291 31263 14297
rect 25240 14232 27476 14260
rect 28537 14263 28595 14269
rect 28537 14229 28549 14263
rect 28583 14229 28595 14263
rect 28537 14223 28595 14229
rect 28994 14220 29000 14272
rect 29052 14220 29058 14272
rect 29362 14220 29368 14272
rect 29420 14260 29426 14272
rect 30009 14263 30067 14269
rect 30009 14260 30021 14263
rect 29420 14232 30021 14260
rect 29420 14220 29426 14232
rect 30009 14229 30021 14232
rect 30055 14229 30067 14263
rect 30009 14223 30067 14229
rect 30098 14220 30104 14272
rect 30156 14220 30162 14272
rect 30558 14220 30564 14272
rect 30616 14260 30622 14272
rect 31404 14260 31432 14368
rect 32401 14365 32413 14368
rect 32447 14365 32459 14399
rect 32401 14359 32459 14365
rect 32858 14356 32864 14408
rect 32916 14396 32922 14408
rect 33597 14399 33655 14405
rect 33597 14396 33609 14399
rect 32916 14368 33609 14396
rect 32916 14356 32922 14368
rect 33597 14365 33609 14368
rect 33643 14365 33655 14399
rect 33597 14359 33655 14365
rect 33686 14356 33692 14408
rect 33744 14356 33750 14408
rect 39298 14356 39304 14408
rect 39356 14356 39362 14408
rect 47946 14356 47952 14408
rect 48004 14356 48010 14408
rect 49326 14356 49332 14408
rect 49384 14356 49390 14408
rect 33318 14328 33324 14340
rect 31680 14300 33324 14328
rect 31680 14269 31708 14300
rect 33318 14288 33324 14300
rect 33376 14288 33382 14340
rect 34790 14288 34796 14340
rect 34848 14328 34854 14340
rect 35158 14328 35164 14340
rect 34848 14300 35164 14328
rect 34848 14288 34854 14300
rect 35158 14288 35164 14300
rect 35216 14288 35222 14340
rect 36446 14328 36452 14340
rect 36386 14300 36452 14328
rect 36446 14288 36452 14300
rect 36504 14288 36510 14340
rect 38838 14328 38844 14340
rect 38134 14300 38844 14328
rect 38838 14288 38844 14300
rect 38896 14288 38902 14340
rect 48133 14331 48191 14337
rect 48133 14297 48145 14331
rect 48179 14328 48191 14331
rect 48685 14331 48743 14337
rect 48685 14328 48697 14331
rect 48179 14300 48697 14328
rect 48179 14297 48191 14300
rect 48133 14291 48191 14297
rect 48685 14297 48697 14300
rect 48731 14297 48743 14331
rect 48685 14291 48743 14297
rect 30616 14232 31432 14260
rect 31665 14263 31723 14269
rect 30616 14220 30622 14232
rect 31665 14229 31677 14263
rect 31711 14229 31723 14263
rect 31665 14223 31723 14229
rect 32493 14263 32551 14269
rect 32493 14229 32505 14263
rect 32539 14260 32551 14263
rect 32582 14260 32588 14272
rect 32539 14232 32588 14260
rect 32539 14229 32551 14232
rect 32493 14223 32551 14229
rect 32582 14220 32588 14232
rect 32640 14220 32646 14272
rect 32766 14220 32772 14272
rect 32824 14260 32830 14272
rect 32861 14263 32919 14269
rect 32861 14260 32873 14263
rect 32824 14232 32873 14260
rect 32824 14220 32830 14232
rect 32861 14229 32873 14232
rect 32907 14229 32919 14263
rect 32861 14223 32919 14229
rect 33410 14220 33416 14272
rect 33468 14260 33474 14272
rect 34238 14260 34244 14272
rect 33468 14232 34244 14260
rect 33468 14220 33474 14232
rect 34238 14220 34244 14232
rect 34296 14260 34302 14272
rect 34333 14263 34391 14269
rect 34333 14260 34345 14263
rect 34296 14232 34345 14260
rect 34296 14220 34302 14232
rect 34333 14229 34345 14232
rect 34379 14229 34391 14263
rect 34333 14223 34391 14229
rect 35434 14220 35440 14272
rect 35492 14260 35498 14272
rect 36814 14260 36820 14272
rect 35492 14232 36820 14260
rect 35492 14220 35498 14232
rect 36814 14220 36820 14232
rect 36872 14220 36878 14272
rect 37093 14263 37151 14269
rect 37093 14229 37105 14263
rect 37139 14260 37151 14263
rect 37182 14260 37188 14272
rect 37139 14232 37188 14260
rect 37139 14229 37151 14232
rect 37093 14223 37151 14229
rect 37182 14220 37188 14232
rect 37240 14220 37246 14272
rect 37550 14220 37556 14272
rect 37608 14260 37614 14272
rect 38470 14260 38476 14272
rect 37608 14232 38476 14260
rect 37608 14220 37614 14232
rect 38470 14220 38476 14232
rect 38528 14220 38534 14272
rect 39482 14220 39488 14272
rect 39540 14220 39546 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 9858 14056 9864 14068
rect 3651 14028 9864 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 9950 14016 9956 14068
rect 10008 14016 10014 14068
rect 10689 14059 10747 14065
rect 10689 14025 10701 14059
rect 10735 14056 10747 14059
rect 11238 14056 11244 14068
rect 10735 14028 11244 14056
rect 10735 14025 10747 14028
rect 10689 14019 10747 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11940 14028 11989 14056
rect 11940 14016 11946 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 14332 14028 15577 14056
rect 14332 14016 14338 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 16758 14056 16764 14068
rect 15712 14028 16764 14056
rect 15712 14016 15718 14028
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 16850 14016 16856 14068
rect 16908 14056 16914 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 16908 14028 17141 14056
rect 16908 14016 16914 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17129 14019 17187 14025
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19426 14056 19432 14068
rect 18739 14028 19432 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 20162 14016 20168 14068
rect 20220 14016 20226 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21416 14028 21465 14056
rect 21416 14016 21422 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 22005 14059 22063 14065
rect 22005 14025 22017 14059
rect 22051 14056 22063 14059
rect 22094 14056 22100 14068
rect 22051 14028 22100 14056
rect 22051 14025 22063 14028
rect 22005 14019 22063 14025
rect 22094 14016 22100 14028
rect 22152 14016 22158 14068
rect 23198 14056 23204 14068
rect 22388 14028 23204 14056
rect 1026 13948 1032 14000
rect 1084 13988 1090 14000
rect 1765 13991 1823 13997
rect 1765 13988 1777 13991
rect 1084 13960 1777 13988
rect 1084 13948 1090 13960
rect 1765 13957 1777 13960
rect 1811 13957 1823 13991
rect 10502 13988 10508 14000
rect 1765 13951 1823 13957
rect 2976 13960 10508 13988
rect 2976 13929 3004 13960
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 13262 13948 13268 14000
rect 13320 13948 13326 14000
rect 15010 13988 15016 14000
rect 14490 13960 15016 13988
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 16025 13991 16083 13997
rect 16025 13957 16037 13991
rect 16071 13988 16083 13991
rect 19518 13988 19524 14000
rect 16071 13960 19524 13988
rect 16071 13957 16083 13960
rect 16025 13951 16083 13957
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 20180 13988 20208 14016
rect 22186 13988 22192 14000
rect 20180 13960 20470 13988
rect 21284 13960 22192 13988
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3568 13892 3985 13920
rect 3568 13880 3574 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11195 13892 12081 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 14642 13880 14648 13932
rect 14700 13920 14706 13932
rect 15197 13923 15255 13929
rect 15197 13920 15209 13923
rect 14700 13892 15209 13920
rect 14700 13880 14706 13892
rect 15197 13889 15209 13892
rect 15243 13889 15255 13923
rect 15197 13883 15255 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16206 13920 16212 13932
rect 15979 13892 16212 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 18598 13920 18604 13932
rect 16816 13892 18604 13920
rect 16816 13880 16822 13892
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 19429 13923 19487 13929
rect 19429 13889 19441 13923
rect 19475 13920 19487 13923
rect 19610 13920 19616 13932
rect 19475 13892 19616 13920
rect 19475 13889 19487 13892
rect 19429 13883 19487 13889
rect 19610 13880 19616 13892
rect 19668 13880 19674 13932
rect 10502 13812 10508 13864
rect 10560 13812 10566 13864
rect 11885 13855 11943 13861
rect 11885 13852 11897 13855
rect 10612 13824 11897 13852
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10612 13784 10640 13824
rect 11885 13821 11897 13824
rect 11931 13852 11943 13855
rect 12526 13852 12532 13864
rect 11931 13824 12532 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13852 13047 13855
rect 16117 13855 16175 13861
rect 13035 13824 13124 13852
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 9824 13756 10640 13784
rect 9824 13744 9830 13756
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 13096 13784 13124 13824
rect 16117 13821 16129 13855
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 10836 13756 13124 13784
rect 10836 13744 10842 13756
rect 12066 13676 12072 13728
rect 12124 13716 12130 13728
rect 12437 13719 12495 13725
rect 12437 13716 12449 13719
rect 12124 13688 12449 13716
rect 12124 13676 12130 13688
rect 12437 13685 12449 13688
rect 12483 13685 12495 13719
rect 13096 13716 13124 13756
rect 14458 13744 14464 13796
rect 14516 13784 14522 13796
rect 16132 13784 16160 13815
rect 17034 13812 17040 13864
rect 17092 13852 17098 13864
rect 17494 13852 17500 13864
rect 17092 13824 17500 13852
rect 17092 13812 17098 13824
rect 17494 13812 17500 13824
rect 17552 13812 17558 13864
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 14516 13756 16160 13784
rect 14516 13744 14522 13756
rect 16298 13744 16304 13796
rect 16356 13784 16362 13796
rect 17788 13784 17816 13815
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 17920 13824 18797 13852
rect 17920 13812 17926 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 17954 13784 17960 13796
rect 16356 13756 17724 13784
rect 17788 13756 17960 13784
rect 16356 13744 16362 13756
rect 13630 13716 13636 13728
rect 13096 13688 13636 13716
rect 12437 13679 12495 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 14737 13719 14795 13725
rect 14737 13685 14749 13719
rect 14783 13716 14795 13719
rect 16022 13716 16028 13728
rect 14783 13688 16028 13716
rect 14783 13685 14795 13688
rect 14737 13679 14795 13685
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 16114 13676 16120 13728
rect 16172 13716 16178 13728
rect 17402 13716 17408 13728
rect 16172 13688 17408 13716
rect 16172 13676 16178 13688
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17696 13716 17724 13756
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 18800 13784 18828 13815
rect 18874 13812 18880 13864
rect 18932 13812 18938 13864
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19024 13824 19717 13852
rect 19024 13812 19030 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 21284 13852 21312 13960
rect 22186 13948 22192 13960
rect 22244 13948 22250 14000
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 22388 13920 22416 14028
rect 23198 14016 23204 14028
rect 23256 14016 23262 14068
rect 24857 14059 24915 14065
rect 24857 14025 24869 14059
rect 24903 14056 24915 14059
rect 25314 14056 25320 14068
rect 24903 14028 25320 14056
rect 24903 14025 24915 14028
rect 24857 14019 24915 14025
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 25556 14028 26004 14056
rect 25556 14016 25562 14028
rect 25682 13948 25688 14000
rect 25740 13948 25746 14000
rect 25976 13988 26004 14028
rect 26510 14016 26516 14068
rect 26568 14016 26574 14068
rect 27614 14016 27620 14068
rect 27672 14016 27678 14068
rect 27798 14016 27804 14068
rect 27856 14056 27862 14068
rect 29365 14059 29423 14065
rect 29365 14056 29377 14059
rect 27856 14028 29377 14056
rect 27856 14016 27862 14028
rect 29365 14025 29377 14028
rect 29411 14025 29423 14059
rect 29365 14019 29423 14025
rect 30006 14016 30012 14068
rect 30064 14056 30070 14068
rect 31110 14056 31116 14068
rect 30064 14028 31116 14056
rect 30064 14016 30070 14028
rect 31110 14016 31116 14028
rect 31168 14016 31174 14068
rect 31757 14059 31815 14065
rect 31757 14025 31769 14059
rect 31803 14056 31815 14059
rect 36081 14059 36139 14065
rect 36081 14056 36093 14059
rect 31803 14028 36093 14056
rect 31803 14025 31815 14028
rect 31757 14019 31815 14025
rect 36081 14025 36093 14028
rect 36127 14025 36139 14059
rect 36081 14019 36139 14025
rect 36449 14059 36507 14065
rect 36449 14025 36461 14059
rect 36495 14056 36507 14059
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 36495 14028 37841 14056
rect 36495 14025 36507 14028
rect 36449 14019 36507 14025
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 37829 14019 37887 14025
rect 38197 14059 38255 14065
rect 38197 14025 38209 14059
rect 38243 14056 38255 14059
rect 41322 14056 41328 14068
rect 38243 14028 41328 14056
rect 38243 14025 38255 14028
rect 38197 14019 38255 14025
rect 41322 14016 41328 14028
rect 41380 14016 41386 14068
rect 45833 14059 45891 14065
rect 45833 14025 45845 14059
rect 45879 14056 45891 14059
rect 47210 14056 47216 14068
rect 45879 14028 47216 14056
rect 45879 14025 45891 14028
rect 45833 14019 45891 14025
rect 47210 14016 47216 14028
rect 47268 14016 47274 14068
rect 26329 13991 26387 13997
rect 26329 13988 26341 13991
rect 25976 13960 26341 13988
rect 26329 13957 26341 13960
rect 26375 13957 26387 13991
rect 26528 13988 26556 14016
rect 28810 13988 28816 14000
rect 26528 13960 28816 13988
rect 26329 13951 26387 13957
rect 28810 13948 28816 13960
rect 28868 13948 28874 14000
rect 30406 13960 31524 13988
rect 31496 13932 31524 13960
rect 34698 13948 34704 14000
rect 34756 13988 34762 14000
rect 34793 13991 34851 13997
rect 34793 13988 34805 13991
rect 34756 13960 34805 13988
rect 34756 13948 34762 13960
rect 34793 13957 34805 13960
rect 34839 13957 34851 13991
rect 34793 13951 34851 13957
rect 34882 13948 34888 14000
rect 34940 13948 34946 14000
rect 35158 13948 35164 14000
rect 35216 13988 35222 14000
rect 36909 13991 36967 13997
rect 36909 13988 36921 13991
rect 35216 13960 36921 13988
rect 35216 13948 35222 13960
rect 36909 13957 36921 13960
rect 36955 13988 36967 13991
rect 36998 13988 37004 14000
rect 36955 13960 37004 13988
rect 36955 13957 36967 13960
rect 36909 13951 36967 13957
rect 36998 13948 37004 13960
rect 37056 13948 37062 14000
rect 37274 13948 37280 14000
rect 37332 13988 37338 14000
rect 37737 13991 37795 13997
rect 37737 13988 37749 13991
rect 37332 13960 37749 13988
rect 37332 13948 37338 13960
rect 37737 13957 37749 13960
rect 37783 13957 37795 13991
rect 37737 13951 37795 13957
rect 38565 13991 38623 13997
rect 38565 13957 38577 13991
rect 38611 13988 38623 13991
rect 38838 13988 38844 14000
rect 38611 13960 38844 13988
rect 38611 13957 38623 13960
rect 38565 13951 38623 13957
rect 38838 13948 38844 13960
rect 38896 13988 38902 14000
rect 38933 13991 38991 13997
rect 38933 13988 38945 13991
rect 38896 13960 38945 13988
rect 38896 13948 38902 13960
rect 38933 13957 38945 13960
rect 38979 13957 38991 13991
rect 38933 13951 38991 13957
rect 39482 13948 39488 14000
rect 39540 13988 39546 14000
rect 45005 13991 45063 13997
rect 45005 13988 45017 13991
rect 39540 13960 45017 13988
rect 39540 13948 39546 13960
rect 45005 13957 45017 13960
rect 45051 13957 45063 13991
rect 45005 13951 45063 13957
rect 47854 13948 47860 14000
rect 47912 13988 47918 14000
rect 47949 13991 48007 13997
rect 47949 13988 47961 13991
rect 47912 13960 47961 13988
rect 47912 13948 47918 13960
rect 47949 13957 47961 13960
rect 47995 13957 48007 13991
rect 47949 13951 48007 13957
rect 21692 13906 22416 13920
rect 23753 13923 23811 13929
rect 21692 13892 22402 13906
rect 21692 13880 21698 13892
rect 23753 13889 23765 13923
rect 23799 13920 23811 13923
rect 24486 13920 24492 13932
rect 23799 13892 24492 13920
rect 23799 13889 23811 13892
rect 23753 13883 23811 13889
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 28902 13880 28908 13932
rect 28960 13880 28966 13932
rect 31110 13880 31116 13932
rect 31168 13880 31174 13932
rect 31478 13880 31484 13932
rect 31536 13920 31542 13932
rect 31754 13920 31760 13932
rect 31536 13892 31760 13920
rect 31536 13880 31542 13892
rect 31754 13880 31760 13892
rect 31812 13920 31818 13932
rect 31812 13892 32706 13920
rect 31812 13880 31818 13892
rect 35250 13880 35256 13932
rect 35308 13880 35314 13932
rect 35618 13880 35624 13932
rect 35676 13920 35682 13932
rect 35989 13923 36047 13929
rect 35989 13920 36001 13923
rect 35676 13892 36001 13920
rect 35676 13880 35682 13892
rect 35989 13889 36001 13892
rect 36035 13889 36047 13923
rect 35989 13883 36047 13889
rect 36170 13880 36176 13932
rect 36228 13920 36234 13932
rect 37182 13920 37188 13932
rect 36228 13892 37188 13920
rect 36228 13880 36234 13892
rect 37182 13880 37188 13892
rect 37240 13920 37246 13932
rect 40218 13920 40224 13932
rect 37240 13892 40224 13920
rect 37240 13880 37246 13892
rect 40218 13880 40224 13892
rect 40276 13880 40282 13932
rect 45646 13880 45652 13932
rect 45704 13880 45710 13932
rect 47213 13923 47271 13929
rect 47213 13889 47225 13923
rect 47259 13889 47271 13923
rect 47213 13883 47271 13889
rect 48133 13923 48191 13929
rect 48133 13889 48145 13923
rect 48179 13920 48191 13923
rect 48685 13923 48743 13929
rect 48685 13920 48697 13923
rect 48179 13892 48697 13920
rect 48179 13889 48191 13892
rect 48133 13883 48191 13889
rect 48685 13889 48697 13892
rect 48731 13889 48743 13923
rect 48685 13883 48743 13889
rect 19705 13815 19763 13821
rect 19812 13824 21312 13852
rect 19812 13784 19840 13824
rect 21910 13812 21916 13864
rect 21968 13852 21974 13864
rect 23477 13855 23535 13861
rect 23477 13852 23489 13855
rect 21968 13824 23489 13852
rect 21968 13812 21974 13824
rect 23477 13821 23489 13824
rect 23523 13852 23535 13855
rect 23523 13824 23704 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 22002 13784 22008 13796
rect 18800 13756 19840 13784
rect 21008 13756 22008 13784
rect 19702 13716 19708 13728
rect 17696 13688 19708 13716
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 19978 13725 19984 13728
rect 19968 13719 19984 13725
rect 19968 13685 19980 13719
rect 20036 13716 20042 13728
rect 21008 13716 21036 13756
rect 22002 13744 22008 13756
rect 22060 13744 22066 13796
rect 23676 13784 23704 13824
rect 23934 13812 23940 13864
rect 23992 13852 23998 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23992 13824 24225 13852
rect 23992 13812 23998 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 26605 13855 26663 13861
rect 26605 13821 26617 13855
rect 26651 13852 26663 13855
rect 27338 13852 27344 13864
rect 26651 13824 27344 13852
rect 26651 13821 26663 13824
rect 26605 13815 26663 13821
rect 27338 13812 27344 13824
rect 27396 13812 27402 13864
rect 30837 13855 30895 13861
rect 30837 13821 30849 13855
rect 30883 13852 30895 13855
rect 32309 13855 32367 13861
rect 32309 13852 32321 13855
rect 30883 13824 31064 13852
rect 30883 13821 30895 13824
rect 30837 13815 30895 13821
rect 24302 13784 24308 13796
rect 23676 13756 24308 13784
rect 24302 13744 24308 13756
rect 24360 13744 24366 13796
rect 28442 13744 28448 13796
rect 28500 13784 28506 13796
rect 29086 13784 29092 13796
rect 28500 13756 29092 13784
rect 28500 13744 28506 13756
rect 29086 13744 29092 13756
rect 29144 13744 29150 13796
rect 31036 13784 31064 13824
rect 31726 13824 32321 13852
rect 31726 13784 31754 13824
rect 32309 13821 32321 13824
rect 32355 13852 32367 13855
rect 32490 13852 32496 13864
rect 32355 13824 32496 13852
rect 32355 13821 32367 13824
rect 32309 13815 32367 13821
rect 32490 13812 32496 13824
rect 32548 13812 32554 13864
rect 32582 13812 32588 13864
rect 32640 13852 32646 13864
rect 33410 13852 33416 13864
rect 32640 13824 33416 13852
rect 32640 13812 32646 13824
rect 33410 13812 33416 13824
rect 33468 13812 33474 13864
rect 34054 13812 34060 13864
rect 34112 13812 34118 13864
rect 34609 13855 34667 13861
rect 34609 13821 34621 13855
rect 34655 13821 34667 13855
rect 34609 13815 34667 13821
rect 31036 13756 31754 13784
rect 34624 13784 34652 13815
rect 34698 13784 34704 13796
rect 34624 13756 34704 13784
rect 34698 13744 34704 13756
rect 34756 13744 34762 13796
rect 35268 13793 35296 13880
rect 35897 13855 35955 13861
rect 35897 13821 35909 13855
rect 35943 13852 35955 13855
rect 36630 13852 36636 13864
rect 35943 13824 36636 13852
rect 35943 13821 35955 13824
rect 35897 13815 35955 13821
rect 36630 13812 36636 13824
rect 36688 13812 36694 13864
rect 37645 13855 37703 13861
rect 37645 13821 37657 13855
rect 37691 13821 37703 13855
rect 37645 13815 37703 13821
rect 45189 13855 45247 13861
rect 45189 13821 45201 13855
rect 45235 13852 45247 13855
rect 46750 13852 46756 13864
rect 45235 13824 46756 13852
rect 45235 13821 45247 13824
rect 45189 13815 45247 13821
rect 35253 13787 35311 13793
rect 35253 13753 35265 13787
rect 35299 13753 35311 13787
rect 35253 13747 35311 13753
rect 36446 13744 36452 13796
rect 36504 13784 36510 13796
rect 36725 13787 36783 13793
rect 36725 13784 36737 13787
rect 36504 13756 36737 13784
rect 36504 13744 36510 13756
rect 36725 13753 36737 13756
rect 36771 13753 36783 13787
rect 37660 13784 37688 13815
rect 46750 13812 46756 13824
rect 46808 13812 46814 13864
rect 46934 13812 46940 13864
rect 46992 13812 46998 13864
rect 47228 13852 47256 13883
rect 49326 13880 49332 13932
rect 49384 13880 49390 13932
rect 47670 13852 47676 13864
rect 47228 13824 47676 13852
rect 47670 13812 47676 13824
rect 47728 13812 47734 13864
rect 47762 13812 47768 13864
rect 47820 13852 47826 13864
rect 49344 13852 49372 13880
rect 47820 13824 49372 13852
rect 47820 13812 47826 13824
rect 38194 13784 38200 13796
rect 37660 13756 38200 13784
rect 36725 13747 36783 13753
rect 38194 13744 38200 13756
rect 38252 13744 38258 13796
rect 46952 13784 46980 13812
rect 47029 13787 47087 13793
rect 47029 13784 47041 13787
rect 46952 13756 47041 13784
rect 47029 13753 47041 13756
rect 47075 13753 47087 13787
rect 47029 13747 47087 13753
rect 20036 13688 21036 13716
rect 19968 13679 19984 13685
rect 19978 13676 19984 13679
rect 20036 13676 20042 13688
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 27430 13716 27436 13728
rect 22796 13688 27436 13716
rect 22796 13676 22802 13688
rect 27430 13676 27436 13688
rect 27488 13676 27494 13728
rect 30834 13676 30840 13728
rect 30892 13716 30898 13728
rect 33799 13719 33857 13725
rect 33799 13716 33811 13719
rect 30892 13688 33811 13716
rect 30892 13676 30898 13688
rect 33799 13685 33811 13688
rect 33845 13716 33857 13719
rect 36170 13716 36176 13728
rect 33845 13688 36176 13716
rect 33845 13685 33857 13688
rect 33799 13679 33857 13685
rect 36170 13676 36176 13688
rect 36228 13676 36234 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 9646 13484 12112 13512
rect 9646 13444 9674 13484
rect 2976 13416 9674 13444
rect 12084 13444 12112 13484
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13504 13484 13645 13512
rect 13504 13472 13510 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 13998 13512 14004 13524
rect 13955 13484 14004 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 13998 13472 14004 13484
rect 14056 13512 14062 13524
rect 14918 13512 14924 13524
rect 14056 13484 14924 13512
rect 14056 13472 14062 13484
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 17954 13512 17960 13524
rect 15396 13484 17960 13512
rect 14277 13447 14335 13453
rect 14277 13444 14289 13447
rect 12084 13416 14289 13444
rect 1762 13336 1768 13388
rect 1820 13336 1826 13388
rect 2976 13317 3004 13416
rect 14277 13413 14289 13416
rect 14323 13413 14335 13447
rect 14277 13407 14335 13413
rect 10778 13336 10784 13388
rect 10836 13336 10842 13388
rect 12526 13336 12532 13388
rect 12584 13336 12590 13388
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12860 13348 13093 13376
rect 12860 13336 12866 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 14826 13376 14832 13388
rect 13081 13339 13139 13345
rect 13188 13348 14832 13376
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13277 3019 13311
rect 12544 13308 12572 13336
rect 13188 13308 13216 13348
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 15396 13385 15424 13484
rect 17954 13472 17960 13484
rect 18012 13512 18018 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 18012 13484 18153 13512
rect 18012 13472 18018 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 18322 13512 18328 13524
rect 18187 13484 18328 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18322 13472 18328 13484
rect 18380 13472 18386 13524
rect 19426 13472 19432 13524
rect 19484 13512 19490 13524
rect 20070 13512 20076 13524
rect 19484 13484 20076 13512
rect 19484 13472 19490 13484
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20254 13472 20260 13524
rect 20312 13512 20318 13524
rect 20441 13515 20499 13521
rect 20441 13512 20453 13515
rect 20312 13484 20453 13512
rect 20312 13472 20318 13484
rect 20441 13481 20453 13484
rect 20487 13481 20499 13515
rect 20441 13475 20499 13481
rect 20898 13472 20904 13524
rect 20956 13472 20962 13524
rect 22738 13512 22744 13524
rect 22572 13484 22744 13512
rect 20346 13404 20352 13456
rect 20404 13444 20410 13456
rect 22097 13447 22155 13453
rect 22097 13444 22109 13447
rect 20404 13416 22109 13444
rect 20404 13404 20410 13416
rect 22097 13413 22109 13416
rect 22143 13413 22155 13447
rect 22097 13407 22155 13413
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 15470 13336 15476 13388
rect 15528 13336 15534 13388
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 15804 13348 16405 13376
rect 15804 13336 15810 13348
rect 16393 13345 16405 13348
rect 16439 13376 16451 13379
rect 18966 13376 18972 13388
rect 16439 13348 18972 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13376 19947 13379
rect 19978 13376 19984 13388
rect 19935 13348 19984 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 20990 13336 20996 13388
rect 21048 13376 21054 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 21048 13348 21373 13376
rect 21048 13336 21054 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 21542 13336 21548 13388
rect 21600 13336 21606 13388
rect 22572 13385 22600 13484
rect 22738 13472 22744 13484
rect 22796 13472 22802 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 24029 13515 24087 13521
rect 24029 13512 24041 13515
rect 23716 13484 24041 13512
rect 23716 13472 23722 13484
rect 24029 13481 24041 13484
rect 24075 13481 24087 13515
rect 24029 13475 24087 13481
rect 25590 13472 25596 13524
rect 25648 13472 25654 13524
rect 28169 13515 28227 13521
rect 28169 13481 28181 13515
rect 28215 13512 28227 13515
rect 28350 13512 28356 13524
rect 28215 13484 28356 13512
rect 28215 13481 28227 13484
rect 28169 13475 28227 13481
rect 28350 13472 28356 13484
rect 28408 13512 28414 13524
rect 28902 13512 28908 13524
rect 28408 13484 28908 13512
rect 28408 13472 28414 13484
rect 28902 13472 28908 13484
rect 28960 13472 28966 13524
rect 29181 13515 29239 13521
rect 29181 13481 29193 13515
rect 29227 13512 29239 13515
rect 33778 13512 33784 13524
rect 29227 13484 33784 13512
rect 29227 13481 29239 13484
rect 29181 13475 29239 13481
rect 33778 13472 33784 13484
rect 33836 13472 33842 13524
rect 35621 13515 35679 13521
rect 35621 13481 35633 13515
rect 35667 13512 35679 13515
rect 36262 13512 36268 13524
rect 35667 13484 36268 13512
rect 35667 13481 35679 13484
rect 35621 13475 35679 13481
rect 36262 13472 36268 13484
rect 36320 13472 36326 13524
rect 37826 13512 37832 13524
rect 36556 13484 37832 13512
rect 24302 13444 24308 13456
rect 22756 13416 24308 13444
rect 22756 13385 22784 13416
rect 24302 13404 24308 13416
rect 24360 13404 24366 13456
rect 25222 13444 25228 13456
rect 24964 13416 25228 13444
rect 22557 13379 22615 13385
rect 22557 13345 22569 13379
rect 22603 13345 22615 13379
rect 22557 13339 22615 13345
rect 22741 13379 22799 13385
rect 22741 13345 22753 13379
rect 22787 13345 22799 13379
rect 22741 13339 22799 13345
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13376 23535 13379
rect 23523 13348 23980 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 12544 13280 13216 13308
rect 2961 13271 3019 13277
rect 14458 13268 14464 13320
rect 14516 13268 14522 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 14976 13280 15516 13308
rect 14976 13268 14982 13280
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 10505 13243 10563 13249
rect 10505 13240 10517 13243
rect 9088 13212 10517 13240
rect 9088 13200 9094 13212
rect 10505 13209 10517 13212
rect 10551 13240 10563 13243
rect 11054 13240 11060 13252
rect 10551 13212 11060 13240
rect 10551 13209 10563 13212
rect 10505 13203 10563 13209
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 14829 13243 14887 13249
rect 14829 13240 14841 13243
rect 12282 13212 13768 13240
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 12360 13172 12388 13212
rect 13740 13184 13768 13212
rect 14016 13212 14841 13240
rect 14016 13184 14044 13212
rect 14829 13209 14841 13212
rect 14875 13240 14887 13243
rect 15010 13240 15016 13252
rect 14875 13212 15016 13240
rect 14875 13209 14887 13212
rect 14829 13203 14887 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 15488 13240 15516 13280
rect 15562 13268 15568 13320
rect 15620 13268 15626 13320
rect 16298 13308 16304 13320
rect 15672 13280 16304 13308
rect 15672 13240 15700 13280
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 18046 13268 18052 13320
rect 18104 13308 18110 13320
rect 22465 13311 22523 13317
rect 18104 13280 22094 13308
rect 18104 13268 18110 13280
rect 16669 13243 16727 13249
rect 15488 13212 15700 13240
rect 15764 13212 16620 13240
rect 11756 13144 12388 13172
rect 11756 13132 11762 13144
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 13998 13172 14004 13184
rect 13780 13144 14004 13172
rect 13780 13132 13786 13144
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 15764 13172 15792 13212
rect 14148 13144 15792 13172
rect 14148 13132 14154 13144
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 15933 13175 15991 13181
rect 15933 13172 15945 13175
rect 15896 13144 15945 13172
rect 15896 13132 15902 13144
rect 15933 13141 15945 13144
rect 15979 13141 15991 13175
rect 16592 13172 16620 13212
rect 16669 13209 16681 13243
rect 16715 13240 16727 13243
rect 16758 13240 16764 13252
rect 16715 13212 16764 13240
rect 16715 13209 16727 13212
rect 16669 13203 16727 13209
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 17126 13200 17132 13252
rect 17184 13200 17190 13252
rect 18877 13243 18935 13249
rect 18877 13209 18889 13243
rect 18923 13240 18935 13243
rect 20073 13243 20131 13249
rect 20073 13240 20085 13243
rect 18923 13212 20085 13240
rect 18923 13209 18935 13212
rect 18877 13203 18935 13209
rect 20073 13209 20085 13212
rect 20119 13209 20131 13243
rect 20073 13203 20131 13209
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 21634 13240 21640 13252
rect 21048 13212 21640 13240
rect 21048 13200 21054 13212
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 22066 13240 22094 13280
rect 22465 13277 22477 13311
rect 22511 13308 22523 13311
rect 23661 13311 23719 13317
rect 22511 13280 23612 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 23382 13240 23388 13252
rect 22066 13212 23388 13240
rect 23382 13200 23388 13212
rect 23440 13200 23446 13252
rect 23584 13240 23612 13280
rect 23661 13277 23673 13311
rect 23707 13308 23719 13311
rect 23842 13308 23848 13320
rect 23707 13280 23848 13308
rect 23707 13277 23719 13280
rect 23661 13271 23719 13277
rect 23842 13268 23848 13280
rect 23900 13268 23906 13320
rect 23952 13308 23980 13348
rect 24964 13308 24992 13416
rect 25222 13404 25228 13416
rect 25280 13404 25286 13456
rect 29914 13444 29920 13456
rect 28552 13416 29920 13444
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13376 25099 13379
rect 26050 13376 26056 13388
rect 25087 13348 26056 13376
rect 25087 13345 25099 13348
rect 25041 13339 25099 13345
rect 26050 13336 26056 13348
rect 26108 13336 26114 13388
rect 28552 13385 28580 13416
rect 29914 13404 29920 13416
rect 29972 13404 29978 13456
rect 33321 13447 33379 13453
rect 33321 13413 33333 13447
rect 33367 13413 33379 13447
rect 33321 13407 33379 13413
rect 28537 13379 28595 13385
rect 28537 13345 28549 13379
rect 28583 13345 28595 13379
rect 28537 13339 28595 13345
rect 29822 13336 29828 13388
rect 29880 13336 29886 13388
rect 30009 13379 30067 13385
rect 30009 13345 30021 13379
rect 30055 13376 30067 13379
rect 30374 13376 30380 13388
rect 30055 13348 30380 13376
rect 30055 13345 30067 13348
rect 30009 13339 30067 13345
rect 30374 13336 30380 13348
rect 30432 13336 30438 13388
rect 31113 13379 31171 13385
rect 31113 13345 31125 13379
rect 31159 13345 31171 13379
rect 31113 13339 31171 13345
rect 23952 13280 24992 13308
rect 25130 13268 25136 13320
rect 25188 13308 25194 13320
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 25188 13280 25237 13308
rect 25188 13268 25194 13280
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 27798 13268 27804 13320
rect 27856 13308 27862 13320
rect 28813 13311 28871 13317
rect 27856 13280 28764 13308
rect 27856 13268 27862 13280
rect 24210 13240 24216 13252
rect 23584 13212 24216 13240
rect 24210 13200 24216 13212
rect 24268 13200 24274 13252
rect 25866 13240 25872 13252
rect 24320 13212 25872 13240
rect 19794 13172 19800 13184
rect 16592 13144 19800 13172
rect 15933 13135 15991 13141
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 19978 13132 19984 13184
rect 20036 13132 20042 13184
rect 21266 13132 21272 13184
rect 21324 13132 21330 13184
rect 23569 13175 23627 13181
rect 23569 13141 23581 13175
rect 23615 13172 23627 13175
rect 23658 13172 23664 13184
rect 23615 13144 23664 13172
rect 23615 13141 23627 13144
rect 23569 13135 23627 13141
rect 23658 13132 23664 13144
rect 23716 13132 23722 13184
rect 23842 13132 23848 13184
rect 23900 13172 23906 13184
rect 24320 13172 24348 13212
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 26694 13200 26700 13252
rect 26752 13240 26758 13252
rect 26789 13243 26847 13249
rect 26789 13240 26801 13243
rect 26752 13212 26801 13240
rect 26752 13200 26758 13212
rect 26789 13209 26801 13212
rect 26835 13240 26847 13243
rect 27525 13243 27583 13249
rect 27525 13240 27537 13243
rect 26835 13212 27537 13240
rect 26835 13209 26847 13212
rect 26789 13203 26847 13209
rect 27525 13209 27537 13212
rect 27571 13240 27583 13243
rect 28442 13240 28448 13252
rect 27571 13212 28448 13240
rect 27571 13209 27583 13212
rect 27525 13203 27583 13209
rect 28442 13200 28448 13212
rect 28500 13200 28506 13252
rect 28736 13240 28764 13280
rect 28813 13277 28825 13311
rect 28859 13308 28871 13311
rect 28994 13308 29000 13320
rect 28859 13280 29000 13308
rect 28859 13277 28871 13280
rect 28813 13271 28871 13277
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30190 13308 30196 13320
rect 30147 13280 30196 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 31128 13308 31156 13339
rect 31570 13336 31576 13388
rect 31628 13376 31634 13388
rect 33336 13376 33364 13407
rect 34422 13404 34428 13456
rect 34480 13444 34486 13456
rect 36173 13447 36231 13453
rect 36173 13444 36185 13447
rect 34480 13416 36185 13444
rect 34480 13404 34486 13416
rect 36173 13413 36185 13416
rect 36219 13413 36231 13447
rect 36173 13407 36231 13413
rect 31628 13348 33364 13376
rect 31628 13336 31634 13348
rect 33686 13336 33692 13388
rect 33744 13376 33750 13388
rect 33873 13379 33931 13385
rect 33873 13376 33885 13379
rect 33744 13348 33885 13376
rect 33744 13336 33750 13348
rect 33873 13345 33885 13348
rect 33919 13376 33931 13379
rect 34333 13379 34391 13385
rect 34333 13376 34345 13379
rect 33919 13348 34345 13376
rect 33919 13345 33931 13348
rect 33873 13339 33931 13345
rect 34333 13345 34345 13348
rect 34379 13345 34391 13379
rect 34333 13339 34391 13345
rect 35069 13379 35127 13385
rect 35069 13345 35081 13379
rect 35115 13376 35127 13379
rect 36556 13376 36584 13484
rect 37826 13472 37832 13484
rect 37884 13472 37890 13524
rect 38194 13472 38200 13524
rect 38252 13472 38258 13524
rect 38565 13515 38623 13521
rect 38565 13481 38577 13515
rect 38611 13512 38623 13515
rect 38838 13512 38844 13524
rect 38611 13484 38844 13512
rect 38611 13481 38623 13484
rect 38565 13475 38623 13481
rect 38838 13472 38844 13484
rect 38896 13512 38902 13524
rect 39482 13512 39488 13524
rect 38896 13484 39488 13512
rect 38896 13472 38902 13484
rect 39482 13472 39488 13484
rect 39540 13512 39546 13524
rect 39577 13515 39635 13521
rect 39577 13512 39589 13515
rect 39540 13484 39589 13512
rect 39540 13472 39546 13484
rect 39577 13481 39589 13484
rect 39623 13481 39635 13515
rect 39577 13475 39635 13481
rect 47673 13515 47731 13521
rect 47673 13481 47685 13515
rect 47719 13512 47731 13515
rect 47762 13512 47768 13524
rect 47719 13484 47768 13512
rect 47719 13481 47731 13484
rect 47673 13475 47731 13481
rect 47762 13472 47768 13484
rect 47820 13472 47826 13524
rect 35115 13348 36584 13376
rect 35115 13345 35127 13348
rect 35069 13339 35127 13345
rect 36722 13336 36728 13388
rect 36780 13376 36786 13388
rect 39574 13376 39580 13388
rect 36780 13348 39580 13376
rect 36780 13336 36786 13348
rect 39574 13336 39580 13348
rect 39632 13336 39638 13388
rect 30300 13280 31156 13308
rect 29730 13240 29736 13252
rect 28736 13212 29736 13240
rect 29730 13200 29736 13212
rect 29788 13240 29794 13252
rect 30300 13240 30328 13280
rect 31478 13268 31484 13320
rect 31536 13268 31542 13320
rect 32861 13311 32919 13317
rect 32861 13277 32873 13311
rect 32907 13308 32919 13311
rect 34054 13308 34060 13320
rect 32907 13280 34060 13308
rect 32907 13277 32919 13280
rect 32861 13271 32919 13277
rect 34054 13268 34060 13280
rect 34112 13268 34118 13320
rect 34882 13268 34888 13320
rect 34940 13308 34946 13320
rect 36449 13311 36507 13317
rect 36449 13308 36461 13311
rect 34940 13280 36461 13308
rect 34940 13268 34946 13280
rect 36449 13277 36461 13280
rect 36495 13277 36507 13311
rect 36449 13271 36507 13277
rect 32585 13243 32643 13249
rect 29788 13212 30328 13240
rect 30484 13212 31340 13240
rect 29788 13200 29794 13212
rect 23900 13144 24348 13172
rect 23900 13132 23906 13144
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 25133 13175 25191 13181
rect 25133 13172 25145 13175
rect 24544 13144 25145 13172
rect 24544 13132 24550 13144
rect 25133 13141 25145 13144
rect 25179 13172 25191 13175
rect 25958 13172 25964 13184
rect 25179 13144 25964 13172
rect 25179 13141 25191 13144
rect 25133 13135 25191 13141
rect 25958 13132 25964 13144
rect 26016 13132 26022 13184
rect 26050 13132 26056 13184
rect 26108 13132 26114 13184
rect 27706 13132 27712 13184
rect 27764 13132 27770 13184
rect 27893 13175 27951 13181
rect 27893 13141 27905 13175
rect 27939 13172 27951 13175
rect 28534 13172 28540 13184
rect 27939 13144 28540 13172
rect 27939 13141 27951 13144
rect 27893 13135 27951 13141
rect 28534 13132 28540 13144
rect 28592 13132 28598 13184
rect 28718 13132 28724 13184
rect 28776 13132 28782 13184
rect 30484 13181 30512 13212
rect 30469 13175 30527 13181
rect 30469 13141 30481 13175
rect 30515 13141 30527 13175
rect 31312 13172 31340 13212
rect 32585 13209 32597 13243
rect 32631 13240 32643 13243
rect 33962 13240 33968 13252
rect 32631 13212 33968 13240
rect 32631 13209 32643 13212
rect 32585 13203 32643 13209
rect 33962 13200 33968 13212
rect 34020 13200 34026 13252
rect 35253 13243 35311 13249
rect 35253 13209 35265 13243
rect 35299 13240 35311 13243
rect 35894 13240 35900 13252
rect 35299 13212 35900 13240
rect 35299 13209 35311 13212
rect 35253 13203 35311 13209
rect 35894 13200 35900 13212
rect 35952 13200 35958 13252
rect 31662 13172 31668 13184
rect 31312 13144 31668 13172
rect 30469 13135 30527 13141
rect 31662 13132 31668 13144
rect 31720 13132 31726 13184
rect 33410 13132 33416 13184
rect 33468 13172 33474 13184
rect 33689 13175 33747 13181
rect 33689 13172 33701 13175
rect 33468 13144 33701 13172
rect 33468 13132 33474 13144
rect 33689 13141 33701 13144
rect 33735 13141 33747 13175
rect 33689 13135 33747 13141
rect 33781 13175 33839 13181
rect 33781 13141 33793 13175
rect 33827 13172 33839 13175
rect 34146 13172 34152 13184
rect 33827 13144 34152 13172
rect 33827 13141 33839 13144
rect 33781 13135 33839 13141
rect 34146 13132 34152 13144
rect 34204 13132 34210 13184
rect 35158 13132 35164 13184
rect 35216 13132 35222 13184
rect 35710 13132 35716 13184
rect 35768 13172 35774 13184
rect 35989 13175 36047 13181
rect 35989 13172 36001 13175
rect 35768 13144 36001 13172
rect 35768 13132 35774 13144
rect 35989 13141 36001 13144
rect 36035 13141 36047 13175
rect 36464 13172 36492 13271
rect 41322 13268 41328 13320
rect 41380 13268 41386 13320
rect 46750 13268 46756 13320
rect 46808 13308 46814 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 46808 13280 47961 13308
rect 46808 13268 46814 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 49142 13268 49148 13320
rect 49200 13268 49206 13320
rect 36630 13200 36636 13252
rect 36688 13240 36694 13252
rect 36725 13243 36783 13249
rect 36725 13240 36737 13243
rect 36688 13212 36737 13240
rect 36688 13200 36694 13212
rect 36725 13209 36737 13212
rect 36771 13209 36783 13243
rect 38838 13240 38844 13252
rect 37950 13212 38844 13240
rect 36725 13203 36783 13209
rect 38838 13200 38844 13212
rect 38896 13200 38902 13252
rect 37458 13172 37464 13184
rect 36464 13144 37464 13172
rect 35989 13135 36047 13141
rect 37458 13132 37464 13144
rect 37516 13132 37522 13184
rect 37642 13132 37648 13184
rect 37700 13172 37706 13184
rect 39298 13172 39304 13184
rect 37700 13144 39304 13172
rect 37700 13132 37706 13144
rect 39298 13132 39304 13144
rect 39356 13132 39362 13184
rect 41509 13175 41567 13181
rect 41509 13141 41521 13175
rect 41555 13172 41567 13175
rect 45922 13172 45928 13184
rect 41555 13144 45928 13172
rect 41555 13141 41567 13144
rect 41509 13135 41567 13141
rect 45922 13132 45928 13144
rect 45980 13132 45986 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 1765 12971 1823 12977
rect 1765 12937 1777 12971
rect 1811 12968 1823 12971
rect 9490 12968 9496 12980
rect 1811 12940 9496 12968
rect 1811 12937 1823 12940
rect 1765 12931 1823 12937
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 11330 12928 11336 12980
rect 11388 12928 11394 12980
rect 11974 12928 11980 12980
rect 12032 12928 12038 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12805 12971 12863 12977
rect 12805 12968 12817 12971
rect 12584 12940 12817 12968
rect 12584 12928 12590 12940
rect 12805 12937 12817 12940
rect 12851 12968 12863 12971
rect 12894 12968 12900 12980
rect 12851 12940 12900 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13262 12968 13268 12980
rect 13127 12940 13268 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13630 12928 13636 12980
rect 13688 12968 13694 12980
rect 13688 12940 14872 12968
rect 13688 12928 13694 12940
rect 1302 12860 1308 12912
rect 1360 12900 1366 12912
rect 1673 12903 1731 12909
rect 1673 12900 1685 12903
rect 1360 12872 1685 12900
rect 1360 12860 1366 12872
rect 1673 12869 1685 12872
rect 1719 12900 1731 12903
rect 2133 12903 2191 12909
rect 2133 12900 2145 12903
rect 1719 12872 2145 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 2133 12869 2145 12872
rect 2179 12869 2191 12903
rect 2133 12863 2191 12869
rect 11149 12903 11207 12909
rect 11149 12869 11161 12903
rect 11195 12900 11207 12903
rect 11698 12900 11704 12912
rect 11195 12872 11704 12900
rect 11195 12869 11207 12872
rect 11149 12863 11207 12869
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 13998 12860 14004 12912
rect 14056 12860 14062 12912
rect 14550 12860 14556 12912
rect 14608 12860 14614 12912
rect 14844 12841 14872 12940
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15252 12940 15853 12968
rect 15252 12928 15258 12940
rect 15841 12937 15853 12940
rect 15887 12968 15899 12971
rect 20717 12971 20775 12977
rect 15887 12940 19104 12968
rect 15887 12937 15899 12940
rect 15841 12931 15899 12937
rect 15933 12903 15991 12909
rect 15933 12869 15945 12903
rect 15979 12900 15991 12903
rect 16390 12900 16396 12912
rect 15979 12872 16396 12900
rect 15979 12869 15991 12872
rect 15933 12863 15991 12869
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 16666 12860 16672 12912
rect 16724 12900 16730 12912
rect 17034 12900 17040 12912
rect 16724 12872 17040 12900
rect 16724 12860 16730 12872
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 18693 12903 18751 12909
rect 18693 12869 18705 12903
rect 18739 12900 18751 12903
rect 18966 12900 18972 12912
rect 18739 12872 18972 12900
rect 18739 12869 18751 12872
rect 18693 12863 18751 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 19076 12900 19104 12940
rect 20717 12937 20729 12971
rect 20763 12968 20775 12971
rect 20898 12968 20904 12980
rect 20763 12940 20904 12968
rect 20763 12937 20775 12940
rect 20717 12931 20775 12937
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21177 12971 21235 12977
rect 21177 12937 21189 12971
rect 21223 12968 21235 12971
rect 23385 12971 23443 12977
rect 21223 12940 23336 12968
rect 21223 12937 21235 12940
rect 21177 12931 21235 12937
rect 23308 12900 23336 12940
rect 23385 12937 23397 12971
rect 23431 12968 23443 12971
rect 23474 12968 23480 12980
rect 23431 12940 23480 12968
rect 23431 12937 23443 12940
rect 23385 12931 23443 12937
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 23658 12928 23664 12980
rect 23716 12968 23722 12980
rect 24394 12968 24400 12980
rect 23716 12940 24400 12968
rect 23716 12928 23722 12940
rect 23842 12900 23848 12912
rect 19076 12872 23244 12900
rect 23308 12872 23848 12900
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2516 12804 2881 12832
rect 1302 12656 1308 12708
rect 1360 12696 1366 12708
rect 2516 12705 2544 12804
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 14829 12835 14887 12841
rect 12115 12804 12434 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 12406 12764 12434 12804
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15746 12832 15752 12844
rect 14875 12804 15752 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 16758 12832 16764 12844
rect 15948 12804 16764 12832
rect 15948 12776 15976 12804
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 16942 12792 16948 12844
rect 17000 12792 17006 12844
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17368 12804 17877 12832
rect 17368 12792 17374 12804
rect 17865 12801 17877 12804
rect 17911 12832 17923 12835
rect 18874 12832 18880 12844
rect 17911 12804 18880 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19610 12792 19616 12844
rect 19668 12792 19674 12844
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 19852 12804 20361 12832
rect 19852 12792 19858 12804
rect 20349 12801 20361 12804
rect 20395 12832 20407 12835
rect 20990 12832 20996 12844
rect 20395 12804 20996 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 21910 12832 21916 12844
rect 21131 12804 21916 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 23017 12835 23075 12841
rect 23017 12801 23029 12835
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 13814 12764 13820 12776
rect 12406 12736 13820 12764
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 15657 12767 15715 12773
rect 15657 12733 15669 12767
rect 15703 12764 15715 12767
rect 15930 12764 15936 12776
rect 15703 12736 15936 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16574 12724 16580 12776
rect 16632 12724 16638 12776
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12764 17463 12767
rect 19518 12764 19524 12776
rect 17451 12736 19524 12764
rect 17451 12733 17463 12736
rect 17405 12727 17463 12733
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 19702 12724 19708 12776
rect 19760 12724 19766 12776
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20254 12764 20260 12776
rect 19935 12736 20260 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 20496 12736 21281 12764
rect 20496 12724 20502 12736
rect 21269 12733 21281 12736
rect 21315 12733 21327 12767
rect 21269 12727 21327 12733
rect 22002 12724 22008 12776
rect 22060 12724 22066 12776
rect 22738 12724 22744 12776
rect 22796 12724 22802 12776
rect 22922 12724 22928 12776
rect 22980 12724 22986 12776
rect 2501 12699 2559 12705
rect 2501 12696 2513 12699
rect 1360 12668 2513 12696
rect 1360 12656 1366 12668
rect 2501 12665 2513 12668
rect 2547 12665 2559 12699
rect 2501 12659 2559 12665
rect 15286 12656 15292 12708
rect 15344 12696 15350 12708
rect 16390 12696 16396 12708
rect 15344 12668 16396 12696
rect 15344 12656 15350 12668
rect 16390 12656 16396 12668
rect 16448 12656 16454 12708
rect 16592 12696 16620 12724
rect 19245 12699 19303 12705
rect 19245 12696 19257 12699
rect 16592 12668 19257 12696
rect 19245 12665 19257 12668
rect 19291 12665 19303 12699
rect 19245 12659 19303 12665
rect 20272 12668 20576 12696
rect 2314 12588 2320 12640
rect 2372 12588 2378 12640
rect 2866 12588 2872 12640
rect 2924 12628 2930 12640
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 2924 12600 3525 12628
rect 2924 12588 2930 12600
rect 3513 12597 3525 12600
rect 3559 12597 3571 12631
rect 3513 12591 3571 12597
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 12618 12628 12624 12640
rect 12483 12600 12624 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14090 12628 14096 12640
rect 13872 12600 14096 12628
rect 13872 12588 13878 12600
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 14182 12588 14188 12640
rect 14240 12628 14246 12640
rect 15010 12628 15016 12640
rect 14240 12600 15016 12628
rect 14240 12588 14246 12600
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 16301 12631 16359 12637
rect 16301 12597 16313 12631
rect 16347 12628 16359 12631
rect 16574 12628 16580 12640
rect 16347 12600 16580 12628
rect 16347 12597 16359 12600
rect 16301 12591 16359 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 20272 12628 20300 12668
rect 17092 12600 20300 12628
rect 20548 12628 20576 12668
rect 20990 12656 20996 12708
rect 21048 12696 21054 12708
rect 21450 12696 21456 12708
rect 21048 12668 21456 12696
rect 21048 12656 21054 12668
rect 21450 12656 21456 12668
rect 21508 12696 21514 12708
rect 23032 12696 23060 12795
rect 23216 12764 23244 12872
rect 23842 12860 23848 12872
rect 23900 12860 23906 12912
rect 23566 12764 23572 12776
rect 23216 12736 23572 12764
rect 23566 12724 23572 12736
rect 23624 12724 23630 12776
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 23952 12764 23980 12940
rect 24394 12928 24400 12940
rect 24452 12928 24458 12980
rect 24578 12928 24584 12980
rect 24636 12968 24642 12980
rect 24636 12940 25544 12968
rect 24636 12928 24642 12940
rect 24854 12860 24860 12912
rect 24912 12860 24918 12912
rect 25314 12860 25320 12912
rect 25372 12860 25378 12912
rect 25516 12900 25544 12940
rect 25958 12928 25964 12980
rect 26016 12968 26022 12980
rect 26697 12971 26755 12977
rect 26697 12968 26709 12971
rect 26016 12940 26709 12968
rect 26016 12928 26022 12940
rect 26697 12937 26709 12940
rect 26743 12968 26755 12971
rect 27062 12968 27068 12980
rect 26743 12940 27068 12968
rect 26743 12937 26755 12940
rect 26697 12931 26755 12937
rect 27062 12928 27068 12940
rect 27120 12928 27126 12980
rect 28534 12928 28540 12980
rect 28592 12968 28598 12980
rect 28592 12940 31616 12968
rect 28592 12928 28598 12940
rect 26145 12903 26203 12909
rect 25516 12872 25636 12900
rect 25608 12841 25636 12872
rect 26145 12869 26157 12903
rect 26191 12900 26203 12903
rect 26234 12900 26240 12912
rect 26191 12872 26240 12900
rect 26191 12869 26203 12872
rect 26145 12863 26203 12869
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 24946 12764 24952 12776
rect 23716 12736 23980 12764
rect 24136 12736 24952 12764
rect 23716 12724 23722 12736
rect 24136 12708 24164 12736
rect 24946 12724 24952 12736
rect 25004 12724 25010 12776
rect 25222 12724 25228 12776
rect 25280 12764 25286 12776
rect 26160 12764 26188 12863
rect 26234 12860 26240 12872
rect 26292 12860 26298 12912
rect 27154 12860 27160 12912
rect 27212 12860 27218 12912
rect 28442 12860 28448 12912
rect 28500 12860 28506 12912
rect 28920 12909 28948 12940
rect 28905 12903 28963 12909
rect 28905 12869 28917 12903
rect 28951 12869 28963 12903
rect 28905 12863 28963 12869
rect 29362 12860 29368 12912
rect 29420 12900 29426 12912
rect 29549 12903 29607 12909
rect 29549 12900 29561 12903
rect 29420 12872 29561 12900
rect 29420 12860 29426 12872
rect 29549 12869 29561 12872
rect 29595 12900 29607 12903
rect 29730 12900 29736 12912
rect 29595 12872 29736 12900
rect 29595 12869 29607 12872
rect 29549 12863 29607 12869
rect 29730 12860 29736 12872
rect 29788 12860 29794 12912
rect 31588 12900 31616 12940
rect 31754 12928 31760 12980
rect 31812 12968 31818 12980
rect 32585 12971 32643 12977
rect 32585 12968 32597 12971
rect 31812 12940 32597 12968
rect 31812 12928 31818 12940
rect 32585 12937 32597 12940
rect 32631 12937 32643 12971
rect 32585 12931 32643 12937
rect 34054 12928 34060 12980
rect 34112 12968 34118 12980
rect 34112 12940 34836 12968
rect 34112 12928 34118 12940
rect 32030 12900 32036 12912
rect 31588 12872 32036 12900
rect 32030 12860 32036 12872
rect 32088 12860 32094 12912
rect 32122 12860 32128 12912
rect 32180 12900 32186 12912
rect 32766 12900 32772 12912
rect 32180 12872 32772 12900
rect 32180 12860 32186 12872
rect 32766 12860 32772 12872
rect 32824 12860 32830 12912
rect 33410 12860 33416 12912
rect 33468 12900 33474 12912
rect 34422 12900 34428 12912
rect 33468 12872 34428 12900
rect 33468 12860 33474 12872
rect 34422 12860 34428 12872
rect 34480 12860 34486 12912
rect 34808 12909 34836 12940
rect 34974 12928 34980 12980
rect 35032 12968 35038 12980
rect 35805 12971 35863 12977
rect 35805 12968 35817 12971
rect 35032 12940 35817 12968
rect 35032 12928 35038 12940
rect 35805 12937 35817 12940
rect 35851 12968 35863 12971
rect 36633 12971 36691 12977
rect 36633 12968 36645 12971
rect 35851 12940 36645 12968
rect 35851 12937 35863 12940
rect 35805 12931 35863 12937
rect 36633 12937 36645 12940
rect 36679 12968 36691 12971
rect 36722 12968 36728 12980
rect 36679 12940 36728 12968
rect 36679 12937 36691 12940
rect 36633 12931 36691 12937
rect 36722 12928 36728 12940
rect 36780 12928 36786 12980
rect 37182 12928 37188 12980
rect 37240 12968 37246 12980
rect 40310 12968 40316 12980
rect 37240 12940 40316 12968
rect 37240 12928 37246 12940
rect 40310 12928 40316 12940
rect 40368 12928 40374 12980
rect 34793 12903 34851 12909
rect 34793 12869 34805 12903
rect 34839 12900 34851 12903
rect 34882 12900 34888 12912
rect 34839 12872 34888 12900
rect 34839 12869 34851 12872
rect 34793 12863 34851 12869
rect 34882 12860 34888 12872
rect 34940 12860 34946 12912
rect 36906 12860 36912 12912
rect 36964 12900 36970 12912
rect 37001 12903 37059 12909
rect 37001 12900 37013 12903
rect 36964 12872 37013 12900
rect 36964 12860 36970 12872
rect 37001 12869 37013 12872
rect 37047 12869 37059 12903
rect 37642 12900 37648 12912
rect 37001 12863 37059 12869
rect 37310 12872 37648 12900
rect 29181 12835 29239 12841
rect 29181 12801 29193 12835
rect 29227 12832 29239 12835
rect 30006 12832 30012 12844
rect 29227 12804 30012 12832
rect 29227 12801 29239 12804
rect 29181 12795 29239 12801
rect 30006 12792 30012 12804
rect 30064 12792 30070 12844
rect 31386 12792 31392 12844
rect 31444 12792 31450 12844
rect 31754 12792 31760 12844
rect 31812 12832 31818 12844
rect 32677 12835 32735 12841
rect 32677 12832 32689 12835
rect 31812 12804 32689 12832
rect 31812 12792 31818 12804
rect 32677 12801 32689 12804
rect 32723 12801 32735 12835
rect 32677 12795 32735 12801
rect 33318 12792 33324 12844
rect 33376 12832 33382 12844
rect 34057 12835 34115 12841
rect 34057 12832 34069 12835
rect 33376 12804 34069 12832
rect 33376 12792 33382 12804
rect 34057 12801 34069 12804
rect 34103 12801 34115 12835
rect 34057 12795 34115 12801
rect 34606 12792 34612 12844
rect 34664 12832 34670 12844
rect 36817 12835 36875 12841
rect 36817 12832 36829 12835
rect 34664 12804 35756 12832
rect 34664 12792 34670 12804
rect 25280 12736 26188 12764
rect 25280 12724 25286 12736
rect 29638 12724 29644 12776
rect 29696 12764 29702 12776
rect 30285 12767 30343 12773
rect 30285 12764 30297 12767
rect 29696 12736 30297 12764
rect 29696 12724 29702 12736
rect 30285 12733 30297 12736
rect 30331 12733 30343 12767
rect 30285 12727 30343 12733
rect 32030 12724 32036 12776
rect 32088 12764 32094 12776
rect 32401 12767 32459 12773
rect 32401 12764 32413 12767
rect 32088 12736 32413 12764
rect 32088 12724 32094 12736
rect 32401 12733 32413 12736
rect 32447 12733 32459 12767
rect 33686 12764 33692 12776
rect 32401 12727 32459 12733
rect 32968 12736 33692 12764
rect 21508 12668 23060 12696
rect 23845 12699 23903 12705
rect 21508 12656 21514 12668
rect 23845 12665 23857 12699
rect 23891 12696 23903 12699
rect 24118 12696 24124 12708
rect 23891 12668 24124 12696
rect 23891 12665 23903 12668
rect 23845 12659 23903 12665
rect 24118 12656 24124 12668
rect 24176 12656 24182 12708
rect 32968 12696 32996 12736
rect 33686 12724 33692 12736
rect 33744 12724 33750 12776
rect 35158 12724 35164 12776
rect 35216 12764 35222 12776
rect 35342 12764 35348 12776
rect 35216 12736 35348 12764
rect 35216 12724 35222 12736
rect 35342 12724 35348 12736
rect 35400 12764 35406 12776
rect 35728 12773 35756 12804
rect 35912 12804 36829 12832
rect 35529 12767 35587 12773
rect 35529 12764 35541 12767
rect 35400 12736 35541 12764
rect 35400 12724 35406 12736
rect 35529 12733 35541 12736
rect 35575 12733 35587 12767
rect 35529 12727 35587 12733
rect 35713 12767 35771 12773
rect 35713 12733 35725 12767
rect 35759 12764 35771 12767
rect 35802 12764 35808 12776
rect 35759 12736 35808 12764
rect 35759 12733 35771 12736
rect 35713 12727 35771 12733
rect 31680 12668 32996 12696
rect 33045 12699 33103 12705
rect 22922 12628 22928 12640
rect 20548 12600 22928 12628
rect 17092 12588 17098 12600
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 24854 12588 24860 12640
rect 24912 12628 24918 12640
rect 25682 12628 25688 12640
rect 24912 12600 25688 12628
rect 24912 12588 24918 12600
rect 25682 12588 25688 12600
rect 25740 12628 25746 12640
rect 25958 12628 25964 12640
rect 25740 12600 25964 12628
rect 25740 12588 25746 12600
rect 25958 12588 25964 12600
rect 26016 12588 26022 12640
rect 28810 12588 28816 12640
rect 28868 12628 28874 12640
rect 31680 12628 31708 12668
rect 33045 12665 33057 12699
rect 33091 12696 33103 12699
rect 34514 12696 34520 12708
rect 33091 12668 34520 12696
rect 33091 12665 33103 12668
rect 33045 12659 33103 12665
rect 34514 12656 34520 12668
rect 34572 12656 34578 12708
rect 35544 12696 35572 12727
rect 35802 12724 35808 12736
rect 35860 12724 35866 12776
rect 35912 12696 35940 12804
rect 36817 12801 36829 12804
rect 36863 12832 36875 12835
rect 37310 12832 37338 12872
rect 37642 12860 37648 12872
rect 37700 12860 37706 12912
rect 36863 12804 37338 12832
rect 36863 12801 36875 12804
rect 36817 12795 36875 12801
rect 37458 12792 37464 12844
rect 37516 12792 37522 12844
rect 38838 12792 38844 12844
rect 38896 12792 38902 12844
rect 40034 12792 40040 12844
rect 40092 12832 40098 12844
rect 40497 12835 40555 12841
rect 40497 12832 40509 12835
rect 40092 12804 40509 12832
rect 40092 12792 40098 12804
rect 40497 12801 40509 12804
rect 40543 12801 40555 12835
rect 40497 12795 40555 12801
rect 45922 12792 45928 12844
rect 45980 12792 45986 12844
rect 47210 12792 47216 12844
rect 47268 12832 47274 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47268 12804 47961 12832
rect 47268 12792 47274 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 49142 12792 49148 12844
rect 49200 12792 49206 12844
rect 36446 12724 36452 12776
rect 36504 12764 36510 12776
rect 37182 12764 37188 12776
rect 36504 12736 37188 12764
rect 36504 12724 36510 12736
rect 37182 12724 37188 12736
rect 37240 12724 37246 12776
rect 37737 12767 37795 12773
rect 37737 12733 37749 12767
rect 37783 12764 37795 12767
rect 38286 12764 38292 12776
rect 37783 12736 38292 12764
rect 37783 12733 37795 12736
rect 37737 12727 37795 12733
rect 38286 12724 38292 12736
rect 38344 12724 38350 12776
rect 39298 12724 39304 12776
rect 39356 12764 39362 12776
rect 39485 12767 39543 12773
rect 39485 12764 39497 12767
rect 39356 12736 39497 12764
rect 39356 12724 39362 12736
rect 39485 12733 39497 12736
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 35544 12668 35940 12696
rect 36173 12699 36231 12705
rect 36173 12665 36185 12699
rect 36219 12696 36231 12699
rect 40221 12699 40279 12705
rect 36219 12668 37596 12696
rect 36219 12665 36231 12668
rect 36173 12659 36231 12665
rect 28868 12600 31708 12628
rect 31757 12631 31815 12637
rect 28868 12588 28874 12600
rect 31757 12597 31769 12631
rect 31803 12628 31815 12631
rect 32306 12628 32312 12640
rect 31803 12600 32312 12628
rect 31803 12597 31815 12600
rect 31757 12591 31815 12597
rect 32306 12588 32312 12600
rect 32364 12628 32370 12640
rect 32582 12628 32588 12640
rect 32364 12600 32588 12628
rect 32364 12588 32370 12600
rect 32582 12588 32588 12600
rect 32640 12588 32646 12640
rect 32858 12588 32864 12640
rect 32916 12628 32922 12640
rect 33505 12631 33563 12637
rect 33505 12628 33517 12631
rect 32916 12600 33517 12628
rect 32916 12588 32922 12600
rect 33505 12597 33517 12600
rect 33551 12628 33563 12631
rect 33689 12631 33747 12637
rect 33689 12628 33701 12631
rect 33551 12600 33701 12628
rect 33551 12597 33563 12600
rect 33505 12591 33563 12597
rect 33689 12597 33701 12600
rect 33735 12597 33747 12631
rect 33689 12591 33747 12597
rect 35802 12588 35808 12640
rect 35860 12628 35866 12640
rect 36906 12628 36912 12640
rect 35860 12600 36912 12628
rect 35860 12588 35866 12600
rect 36906 12588 36912 12600
rect 36964 12588 36970 12640
rect 37568 12628 37596 12668
rect 40221 12665 40233 12699
rect 40267 12696 40279 12699
rect 46934 12696 46940 12708
rect 40267 12668 46940 12696
rect 40267 12665 40279 12668
rect 40221 12659 40279 12665
rect 46934 12656 46940 12668
rect 46992 12656 46998 12708
rect 39114 12628 39120 12640
rect 37568 12600 39120 12628
rect 39114 12588 39120 12600
rect 39172 12588 39178 12640
rect 46109 12631 46167 12637
rect 46109 12597 46121 12631
rect 46155 12628 46167 12631
rect 47946 12628 47952 12640
rect 46155 12600 47952 12628
rect 46155 12597 46167 12600
rect 46109 12591 46167 12597
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 3053 12427 3111 12433
rect 3053 12393 3065 12427
rect 3099 12424 3111 12427
rect 4338 12424 4344 12436
rect 3099 12396 4344 12424
rect 3099 12393 3111 12396
rect 3053 12387 3111 12393
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11790 12424 11796 12436
rect 11287 12396 11796 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 13722 12424 13728 12436
rect 13596 12396 13728 12424
rect 13596 12384 13602 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14240 12396 14381 12424
rect 14240 12384 14246 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 15853 12427 15911 12433
rect 15853 12424 15865 12427
rect 14369 12387 14427 12393
rect 14476 12396 15865 12424
rect 11054 12316 11060 12368
rect 11112 12356 11118 12368
rect 11112 12328 11836 12356
rect 11112 12316 11118 12328
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 5810 12288 5816 12300
rect 2179 12260 5816 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 10778 12288 10784 12300
rect 9539 12260 10784 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 10778 12248 10784 12260
rect 10836 12288 10842 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 10836 12260 11713 12288
rect 10836 12248 10842 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11808 12288 11836 12328
rect 13354 12316 13360 12368
rect 13412 12356 13418 12368
rect 14476 12356 14504 12396
rect 15853 12393 15865 12396
rect 15899 12424 15911 12427
rect 16114 12424 16120 12436
rect 15899 12396 16120 12424
rect 15899 12393 15911 12396
rect 15853 12387 15911 12393
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 17862 12424 17868 12436
rect 16224 12396 17868 12424
rect 16224 12368 16252 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 19392 12396 19441 12424
rect 19392 12384 19398 12396
rect 19429 12393 19441 12396
rect 19475 12393 19487 12427
rect 19429 12387 19487 12393
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 26050 12424 26056 12436
rect 21784 12396 26056 12424
rect 21784 12384 21790 12396
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 26326 12384 26332 12436
rect 26384 12424 26390 12436
rect 26970 12424 26976 12436
rect 26384 12396 26976 12424
rect 26384 12384 26390 12396
rect 26970 12384 26976 12396
rect 27028 12384 27034 12436
rect 27709 12427 27767 12433
rect 27709 12393 27721 12427
rect 27755 12424 27767 12427
rect 31754 12424 31760 12436
rect 27755 12396 31760 12424
rect 27755 12393 27767 12396
rect 27709 12387 27767 12393
rect 31754 12384 31760 12396
rect 31812 12384 31818 12436
rect 31864 12396 39252 12424
rect 13412 12328 14504 12356
rect 13412 12316 13418 12328
rect 16206 12316 16212 12368
rect 16264 12316 16270 12368
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 16448 12328 17356 12356
rect 16448 12316 16454 12328
rect 13722 12288 13728 12300
rect 11808 12260 13728 12288
rect 11701 12251 11759 12257
rect 13722 12248 13728 12260
rect 13780 12288 13786 12300
rect 15286 12288 15292 12300
rect 13780 12260 15292 12288
rect 13780 12248 13786 12260
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 15804 12260 16129 12288
rect 15804 12248 15810 12260
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 16485 12291 16543 12297
rect 16485 12257 16497 12291
rect 16531 12288 16543 12291
rect 16942 12288 16948 12300
rect 16531 12260 16948 12288
rect 16531 12257 16543 12260
rect 16485 12251 16543 12257
rect 2222 12180 2228 12232
rect 2280 12220 2286 12232
rect 2409 12223 2467 12229
rect 2409 12220 2421 12223
rect 2280 12192 2421 12220
rect 2280 12180 2286 12192
rect 2409 12189 2421 12192
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2866 12180 2872 12232
rect 2924 12180 2930 12232
rect 11606 12220 11612 12232
rect 10902 12192 11612 12220
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 9766 12112 9772 12164
rect 9824 12112 9830 12164
rect 11054 12112 11060 12164
rect 11112 12152 11118 12164
rect 11977 12155 12035 12161
rect 11977 12152 11989 12155
rect 11112 12124 11989 12152
rect 11112 12112 11118 12124
rect 11977 12121 11989 12124
rect 12023 12121 12035 12155
rect 13538 12152 13544 12164
rect 13202 12124 13544 12152
rect 11977 12115 12035 12121
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 13725 12155 13783 12161
rect 13725 12121 13737 12155
rect 13771 12152 13783 12155
rect 14458 12152 14464 12164
rect 13771 12124 14464 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 14458 12112 14464 12124
rect 14516 12112 14522 12164
rect 16500 12152 16528 12251
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17328 12297 17356 12328
rect 17402 12316 17408 12368
rect 17460 12356 17466 12368
rect 21266 12356 21272 12368
rect 17460 12328 19472 12356
rect 17460 12316 17466 12328
rect 19444 12300 19472 12328
rect 19536 12328 21272 12356
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12288 17371 12291
rect 17494 12288 17500 12300
rect 17359 12260 17500 12288
rect 17359 12257 17371 12260
rect 17313 12251 17371 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 19426 12248 19432 12300
rect 19484 12248 19490 12300
rect 17034 12180 17040 12232
rect 17092 12220 17098 12232
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 17092 12192 17141 12220
rect 17092 12180 17098 12192
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 19058 12180 19064 12232
rect 19116 12220 19122 12232
rect 19536 12220 19564 12328
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 21637 12359 21695 12365
rect 21637 12325 21649 12359
rect 21683 12356 21695 12359
rect 23750 12356 23756 12368
rect 21683 12328 23756 12356
rect 21683 12325 21695 12328
rect 21637 12319 21695 12325
rect 23750 12316 23756 12328
rect 23808 12316 23814 12368
rect 25958 12316 25964 12368
rect 26016 12356 26022 12368
rect 26694 12356 26700 12368
rect 26016 12328 26700 12356
rect 26016 12316 26022 12328
rect 26694 12316 26700 12328
rect 26752 12316 26758 12368
rect 31018 12316 31024 12368
rect 31076 12356 31082 12368
rect 31864 12356 31892 12396
rect 31076 12328 31892 12356
rect 39025 12359 39083 12365
rect 31076 12316 31082 12328
rect 39025 12325 39037 12359
rect 39071 12325 39083 12359
rect 39224 12356 39252 12396
rect 39298 12384 39304 12436
rect 39356 12384 39362 12436
rect 39482 12384 39488 12436
rect 39540 12384 39546 12436
rect 39942 12356 39948 12368
rect 39224 12328 39948 12356
rect 39025 12319 39083 12325
rect 19886 12248 19892 12300
rect 19944 12288 19950 12300
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19944 12260 19993 12288
rect 19944 12248 19950 12260
rect 19981 12257 19993 12260
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20625 12291 20683 12297
rect 20625 12257 20637 12291
rect 20671 12288 20683 12291
rect 20990 12288 20996 12300
rect 20671 12260 20996 12288
rect 20671 12257 20683 12260
rect 20625 12251 20683 12257
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 19116 12192 19564 12220
rect 19720 12192 19809 12220
rect 19116 12180 19122 12192
rect 15410 12124 16528 12152
rect 18141 12155 18199 12161
rect 18141 12121 18153 12155
rect 18187 12152 18199 12155
rect 18782 12152 18788 12164
rect 18187 12124 18788 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 18874 12112 18880 12164
rect 18932 12112 18938 12164
rect 19518 12112 19524 12164
rect 19576 12152 19582 12164
rect 19720 12152 19748 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 20530 12220 20536 12232
rect 19797 12183 19855 12189
rect 19996 12192 20536 12220
rect 19996 12152 20024 12192
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 21174 12180 21180 12232
rect 21232 12180 21238 12232
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 21726 12220 21732 12232
rect 21315 12192 21732 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21726 12180 21732 12192
rect 21784 12180 21790 12232
rect 22296 12220 22324 12251
rect 22370 12248 22376 12300
rect 22428 12248 22434 12300
rect 23474 12288 23480 12300
rect 22480 12260 23480 12288
rect 22480 12220 22508 12260
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 23658 12248 23664 12300
rect 23716 12248 23722 12300
rect 23937 12291 23995 12297
rect 23937 12257 23949 12291
rect 23983 12288 23995 12291
rect 24486 12288 24492 12300
rect 23983 12260 24492 12288
rect 23983 12257 23995 12260
rect 23937 12251 23995 12257
rect 24486 12248 24492 12260
rect 24544 12248 24550 12300
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 24946 12288 24952 12300
rect 24903 12260 24952 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 23676 12220 23704 12248
rect 22296 12192 22508 12220
rect 22756 12192 23704 12220
rect 19576 12124 19748 12152
rect 19812 12124 20024 12152
rect 19576 12112 19582 12124
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 14366 12084 14372 12096
rect 13044 12056 14372 12084
rect 13044 12044 13050 12056
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 14476 12084 14504 12112
rect 15654 12084 15660 12096
rect 14476 12056 15660 12084
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16758 12044 16764 12096
rect 16816 12044 16822 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 19812 12084 19840 12124
rect 20070 12112 20076 12164
rect 20128 12152 20134 12164
rect 21192 12152 21220 12180
rect 20128 12124 21220 12152
rect 20128 12112 20134 12124
rect 21450 12112 21456 12164
rect 21508 12152 21514 12164
rect 22465 12155 22523 12161
rect 22465 12152 22477 12155
rect 21508 12124 22477 12152
rect 21508 12112 21514 12124
rect 22465 12121 22477 12124
rect 22511 12121 22523 12155
rect 22465 12115 22523 12121
rect 17276 12056 19840 12084
rect 19889 12087 19947 12093
rect 17276 12044 17282 12056
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 20898 12084 20904 12096
rect 19935 12056 20904 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 21174 12044 21180 12096
rect 21232 12084 21238 12096
rect 22756 12084 22784 12192
rect 24118 12180 24124 12232
rect 24176 12220 24182 12232
rect 24578 12220 24584 12232
rect 24176 12192 24584 12220
rect 24176 12180 24182 12192
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 25976 12206 26004 12316
rect 27154 12248 27160 12300
rect 27212 12248 27218 12300
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 28353 12291 28411 12297
rect 28353 12288 28365 12291
rect 27396 12260 28365 12288
rect 27396 12248 27402 12260
rect 28353 12257 28365 12260
rect 28399 12288 28411 12291
rect 29733 12291 29791 12297
rect 29733 12288 29745 12291
rect 28399 12260 29745 12288
rect 28399 12257 28411 12260
rect 28353 12251 28411 12257
rect 29733 12257 29745 12260
rect 29779 12288 29791 12291
rect 30006 12288 30012 12300
rect 29779 12260 30012 12288
rect 29779 12257 29791 12260
rect 29733 12251 29791 12257
rect 30006 12248 30012 12260
rect 30064 12248 30070 12300
rect 31478 12288 31484 12300
rect 31128 12260 31484 12288
rect 31128 12232 31156 12260
rect 31478 12248 31484 12260
rect 31536 12288 31542 12300
rect 31757 12291 31815 12297
rect 31757 12288 31769 12291
rect 31536 12260 31769 12288
rect 31536 12248 31542 12260
rect 31757 12257 31769 12260
rect 31803 12257 31815 12291
rect 31757 12251 31815 12257
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 28810 12220 28816 12232
rect 27672 12192 28816 12220
rect 27672 12180 27678 12192
rect 28810 12180 28816 12192
rect 28868 12220 28874 12232
rect 29181 12223 29239 12229
rect 29181 12220 29193 12223
rect 28868 12192 29193 12220
rect 28868 12180 28874 12192
rect 29181 12189 29193 12192
rect 29227 12189 29239 12223
rect 29181 12183 29239 12189
rect 31110 12180 31116 12232
rect 31168 12180 31174 12232
rect 23661 12155 23719 12161
rect 23661 12152 23673 12155
rect 22848 12124 23673 12152
rect 22848 12093 22876 12124
rect 23661 12121 23673 12124
rect 23707 12121 23719 12155
rect 26878 12152 26884 12164
rect 23661 12115 23719 12121
rect 26160 12124 26884 12152
rect 21232 12056 22784 12084
rect 22833 12087 22891 12093
rect 21232 12044 21238 12056
rect 22833 12053 22845 12087
rect 22879 12053 22891 12087
rect 22833 12047 22891 12053
rect 23293 12087 23351 12093
rect 23293 12053 23305 12087
rect 23339 12084 23351 12087
rect 23382 12084 23388 12096
rect 23339 12056 23388 12084
rect 23339 12053 23351 12056
rect 23293 12047 23351 12053
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 23753 12087 23811 12093
rect 23753 12053 23765 12087
rect 23799 12084 23811 12087
rect 26160 12084 26188 12124
rect 26878 12112 26884 12124
rect 26936 12112 26942 12164
rect 27062 12112 27068 12164
rect 27120 12152 27126 12164
rect 27249 12155 27307 12161
rect 27249 12152 27261 12155
rect 27120 12124 27261 12152
rect 27120 12112 27126 12124
rect 27249 12121 27261 12124
rect 27295 12152 27307 12155
rect 27522 12152 27528 12164
rect 27295 12124 27528 12152
rect 27295 12121 27307 12124
rect 27249 12115 27307 12121
rect 27522 12112 27528 12124
rect 27580 12112 27586 12164
rect 29914 12112 29920 12164
rect 29972 12152 29978 12164
rect 30009 12155 30067 12161
rect 30009 12152 30021 12155
rect 29972 12124 30021 12152
rect 29972 12112 29978 12124
rect 30009 12121 30021 12124
rect 30055 12121 30067 12155
rect 30009 12115 30067 12121
rect 23799 12056 26188 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 27338 12044 27344 12096
rect 27396 12044 27402 12096
rect 31386 12044 31392 12096
rect 31444 12084 31450 12096
rect 31481 12087 31539 12093
rect 31481 12084 31493 12087
rect 31444 12056 31493 12084
rect 31444 12044 31450 12056
rect 31481 12053 31493 12056
rect 31527 12053 31539 12087
rect 31772 12084 31800 12251
rect 33870 12248 33876 12300
rect 33928 12288 33934 12300
rect 37185 12291 37243 12297
rect 37185 12288 37197 12291
rect 33928 12260 37197 12288
rect 33928 12248 33934 12260
rect 37185 12257 37197 12260
rect 37231 12257 37243 12291
rect 37185 12251 37243 12257
rect 38378 12248 38384 12300
rect 38436 12248 38442 12300
rect 38565 12291 38623 12297
rect 38565 12257 38577 12291
rect 38611 12288 38623 12291
rect 38746 12288 38752 12300
rect 38611 12260 38752 12288
rect 38611 12257 38623 12260
rect 38565 12251 38623 12257
rect 38746 12248 38752 12260
rect 38804 12248 38810 12300
rect 39040 12288 39068 12319
rect 39942 12316 39948 12328
rect 40000 12316 40006 12368
rect 40313 12359 40371 12365
rect 40313 12325 40325 12359
rect 40359 12356 40371 12359
rect 47394 12356 47400 12368
rect 40359 12328 47400 12356
rect 40359 12325 40371 12328
rect 40313 12319 40371 12325
rect 47394 12316 47400 12328
rect 47452 12316 47458 12368
rect 39040 12260 41460 12288
rect 32122 12180 32128 12232
rect 32180 12180 32186 12232
rect 34146 12180 34152 12232
rect 34204 12220 34210 12232
rect 34333 12223 34391 12229
rect 34333 12220 34345 12223
rect 34204 12192 34345 12220
rect 34204 12180 34210 12192
rect 34333 12189 34345 12192
rect 34379 12189 34391 12223
rect 34333 12183 34391 12189
rect 34882 12180 34888 12232
rect 34940 12180 34946 12232
rect 37090 12180 37096 12232
rect 37148 12220 37154 12232
rect 41432 12229 41460 12260
rect 49142 12248 49148 12300
rect 49200 12248 49206 12300
rect 37369 12223 37427 12229
rect 37369 12220 37381 12223
rect 37148 12192 37381 12220
rect 37148 12180 37154 12192
rect 37369 12189 37381 12192
rect 37415 12189 37427 12223
rect 40773 12223 40831 12229
rect 40773 12220 40785 12223
rect 37369 12183 37427 12189
rect 37844 12192 40785 12220
rect 32306 12112 32312 12164
rect 32364 12152 32370 12164
rect 32401 12155 32459 12161
rect 32401 12152 32413 12155
rect 32364 12124 32413 12152
rect 32364 12112 32370 12124
rect 32401 12121 32413 12124
rect 32447 12121 32459 12155
rect 32858 12152 32864 12164
rect 32401 12115 32459 12121
rect 32784 12124 32864 12152
rect 32784 12084 32812 12124
rect 32858 12112 32864 12124
rect 32916 12112 32922 12164
rect 34606 12112 34612 12164
rect 34664 12152 34670 12164
rect 35158 12152 35164 12164
rect 34664 12124 35164 12152
rect 34664 12112 34670 12124
rect 35158 12112 35164 12124
rect 35216 12112 35222 12164
rect 35268 12124 35650 12152
rect 34149 12087 34207 12093
rect 34149 12084 34161 12087
rect 31772 12056 34161 12084
rect 31481 12047 31539 12053
rect 34149 12053 34161 12056
rect 34195 12084 34207 12087
rect 34330 12084 34336 12096
rect 34195 12056 34336 12084
rect 34195 12053 34207 12056
rect 34149 12047 34207 12053
rect 34330 12044 34336 12056
rect 34388 12084 34394 12096
rect 35268 12084 35296 12124
rect 34388 12056 35296 12084
rect 34388 12044 34394 12056
rect 36538 12044 36544 12096
rect 36596 12084 36602 12096
rect 36633 12087 36691 12093
rect 36633 12084 36645 12087
rect 36596 12056 36645 12084
rect 36596 12044 36602 12056
rect 36633 12053 36645 12056
rect 36679 12084 36691 12087
rect 36722 12084 36728 12096
rect 36679 12056 36728 12084
rect 36679 12053 36691 12056
rect 36633 12047 36691 12053
rect 36722 12044 36728 12056
rect 36780 12044 36786 12096
rect 37274 12044 37280 12096
rect 37332 12084 37338 12096
rect 37844 12093 37872 12192
rect 40773 12189 40785 12192
rect 40819 12189 40831 12223
rect 40773 12183 40831 12189
rect 41417 12223 41475 12229
rect 41417 12189 41429 12223
rect 41463 12189 41475 12223
rect 45925 12223 45983 12229
rect 45925 12220 45937 12223
rect 41417 12183 41475 12189
rect 45526 12192 45937 12220
rect 40129 12155 40187 12161
rect 40129 12121 40141 12155
rect 40175 12152 40187 12155
rect 40402 12152 40408 12164
rect 40175 12124 40408 12152
rect 40175 12121 40187 12124
rect 40129 12115 40187 12121
rect 40402 12112 40408 12124
rect 40460 12112 40466 12164
rect 37461 12087 37519 12093
rect 37461 12084 37473 12087
rect 37332 12056 37473 12084
rect 37332 12044 37338 12056
rect 37461 12053 37473 12056
rect 37507 12053 37519 12087
rect 37461 12047 37519 12053
rect 37829 12087 37887 12093
rect 37829 12053 37841 12087
rect 37875 12053 37887 12087
rect 37829 12047 37887 12053
rect 38654 12044 38660 12096
rect 38712 12044 38718 12096
rect 40954 12044 40960 12096
rect 41012 12044 41018 12096
rect 41601 12087 41659 12093
rect 41601 12053 41613 12087
rect 41647 12084 41659 12087
rect 45526 12084 45554 12192
rect 45925 12189 45937 12192
rect 45971 12189 45983 12223
rect 45925 12183 45983 12189
rect 47946 12180 47952 12232
rect 48004 12180 48010 12232
rect 41647 12056 45554 12084
rect 41647 12053 41659 12056
rect 41601 12047 41659 12053
rect 46106 12044 46112 12096
rect 46164 12044 46170 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 2222 11840 2228 11892
rect 2280 11840 2286 11892
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 4246 11880 4252 11892
rect 4019 11852 4252 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 11609 11883 11667 11889
rect 11609 11849 11621 11883
rect 11655 11880 11667 11883
rect 11698 11880 11704 11892
rect 11655 11852 11704 11880
rect 11655 11849 11667 11852
rect 11609 11843 11667 11849
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12124 11852 12725 11880
rect 12124 11840 12130 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12713 11843 12771 11849
rect 13538 11840 13544 11892
rect 13596 11840 13602 11892
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 14185 11883 14243 11889
rect 14185 11880 14197 11883
rect 13688 11852 14197 11880
rect 13688 11840 13694 11852
rect 14185 11849 14197 11852
rect 14231 11849 14243 11883
rect 14185 11843 14243 11849
rect 14274 11840 14280 11892
rect 14332 11840 14338 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 16853 11883 16911 11889
rect 16853 11880 16865 11883
rect 14700 11852 16865 11880
rect 14700 11840 14706 11852
rect 16853 11849 16865 11852
rect 16899 11849 16911 11883
rect 16853 11843 16911 11849
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 19889 11883 19947 11889
rect 19889 11880 19901 11883
rect 18012 11852 19901 11880
rect 18012 11840 18018 11852
rect 19889 11849 19901 11852
rect 19935 11849 19947 11883
rect 19889 11843 19947 11849
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20257 11883 20315 11889
rect 20257 11880 20269 11883
rect 20036 11852 20269 11880
rect 20036 11840 20042 11852
rect 20257 11849 20269 11852
rect 20303 11849 20315 11883
rect 20257 11843 20315 11849
rect 20714 11840 20720 11892
rect 20772 11840 20778 11892
rect 21085 11883 21143 11889
rect 21085 11849 21097 11883
rect 21131 11880 21143 11883
rect 22002 11880 22008 11892
rect 21131 11852 22008 11880
rect 21131 11849 21143 11852
rect 21085 11843 21143 11849
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 22097 11883 22155 11889
rect 22097 11849 22109 11883
rect 22143 11880 22155 11883
rect 22370 11880 22376 11892
rect 22143 11852 22376 11880
rect 22143 11849 22155 11852
rect 22097 11843 22155 11849
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 12805 11815 12863 11821
rect 11296 11784 12434 11812
rect 11296 11772 11302 11784
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1360 11716 1593 11744
rect 1360 11704 1366 11716
rect 1581 11713 1593 11716
rect 1627 11744 1639 11747
rect 2314 11744 2320 11756
rect 1627 11716 2320 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 2682 11704 2688 11756
rect 2740 11704 2746 11756
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 3375 11716 3801 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 12406 11744 12434 11784
rect 12805 11781 12817 11815
rect 12851 11812 12863 11815
rect 14366 11812 14372 11824
rect 12851 11784 14372 11812
rect 12851 11781 12863 11784
rect 12805 11775 12863 11781
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 15378 11812 15384 11824
rect 14476 11784 15384 11812
rect 12986 11744 12992 11756
rect 12406 11716 12992 11744
rect 3789 11707 3847 11713
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 14476 11744 14504 11784
rect 15378 11772 15384 11784
rect 15436 11812 15442 11824
rect 15565 11815 15623 11821
rect 15565 11812 15577 11815
rect 15436 11784 15577 11812
rect 15436 11772 15442 11784
rect 15565 11781 15577 11784
rect 15611 11781 15623 11815
rect 15565 11775 15623 11781
rect 15764 11784 16528 11812
rect 13188 11716 14504 11744
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 11848 11648 12909 11676
rect 11848 11636 11854 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13188 11608 13216 11716
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 14792 11716 15485 11744
rect 14792 11704 14798 11716
rect 15473 11713 15485 11716
rect 15519 11744 15531 11747
rect 15764 11744 15792 11784
rect 16393 11747 16451 11753
rect 16393 11744 16405 11747
rect 15519 11716 15792 11744
rect 16040 11716 16405 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11676 14151 11679
rect 14274 11676 14280 11688
rect 14139 11648 14280 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 14608 11648 15608 11676
rect 14608 11636 14614 11648
rect 11992 11580 13216 11608
rect 14645 11611 14703 11617
rect 11882 11500 11888 11552
rect 11940 11540 11946 11552
rect 11992 11549 12020 11580
rect 14645 11577 14657 11611
rect 14691 11608 14703 11611
rect 15470 11608 15476 11620
rect 14691 11580 15476 11608
rect 14691 11577 14703 11580
rect 14645 11571 14703 11577
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 15580 11608 15608 11648
rect 15654 11636 15660 11688
rect 15712 11636 15718 11688
rect 16040 11608 16068 11716
rect 16393 11713 16405 11716
rect 16439 11713 16451 11747
rect 16393 11707 16451 11713
rect 15580 11580 16068 11608
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 11940 11512 11989 11540
rect 11940 11500 11946 11512
rect 11977 11509 11989 11512
rect 12023 11509 12035 11543
rect 11977 11503 12035 11509
rect 12342 11500 12348 11552
rect 12400 11500 12406 11552
rect 13354 11500 13360 11552
rect 13412 11500 13418 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14884 11512 15117 11540
rect 14884 11500 14890 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 16206 11540 16212 11552
rect 15436 11512 16212 11540
rect 15436 11500 15442 11512
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16408 11540 16436 11707
rect 16500 11676 16528 11784
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 18325 11815 18383 11821
rect 17000 11784 17158 11812
rect 17000 11772 17006 11784
rect 18325 11781 18337 11815
rect 18371 11812 18383 11815
rect 20438 11812 20444 11824
rect 18371 11784 20444 11812
rect 18371 11781 18383 11784
rect 18325 11775 18383 11781
rect 20438 11772 20444 11784
rect 20496 11772 20502 11824
rect 20530 11772 20536 11824
rect 20588 11812 20594 11824
rect 22112 11812 22140 11843
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 24486 11840 24492 11892
rect 24544 11880 24550 11892
rect 25685 11883 25743 11889
rect 25685 11880 25697 11883
rect 24544 11852 25697 11880
rect 24544 11840 24550 11852
rect 25685 11849 25697 11852
rect 25731 11849 25743 11883
rect 25685 11843 25743 11849
rect 26605 11883 26663 11889
rect 26605 11849 26617 11883
rect 26651 11880 26663 11883
rect 27338 11880 27344 11892
rect 26651 11852 27344 11880
rect 26651 11849 26663 11852
rect 26605 11843 26663 11849
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 27893 11883 27951 11889
rect 27893 11849 27905 11883
rect 27939 11880 27951 11883
rect 28626 11880 28632 11892
rect 27939 11852 28632 11880
rect 27939 11849 27951 11852
rect 27893 11843 27951 11849
rect 28626 11840 28632 11852
rect 28684 11840 28690 11892
rect 31110 11880 31116 11892
rect 28736 11852 31116 11880
rect 20588 11784 22140 11812
rect 20588 11772 20594 11784
rect 22186 11772 22192 11824
rect 22244 11812 22250 11824
rect 23385 11815 23443 11821
rect 23385 11812 23397 11815
rect 22244 11784 23397 11812
rect 22244 11772 22250 11784
rect 23385 11781 23397 11784
rect 23431 11812 23443 11815
rect 24118 11812 24124 11824
rect 23431 11784 24124 11812
rect 23431 11781 23443 11784
rect 23385 11775 23443 11781
rect 18690 11704 18696 11756
rect 18748 11744 18754 11756
rect 19794 11744 19800 11756
rect 18748 11716 19800 11744
rect 18748 11704 18754 11716
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 20806 11744 20812 11756
rect 20180 11716 20812 11744
rect 18601 11679 18659 11685
rect 16500 11648 18552 11676
rect 18524 11608 18552 11648
rect 18601 11645 18613 11679
rect 18647 11676 18659 11679
rect 18782 11676 18788 11688
rect 18647 11648 18788 11676
rect 18647 11645 18659 11648
rect 18601 11639 18659 11645
rect 18782 11636 18788 11648
rect 18840 11636 18846 11688
rect 19058 11636 19064 11688
rect 19116 11636 19122 11688
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11676 19763 11679
rect 20180 11676 20208 11716
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 22462 11704 22468 11756
rect 22520 11744 22526 11756
rect 23952 11753 23980 11784
rect 24118 11772 24124 11784
rect 24176 11772 24182 11824
rect 25590 11772 25596 11824
rect 25648 11812 25654 11824
rect 26145 11815 26203 11821
rect 26145 11812 26157 11815
rect 25648 11784 26157 11812
rect 25648 11772 25654 11784
rect 26145 11781 26157 11784
rect 26191 11812 26203 11815
rect 26970 11812 26976 11824
rect 26191 11784 26976 11812
rect 26191 11781 26203 11784
rect 26145 11775 26203 11781
rect 26970 11772 26976 11784
rect 27028 11812 27034 11824
rect 27525 11815 27583 11821
rect 27525 11812 27537 11815
rect 27028 11784 27537 11812
rect 27028 11772 27034 11784
rect 27525 11781 27537 11784
rect 27571 11781 27583 11815
rect 27525 11775 27583 11781
rect 28442 11772 28448 11824
rect 28500 11812 28506 11824
rect 28736 11812 28764 11852
rect 31110 11840 31116 11852
rect 31168 11840 31174 11892
rect 31481 11883 31539 11889
rect 31481 11849 31493 11883
rect 31527 11880 31539 11883
rect 31846 11880 31852 11892
rect 31527 11852 31852 11880
rect 31527 11849 31539 11852
rect 31481 11843 31539 11849
rect 31846 11840 31852 11852
rect 31904 11840 31910 11892
rect 32398 11840 32404 11892
rect 32456 11880 32462 11892
rect 32585 11883 32643 11889
rect 32585 11880 32597 11883
rect 32456 11852 32597 11880
rect 32456 11840 32462 11852
rect 32585 11849 32597 11852
rect 32631 11849 32643 11883
rect 32585 11843 32643 11849
rect 32674 11840 32680 11892
rect 32732 11840 32738 11892
rect 33045 11883 33103 11889
rect 33045 11849 33057 11883
rect 33091 11849 33103 11883
rect 33045 11843 33103 11849
rect 30009 11815 30067 11821
rect 28500 11784 28842 11812
rect 28500 11772 28506 11784
rect 22557 11747 22615 11753
rect 22557 11744 22569 11747
rect 22520 11716 22569 11744
rect 22520 11704 22526 11716
rect 22557 11713 22569 11716
rect 22603 11713 22615 11747
rect 22557 11707 22615 11713
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11713 23995 11747
rect 25682 11744 25688 11756
rect 25346 11716 25688 11744
rect 23937 11707 23995 11713
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 25774 11704 25780 11756
rect 25832 11744 25838 11756
rect 25832 11716 27476 11744
rect 25832 11704 25838 11716
rect 27448 11688 27476 11716
rect 19751 11648 20208 11676
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 20346 11636 20352 11688
rect 20404 11676 20410 11688
rect 21174 11676 21180 11688
rect 20404 11648 21180 11676
rect 20404 11636 20410 11648
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 21361 11679 21419 11685
rect 21361 11645 21373 11679
rect 21407 11676 21419 11679
rect 21542 11676 21548 11688
rect 21407 11648 21548 11676
rect 21407 11645 21419 11648
rect 21361 11639 21419 11645
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 23474 11636 23480 11688
rect 23532 11676 23538 11688
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 23532 11648 24225 11676
rect 23532 11636 23538 11648
rect 24213 11645 24225 11648
rect 24259 11676 24271 11679
rect 26326 11676 26332 11688
rect 24259 11648 26332 11676
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 27341 11679 27399 11685
rect 27341 11645 27353 11679
rect 27387 11645 27399 11679
rect 27341 11639 27399 11645
rect 26142 11608 26148 11620
rect 18524 11580 18828 11608
rect 18690 11540 18696 11552
rect 16408 11512 18696 11540
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 18800 11540 18828 11580
rect 18984 11580 19288 11608
rect 18984 11540 19012 11580
rect 18800 11512 19012 11540
rect 19150 11500 19156 11552
rect 19208 11500 19214 11552
rect 19260 11540 19288 11580
rect 21192 11580 24072 11608
rect 21192 11540 21220 11580
rect 19260 11512 21220 11540
rect 21266 11500 21272 11552
rect 21324 11540 21330 11552
rect 21634 11540 21640 11552
rect 21324 11512 21640 11540
rect 21324 11500 21330 11512
rect 21634 11500 21640 11512
rect 21692 11540 21698 11552
rect 21821 11543 21879 11549
rect 21821 11540 21833 11543
rect 21692 11512 21833 11540
rect 21692 11500 21698 11512
rect 21821 11509 21833 11512
rect 21867 11540 21879 11543
rect 22002 11540 22008 11552
rect 21867 11512 22008 11540
rect 21867 11509 21879 11512
rect 21821 11503 21879 11509
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 22281 11543 22339 11549
rect 22281 11509 22293 11543
rect 22327 11540 22339 11543
rect 22462 11540 22468 11552
rect 22327 11512 22468 11540
rect 22327 11509 22339 11512
rect 22281 11503 22339 11509
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 24044 11540 24072 11580
rect 25240 11580 26148 11608
rect 24670 11540 24676 11552
rect 24044 11512 24676 11540
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 24762 11500 24768 11552
rect 24820 11540 24826 11552
rect 25240 11540 25268 11580
rect 26142 11568 26148 11580
rect 26200 11568 26206 11620
rect 27356 11608 27384 11639
rect 27430 11636 27436 11688
rect 27488 11636 27494 11688
rect 27798 11608 27804 11620
rect 27356 11580 27804 11608
rect 27798 11568 27804 11580
rect 27856 11568 27862 11620
rect 28736 11608 28764 11784
rect 30009 11781 30021 11815
rect 30055 11812 30067 11815
rect 31386 11812 31392 11824
rect 30055 11784 31392 11812
rect 30055 11781 30067 11784
rect 30009 11775 30067 11781
rect 31386 11772 31392 11784
rect 31444 11812 31450 11824
rect 33060 11812 33088 11843
rect 33778 11840 33784 11892
rect 33836 11880 33842 11892
rect 33873 11883 33931 11889
rect 33873 11880 33885 11883
rect 33836 11852 33885 11880
rect 33836 11840 33842 11852
rect 33873 11849 33885 11852
rect 33919 11849 33931 11883
rect 33873 11843 33931 11849
rect 34330 11840 34336 11892
rect 34388 11880 34394 11892
rect 34701 11883 34759 11889
rect 34701 11880 34713 11883
rect 34388 11852 34713 11880
rect 34388 11840 34394 11852
rect 34701 11849 34713 11852
rect 34747 11880 34759 11883
rect 34747 11852 35204 11880
rect 34747 11849 34759 11852
rect 34701 11843 34759 11849
rect 35066 11812 35072 11824
rect 31444 11784 31754 11812
rect 33060 11784 35072 11812
rect 31444 11772 31450 11784
rect 31110 11704 31116 11756
rect 31168 11704 31174 11756
rect 31726 11744 31754 11784
rect 35066 11772 35072 11784
rect 35124 11772 35130 11824
rect 35176 11812 35204 11852
rect 35250 11840 35256 11892
rect 35308 11880 35314 11892
rect 37737 11883 37795 11889
rect 37737 11880 37749 11883
rect 35308 11852 37749 11880
rect 35308 11840 35314 11852
rect 37737 11849 37749 11852
rect 37783 11849 37795 11883
rect 37737 11843 37795 11849
rect 38654 11840 38660 11892
rect 38712 11840 38718 11892
rect 39114 11840 39120 11892
rect 39172 11840 39178 11892
rect 35710 11812 35716 11824
rect 35176 11784 35716 11812
rect 35710 11772 35716 11784
rect 35768 11812 35774 11824
rect 35768 11784 35926 11812
rect 35768 11772 35774 11784
rect 36722 11772 36728 11824
rect 36780 11812 36786 11824
rect 36780 11784 39252 11812
rect 36780 11772 36786 11784
rect 31726 11716 32996 11744
rect 28810 11636 28816 11688
rect 28868 11676 28874 11688
rect 28868 11648 30236 11676
rect 28868 11636 28874 11648
rect 28902 11608 28908 11620
rect 28736 11580 28908 11608
rect 28902 11568 28908 11580
rect 28960 11568 28966 11620
rect 30208 11608 30236 11648
rect 30282 11636 30288 11688
rect 30340 11636 30346 11688
rect 30834 11636 30840 11688
rect 30892 11636 30898 11688
rect 31021 11679 31079 11685
rect 31021 11645 31033 11679
rect 31067 11676 31079 11679
rect 31754 11676 31760 11688
rect 31067 11648 31760 11676
rect 31067 11645 31079 11648
rect 31021 11639 31079 11645
rect 31754 11636 31760 11648
rect 31812 11636 31818 11688
rect 32493 11679 32551 11685
rect 32493 11645 32505 11679
rect 32539 11676 32551 11679
rect 32858 11676 32864 11688
rect 32539 11648 32864 11676
rect 32539 11645 32551 11648
rect 32493 11639 32551 11645
rect 32858 11636 32864 11648
rect 32916 11636 32922 11688
rect 32968 11676 32996 11716
rect 33686 11704 33692 11756
rect 33744 11744 33750 11756
rect 33781 11747 33839 11753
rect 33781 11744 33793 11747
rect 33744 11716 33793 11744
rect 33744 11704 33750 11716
rect 33781 11713 33793 11716
rect 33827 11713 33839 11747
rect 33781 11707 33839 11713
rect 36814 11704 36820 11756
rect 36872 11744 36878 11756
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 36872 11716 37841 11744
rect 36872 11704 36878 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 39022 11704 39028 11756
rect 39080 11704 39086 11756
rect 33597 11679 33655 11685
rect 33597 11676 33609 11679
rect 32968 11648 33609 11676
rect 33597 11645 33609 11648
rect 33643 11645 33655 11679
rect 33597 11639 33655 11645
rect 33962 11636 33968 11688
rect 34020 11676 34026 11688
rect 34238 11676 34244 11688
rect 34020 11648 34244 11676
rect 34020 11636 34026 11648
rect 34238 11636 34244 11648
rect 34296 11636 34302 11688
rect 34882 11636 34888 11688
rect 34940 11676 34946 11688
rect 35161 11679 35219 11685
rect 35161 11676 35173 11679
rect 34940 11648 35173 11676
rect 34940 11636 34946 11648
rect 35161 11645 35173 11648
rect 35207 11645 35219 11679
rect 35161 11639 35219 11645
rect 35437 11679 35495 11685
rect 35437 11645 35449 11679
rect 35483 11676 35495 11679
rect 36446 11676 36452 11688
rect 35483 11648 36452 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 31386 11608 31392 11620
rect 30208 11580 31392 11608
rect 31386 11568 31392 11580
rect 31444 11568 31450 11620
rect 24820 11512 25268 11540
rect 24820 11500 24826 11512
rect 27246 11500 27252 11552
rect 27304 11540 27310 11552
rect 28537 11543 28595 11549
rect 28537 11540 28549 11543
rect 27304 11512 28549 11540
rect 27304 11500 27310 11512
rect 28537 11509 28549 11512
rect 28583 11540 28595 11543
rect 30190 11540 30196 11552
rect 28583 11512 30196 11540
rect 28583 11509 28595 11512
rect 28537 11503 28595 11509
rect 30190 11500 30196 11512
rect 30248 11500 30254 11552
rect 31478 11500 31484 11552
rect 31536 11540 31542 11552
rect 31757 11543 31815 11549
rect 31757 11540 31769 11543
rect 31536 11512 31769 11540
rect 31536 11500 31542 11512
rect 31757 11509 31769 11512
rect 31803 11509 31815 11543
rect 31757 11503 31815 11509
rect 34238 11500 34244 11552
rect 34296 11500 34302 11552
rect 34422 11500 34428 11552
rect 34480 11540 34486 11552
rect 34517 11543 34575 11549
rect 34517 11540 34529 11543
rect 34480 11512 34529 11540
rect 34480 11500 34486 11512
rect 34517 11509 34529 11512
rect 34563 11509 34575 11543
rect 35176 11540 35204 11639
rect 36446 11636 36452 11648
rect 36504 11636 36510 11688
rect 36630 11636 36636 11688
rect 36688 11676 36694 11688
rect 39224 11685 39252 11784
rect 39942 11772 39948 11824
rect 40000 11772 40006 11824
rect 40402 11772 40408 11824
rect 40460 11772 40466 11824
rect 40954 11772 40960 11824
rect 41012 11812 41018 11824
rect 45097 11815 45155 11821
rect 45097 11812 45109 11815
rect 41012 11784 45109 11812
rect 41012 11772 41018 11784
rect 45097 11781 45109 11784
rect 45143 11781 45155 11815
rect 45097 11775 45155 11781
rect 49142 11772 49148 11824
rect 49200 11772 49206 11824
rect 39960 11744 39988 11772
rect 40589 11747 40647 11753
rect 40589 11744 40601 11747
rect 39960 11716 40601 11744
rect 40589 11713 40601 11716
rect 40635 11713 40647 11747
rect 40589 11707 40647 11713
rect 46106 11704 46112 11756
rect 46164 11744 46170 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 46164 11716 47961 11744
rect 46164 11704 46170 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 37553 11679 37611 11685
rect 37553 11676 37565 11679
rect 36688 11648 37565 11676
rect 36688 11636 36694 11648
rect 37553 11645 37565 11648
rect 37599 11645 37611 11679
rect 37553 11639 37611 11645
rect 39209 11679 39267 11685
rect 39209 11645 39221 11679
rect 39255 11645 39267 11679
rect 39209 11639 39267 11645
rect 36909 11611 36967 11617
rect 36909 11577 36921 11611
rect 36955 11608 36967 11611
rect 38378 11608 38384 11620
rect 36955 11580 38384 11608
rect 36955 11577 36967 11580
rect 36909 11571 36967 11577
rect 38378 11568 38384 11580
rect 38436 11568 38442 11620
rect 40129 11611 40187 11617
rect 40129 11577 40141 11611
rect 40175 11608 40187 11611
rect 45281 11611 45339 11617
rect 40175 11580 42840 11608
rect 40175 11577 40187 11580
rect 40129 11571 40187 11577
rect 35618 11540 35624 11552
rect 35176 11512 35624 11540
rect 34517 11503 34575 11509
rect 35618 11500 35624 11512
rect 35676 11500 35682 11552
rect 38197 11543 38255 11549
rect 38197 11509 38209 11543
rect 38243 11540 38255 11543
rect 40218 11540 40224 11552
rect 38243 11512 40224 11540
rect 38243 11509 38255 11512
rect 38197 11503 38255 11509
rect 40218 11500 40224 11512
rect 40276 11500 40282 11552
rect 42812 11540 42840 11580
rect 45281 11577 45293 11611
rect 45327 11608 45339 11611
rect 46658 11608 46664 11620
rect 45327 11580 46664 11608
rect 45327 11577 45339 11580
rect 45281 11571 45339 11577
rect 46658 11568 46664 11580
rect 46716 11568 46722 11620
rect 47026 11540 47032 11552
rect 42812 11512 47032 11540
rect 47026 11500 47032 11512
rect 47084 11500 47090 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 11422 11336 11428 11348
rect 2915 11308 11428 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 13265 11339 13323 11345
rect 12492 11308 13124 11336
rect 12492 11296 12498 11308
rect 1302 11228 1308 11280
rect 1360 11268 1366 11280
rect 2682 11268 2688 11280
rect 1360 11240 2688 11268
rect 1360 11228 1366 11240
rect 2682 11228 2688 11240
rect 2740 11268 2746 11280
rect 3237 11271 3295 11277
rect 3237 11268 3249 11271
rect 2740 11240 3249 11268
rect 2740 11228 2746 11240
rect 3237 11237 3249 11240
rect 3283 11237 3295 11271
rect 3237 11231 3295 11237
rect 4157 11271 4215 11277
rect 4157 11237 4169 11271
rect 4203 11268 4215 11271
rect 11238 11268 11244 11280
rect 4203 11240 11244 11268
rect 4203 11237 4215 11240
rect 4157 11231 4215 11237
rect 11238 11228 11244 11240
rect 11296 11228 11302 11280
rect 3421 11203 3479 11209
rect 3421 11200 3433 11203
rect 1596 11172 3433 11200
rect 1210 11092 1216 11144
rect 1268 11132 1274 11144
rect 1596 11141 1624 11172
rect 3421 11169 3433 11172
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11054 11200 11060 11212
rect 11011 11172 11060 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11790 11160 11796 11212
rect 11848 11200 11854 11212
rect 13096 11209 13124 11308
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13538 11336 13544 11348
rect 13311 11308 13544 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 13964 11308 14381 11336
rect 13964 11296 13970 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 15562 11336 15568 11348
rect 14516 11308 15568 11336
rect 14516 11296 14522 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16724 11308 16773 11336
rect 16724 11296 16730 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 16761 11299 16819 11305
rect 18874 11296 18880 11348
rect 18932 11336 18938 11348
rect 19061 11339 19119 11345
rect 19061 11336 19073 11339
rect 18932 11308 19073 11336
rect 18932 11296 18938 11308
rect 19061 11305 19073 11308
rect 19107 11336 19119 11339
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 19107 11308 19349 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19337 11305 19349 11308
rect 19383 11336 19395 11339
rect 22462 11336 22468 11348
rect 19383 11308 22468 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 23290 11296 23296 11348
rect 23348 11296 23354 11348
rect 25222 11336 25228 11348
rect 24412 11308 25228 11336
rect 16301 11271 16359 11277
rect 16301 11237 16313 11271
rect 16347 11268 16359 11271
rect 18414 11268 18420 11280
rect 16347 11240 18420 11268
rect 16347 11237 16359 11240
rect 16301 11231 16359 11237
rect 18414 11228 18420 11240
rect 18472 11228 18478 11280
rect 19150 11268 19156 11280
rect 18524 11240 19156 11268
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 11848 11172 12449 11200
rect 11848 11160 11854 11172
rect 12437 11169 12449 11172
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11200 13139 11203
rect 14734 11200 14740 11212
rect 13127 11172 14740 11200
rect 13127 11169 13139 11172
rect 13081 11163 13139 11169
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11200 15071 11203
rect 15102 11200 15108 11212
rect 15059 11172 15108 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 15746 11160 15752 11212
rect 15804 11160 15810 11212
rect 15838 11160 15844 11212
rect 15896 11160 15902 11212
rect 17402 11160 17408 11212
rect 17460 11160 17466 11212
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 18524 11200 18552 11240
rect 19150 11228 19156 11240
rect 19208 11268 19214 11280
rect 19521 11271 19579 11277
rect 19521 11268 19533 11271
rect 19208 11240 19533 11268
rect 19208 11228 19214 11240
rect 19521 11237 19533 11240
rect 19567 11268 19579 11271
rect 20346 11268 20352 11280
rect 19567 11240 20352 11268
rect 19567 11237 19579 11240
rect 19521 11231 19579 11237
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 20438 11228 20444 11280
rect 20496 11228 20502 11280
rect 17736 11172 18552 11200
rect 18601 11203 18659 11209
rect 17736 11160 17742 11172
rect 18601 11169 18613 11203
rect 18647 11200 18659 11203
rect 19426 11200 19432 11212
rect 18647 11172 19432 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 19981 11203 20039 11209
rect 19981 11169 19993 11203
rect 20027 11200 20039 11203
rect 20070 11200 20076 11212
rect 20027 11172 20076 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 23750 11200 23756 11212
rect 20640 11172 23756 11200
rect 1581 11135 1639 11141
rect 1581 11132 1593 11135
rect 1268 11104 1593 11132
rect 1268 11092 1274 11104
rect 1581 11101 1593 11104
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2271 11104 2697 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 2832 11104 3985 11132
rect 2832 11092 2838 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 12710 11092 12716 11144
rect 12768 11092 12774 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16850 11132 16856 11144
rect 15979 11104 16856 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 19058 11132 19064 11144
rect 17175 11104 19064 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 20640 11132 20668 11172
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11200 23995 11203
rect 24412 11200 24440 11308
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 26602 11336 26608 11348
rect 26375 11308 26608 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 28534 11296 28540 11348
rect 28592 11336 28598 11348
rect 28629 11339 28687 11345
rect 28629 11336 28641 11339
rect 28592 11308 28641 11336
rect 28592 11296 28598 11308
rect 28629 11305 28641 11308
rect 28675 11305 28687 11339
rect 28629 11299 28687 11305
rect 28810 11296 28816 11348
rect 28868 11336 28874 11348
rect 28997 11339 29055 11345
rect 28997 11336 29009 11339
rect 28868 11308 29009 11336
rect 28868 11296 28874 11308
rect 28997 11305 29009 11308
rect 29043 11305 29055 11339
rect 28997 11299 29055 11305
rect 30466 11296 30472 11348
rect 30524 11296 30530 11348
rect 31386 11296 31392 11348
rect 31444 11336 31450 11348
rect 33318 11336 33324 11348
rect 31444 11308 33324 11336
rect 31444 11296 31450 11308
rect 33318 11296 33324 11308
rect 33376 11336 33382 11348
rect 34422 11336 34428 11348
rect 33376 11308 34428 11336
rect 33376 11296 33382 11308
rect 34422 11296 34428 11308
rect 34480 11336 34486 11348
rect 34701 11339 34759 11345
rect 34701 11336 34713 11339
rect 34480 11308 34713 11336
rect 34480 11296 34486 11308
rect 34701 11305 34713 11308
rect 34747 11305 34759 11339
rect 34701 11299 34759 11305
rect 36464 11308 38240 11336
rect 31018 11268 31024 11280
rect 29840 11240 31024 11268
rect 23983 11172 24440 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24486 11160 24492 11212
rect 24544 11200 24550 11212
rect 24857 11203 24915 11209
rect 24857 11200 24869 11203
rect 24544 11172 24869 11200
rect 24544 11160 24550 11172
rect 24857 11169 24869 11172
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 19306 11104 20668 11132
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13725 11067 13783 11073
rect 13725 11064 13737 11067
rect 13504 11036 13737 11064
rect 13504 11024 13510 11036
rect 13725 11033 13737 11036
rect 13771 11033 13783 11067
rect 13725 11027 13783 11033
rect 14734 11024 14740 11076
rect 14792 11064 14798 11076
rect 16666 11064 16672 11076
rect 14792 11036 16672 11064
rect 14792 11024 14798 11036
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 18325 11067 18383 11073
rect 18325 11033 18337 11067
rect 18371 11064 18383 11067
rect 18506 11064 18512 11076
rect 18371 11036 18512 11064
rect 18371 11033 18383 11036
rect 18325 11027 18383 11033
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 18782 11064 18788 11076
rect 18616 11036 18788 11064
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 12526 10996 12532 11008
rect 11756 10968 12532 10996
rect 11756 10956 11762 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 17126 10996 17132 11008
rect 15344 10968 17132 10996
rect 15344 10956 15350 10968
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17218 10956 17224 11008
rect 17276 10956 17282 11008
rect 17310 10956 17316 11008
rect 17368 10996 17374 11008
rect 17957 10999 18015 11005
rect 17957 10996 17969 10999
rect 17368 10968 17969 10996
rect 17368 10956 17374 10968
rect 17957 10965 17969 10968
rect 18003 10965 18015 10999
rect 17957 10959 18015 10965
rect 18417 10999 18475 11005
rect 18417 10965 18429 10999
rect 18463 10996 18475 10999
rect 18616 10996 18644 11036
rect 18782 11024 18788 11036
rect 18840 11064 18846 11076
rect 19306 11064 19334 11104
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 24578 11092 24584 11144
rect 24636 11092 24642 11144
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 29362 11092 29368 11144
rect 29420 11132 29426 11144
rect 29840 11132 29868 11240
rect 31018 11228 31024 11240
rect 31076 11228 31082 11280
rect 32858 11228 32864 11280
rect 32916 11228 32922 11280
rect 34238 11228 34244 11280
rect 34296 11268 34302 11280
rect 36464 11268 36492 11308
rect 34296 11240 36492 11268
rect 34296 11228 34302 11240
rect 29917 11203 29975 11209
rect 29917 11169 29929 11203
rect 29963 11200 29975 11203
rect 30190 11200 30196 11212
rect 29963 11172 30196 11200
rect 29963 11169 29975 11172
rect 29917 11163 29975 11169
rect 30190 11160 30196 11172
rect 30248 11160 30254 11212
rect 32122 11160 32128 11212
rect 32180 11200 32186 11212
rect 34057 11203 34115 11209
rect 34057 11200 34069 11203
rect 32180 11172 34069 11200
rect 32180 11160 32186 11172
rect 34057 11169 34069 11172
rect 34103 11169 34115 11203
rect 34057 11163 34115 11169
rect 35710 11160 35716 11212
rect 35768 11200 35774 11212
rect 35768 11172 36400 11200
rect 35768 11160 35774 11172
rect 30009 11135 30067 11141
rect 30009 11132 30021 11135
rect 29420 11104 30021 11132
rect 29420 11092 29426 11104
rect 30009 11101 30021 11104
rect 30055 11101 30067 11135
rect 30009 11095 30067 11101
rect 30282 11092 30288 11144
rect 30340 11132 30346 11144
rect 31113 11135 31171 11141
rect 31113 11132 31125 11135
rect 30340 11104 31125 11132
rect 30340 11092 30346 11104
rect 31113 11101 31125 11104
rect 31159 11101 31171 11135
rect 31113 11095 31171 11101
rect 33318 11092 33324 11144
rect 33376 11092 33382 11144
rect 36372 11118 36400 11172
rect 37458 11160 37464 11212
rect 37516 11200 37522 11212
rect 37737 11203 37795 11209
rect 37737 11200 37749 11203
rect 37516 11172 37749 11200
rect 37516 11160 37522 11172
rect 37737 11169 37749 11172
rect 37783 11169 37795 11203
rect 37737 11163 37795 11169
rect 38212 11141 38240 11308
rect 38654 11296 38660 11348
rect 38712 11336 38718 11348
rect 38749 11339 38807 11345
rect 38749 11336 38761 11339
rect 38712 11308 38761 11336
rect 38712 11296 38718 11308
rect 38749 11305 38761 11308
rect 38795 11336 38807 11339
rect 39482 11336 39488 11348
rect 38795 11308 39488 11336
rect 38795 11305 38807 11308
rect 38749 11299 38807 11305
rect 39482 11296 39488 11308
rect 39540 11296 39546 11348
rect 39574 11296 39580 11348
rect 39632 11296 39638 11348
rect 44358 11336 44364 11348
rect 39868 11308 44364 11336
rect 38381 11271 38439 11277
rect 38381 11237 38393 11271
rect 38427 11268 38439 11271
rect 39868 11268 39896 11308
rect 44358 11296 44364 11308
rect 44416 11296 44422 11348
rect 38427 11240 39896 11268
rect 40957 11271 41015 11277
rect 38427 11237 38439 11240
rect 38381 11231 38439 11237
rect 40957 11237 40969 11271
rect 41003 11268 41015 11271
rect 41003 11240 45554 11268
rect 41003 11237 41015 11240
rect 40957 11231 41015 11237
rect 38197 11135 38255 11141
rect 38197 11101 38209 11135
rect 38243 11101 38255 11135
rect 38197 11095 38255 11101
rect 39574 11092 39580 11144
rect 39632 11132 39638 11144
rect 40129 11135 40187 11141
rect 40129 11132 40141 11135
rect 39632 11104 40141 11132
rect 39632 11092 39638 11104
rect 40129 11101 40141 11104
rect 40175 11101 40187 11135
rect 40129 11095 40187 11101
rect 40218 11092 40224 11144
rect 40276 11132 40282 11144
rect 40773 11135 40831 11141
rect 40773 11132 40785 11135
rect 40276 11104 40785 11132
rect 40276 11092 40282 11104
rect 40773 11101 40785 11104
rect 40819 11101 40831 11135
rect 45526 11132 45554 11240
rect 49142 11160 49148 11212
rect 49200 11160 49206 11212
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 45526 11104 45661 11132
rect 40773 11095 40831 11101
rect 45649 11101 45661 11104
rect 45695 11101 45707 11135
rect 45649 11095 45707 11101
rect 46934 11092 46940 11144
rect 46992 11132 46998 11144
rect 47949 11135 48007 11141
rect 47949 11132 47961 11135
rect 46992 11104 47961 11132
rect 46992 11092 46998 11104
rect 47949 11101 47961 11104
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 18840 11036 19334 11064
rect 18840 11024 18846 11036
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 20438 11064 20444 11076
rect 20220 11036 20444 11064
rect 20220 11024 20226 11036
rect 20438 11024 20444 11036
rect 20496 11064 20502 11076
rect 21913 11067 21971 11073
rect 20496 11036 20746 11064
rect 20496 11024 20502 11036
rect 21913 11033 21925 11067
rect 21959 11064 21971 11067
rect 23566 11064 23572 11076
rect 21959 11036 23572 11064
rect 21959 11033 21971 11036
rect 21913 11027 21971 11033
rect 23566 11024 23572 11036
rect 23624 11024 23630 11076
rect 23661 11067 23719 11073
rect 23661 11033 23673 11067
rect 23707 11064 23719 11067
rect 23934 11064 23940 11076
rect 23707 11036 23940 11064
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 26694 11064 26700 11076
rect 26082 11036 26700 11064
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 27154 11024 27160 11076
rect 27212 11024 27218 11076
rect 28534 11064 28540 11076
rect 28382 11036 28540 11064
rect 28534 11024 28540 11036
rect 28592 11064 28598 11076
rect 28902 11064 28908 11076
rect 28592 11036 28908 11064
rect 28592 11024 28598 11036
rect 28902 11024 28908 11036
rect 28960 11024 28966 11076
rect 29454 11024 29460 11076
rect 29512 11064 29518 11076
rect 30101 11067 30159 11073
rect 30101 11064 30113 11067
rect 29512 11036 30113 11064
rect 29512 11024 29518 11036
rect 30101 11033 30113 11036
rect 30147 11033 30159 11067
rect 30101 11027 30159 11033
rect 18463 10968 18644 10996
rect 18463 10965 18475 10968
rect 18417 10959 18475 10965
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 25590 10996 25596 11008
rect 19852 10968 25596 10996
rect 19852 10956 19858 10968
rect 25590 10956 25596 10968
rect 25648 10956 25654 11008
rect 28994 10956 29000 11008
rect 29052 10996 29058 11008
rect 29089 10999 29147 11005
rect 29089 10996 29101 10999
rect 29052 10968 29101 10996
rect 29052 10956 29058 10968
rect 29089 10965 29101 10968
rect 29135 10996 29147 10999
rect 29273 10999 29331 11005
rect 29273 10996 29285 10999
rect 29135 10968 29285 10996
rect 29135 10965 29147 10968
rect 29089 10959 29147 10965
rect 29273 10965 29285 10968
rect 29319 10965 29331 10999
rect 30116 10996 30144 11027
rect 30374 11024 30380 11076
rect 30432 11064 30438 11076
rect 31294 11064 31300 11076
rect 30432 11036 31300 11064
rect 30432 11024 30438 11036
rect 31294 11024 31300 11036
rect 31352 11064 31358 11076
rect 31389 11067 31447 11073
rect 31389 11064 31401 11067
rect 31352 11036 31401 11064
rect 31352 11024 31358 11036
rect 31389 11033 31401 11036
rect 31435 11033 31447 11067
rect 31389 11027 31447 11033
rect 31478 11024 31484 11076
rect 31536 11064 31542 11076
rect 34790 11064 34796 11076
rect 31536 11036 31878 11064
rect 33704 11036 34796 11064
rect 31536 11024 31542 11036
rect 30745 10999 30803 11005
rect 30745 10996 30757 10999
rect 30116 10968 30757 10996
rect 29273 10959 29331 10965
rect 30745 10965 30757 10968
rect 30791 10996 30803 10999
rect 30834 10996 30840 11008
rect 30791 10968 30840 10996
rect 30791 10965 30803 10968
rect 30745 10959 30803 10965
rect 30834 10956 30840 10968
rect 30892 10956 30898 11008
rect 31570 10956 31576 11008
rect 31628 10996 31634 11008
rect 33704 10996 33732 11036
rect 34790 11024 34796 11036
rect 34848 11024 34854 11076
rect 35526 11024 35532 11076
rect 35584 11064 35590 11076
rect 35713 11067 35771 11073
rect 35713 11064 35725 11067
rect 35584 11036 35725 11064
rect 35584 11024 35590 11036
rect 35713 11033 35725 11036
rect 35759 11064 35771 11067
rect 35894 11064 35900 11076
rect 35759 11036 35900 11064
rect 35759 11033 35771 11036
rect 35713 11027 35771 11033
rect 35894 11024 35900 11036
rect 35952 11024 35958 11076
rect 37461 11067 37519 11073
rect 37461 11033 37473 11067
rect 37507 11064 37519 11067
rect 38378 11064 38384 11076
rect 37507 11036 38384 11064
rect 37507 11033 37519 11036
rect 37461 11027 37519 11033
rect 38378 11024 38384 11036
rect 38436 11024 38442 11076
rect 40313 11067 40371 11073
rect 40313 11033 40325 11067
rect 40359 11064 40371 11067
rect 45833 11067 45891 11073
rect 40359 11036 45554 11064
rect 40359 11033 40371 11036
rect 40313 11027 40371 11033
rect 31628 10968 33732 10996
rect 45526 10996 45554 11036
rect 45833 11033 45845 11067
rect 45879 11064 45891 11067
rect 47210 11064 47216 11076
rect 45879 11036 47216 11064
rect 45879 11033 45891 11036
rect 45833 11027 45891 11033
rect 47210 11024 47216 11036
rect 47268 11024 47274 11076
rect 46106 10996 46112 11008
rect 45526 10968 46112 10996
rect 31628 10956 31634 10968
rect 46106 10956 46112 10968
rect 46164 10956 46170 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10792 2283 10795
rect 2774 10792 2780 10804
rect 2271 10764 2780 10792
rect 2271 10761 2283 10764
rect 2225 10755 2283 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4019 10764 6914 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 6886 10724 6914 10764
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 12253 10795 12311 10801
rect 12253 10792 12265 10795
rect 11848 10764 12265 10792
rect 11848 10752 11854 10764
rect 12253 10761 12265 10764
rect 12299 10761 12311 10795
rect 12253 10755 12311 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12860 10764 13185 10792
rect 12860 10752 12866 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 14366 10752 14372 10804
rect 14424 10752 14430 10804
rect 14737 10795 14795 10801
rect 14737 10761 14749 10795
rect 14783 10792 14795 10795
rect 15838 10792 15844 10804
rect 14783 10764 15844 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 13998 10724 14004 10736
rect 6886 10696 14004 10724
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1360 10628 1593 10656
rect 1360 10616 1366 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2731 10628 2765 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 1210 10548 1216 10600
rect 1268 10588 1274 10600
rect 2700 10588 2728 10619
rect 3786 10616 3792 10668
rect 3844 10616 3850 10668
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 12124 10628 13553 10656
rect 12124 10616 12130 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 13630 10616 13636 10668
rect 13688 10616 13694 10668
rect 14752 10656 14780 10755
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 15979 10764 17141 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17494 10752 17500 10804
rect 17552 10752 17558 10804
rect 18138 10752 18144 10804
rect 18196 10792 18202 10804
rect 18325 10795 18383 10801
rect 18325 10792 18337 10795
rect 18196 10764 18337 10792
rect 18196 10752 18202 10764
rect 18325 10761 18337 10764
rect 18371 10761 18383 10795
rect 19521 10795 19579 10801
rect 18325 10755 18383 10761
rect 18616 10764 19012 10792
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 16758 10724 16764 10736
rect 14875 10696 16764 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 16758 10684 16764 10696
rect 16816 10684 16822 10736
rect 17586 10684 17592 10736
rect 17644 10684 17650 10736
rect 13740 10628 14780 10656
rect 3418 10588 3424 10600
rect 1268 10560 3424 10588
rect 1268 10548 1274 10560
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10588 12587 10591
rect 13648 10588 13676 10616
rect 12575 10560 13676 10588
rect 12575 10557 12587 10560
rect 12529 10551 12587 10557
rect 12713 10523 12771 10529
rect 12713 10489 12725 10523
rect 12759 10520 12771 10523
rect 13740 10520 13768 10628
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 15068 10628 16252 10656
rect 15068 10616 15074 10628
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 14642 10588 14648 10600
rect 13863 10560 14648 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16224 10588 16252 10628
rect 16482 10616 16488 10668
rect 16540 10656 16546 10668
rect 18616 10656 18644 10764
rect 18984 10724 19012 10764
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19702 10792 19708 10804
rect 19567 10764 19708 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 20717 10795 20775 10801
rect 20717 10761 20729 10795
rect 20763 10761 20775 10795
rect 20717 10755 20775 10761
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 22646 10792 22652 10804
rect 21131 10764 22652 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 20732 10724 20760 10755
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 24210 10752 24216 10804
rect 24268 10752 24274 10804
rect 26326 10752 26332 10804
rect 26384 10792 26390 10804
rect 27062 10792 27068 10804
rect 26384 10764 27068 10792
rect 26384 10752 26390 10764
rect 27062 10752 27068 10764
rect 27120 10792 27126 10804
rect 27525 10795 27583 10801
rect 27525 10792 27537 10795
rect 27120 10764 27537 10792
rect 27120 10752 27126 10764
rect 27525 10761 27537 10764
rect 27571 10761 27583 10795
rect 27525 10755 27583 10761
rect 28537 10795 28595 10801
rect 28537 10761 28549 10795
rect 28583 10792 28595 10795
rect 28718 10792 28724 10804
rect 28583 10764 28724 10792
rect 28583 10761 28595 10764
rect 28537 10755 28595 10761
rect 28718 10752 28724 10764
rect 28776 10792 28782 10804
rect 28776 10764 28856 10792
rect 28776 10752 28782 10764
rect 18984 10696 20760 10724
rect 21177 10727 21235 10733
rect 21177 10693 21189 10727
rect 21223 10724 21235 10727
rect 22278 10724 22284 10736
rect 21223 10696 22284 10724
rect 21223 10693 21235 10696
rect 21177 10687 21235 10693
rect 22278 10684 22284 10696
rect 22336 10684 22342 10736
rect 23842 10724 23848 10736
rect 23506 10696 23848 10724
rect 23842 10684 23848 10696
rect 23900 10684 23906 10736
rect 24504 10696 27292 10724
rect 16540 10628 18644 10656
rect 16540 10616 16546 10628
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 19794 10616 19800 10668
rect 19852 10656 19858 10668
rect 19889 10659 19947 10665
rect 19889 10656 19901 10659
rect 19852 10628 19901 10656
rect 19852 10616 19858 10628
rect 19889 10625 19901 10628
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 20254 10616 20260 10668
rect 20312 10656 20318 10668
rect 20312 10628 21496 10656
rect 20312 10616 20318 10628
rect 17681 10591 17739 10597
rect 17681 10588 17693 10591
rect 16224 10560 17693 10588
rect 16117 10551 16175 10557
rect 17681 10557 17693 10560
rect 17727 10557 17739 10591
rect 17681 10551 17739 10557
rect 12759 10492 13768 10520
rect 12759 10489 12771 10492
rect 12713 10483 12771 10489
rect 3326 10412 3332 10464
rect 3384 10412 3390 10464
rect 12066 10412 12072 10464
rect 12124 10412 12130 10464
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 12728 10452 12756 10483
rect 15654 10480 15660 10532
rect 15712 10480 15718 10532
rect 15930 10480 15936 10532
rect 15988 10520 15994 10532
rect 16132 10520 16160 10551
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18012 10560 18797 10588
rect 18012 10548 18018 10560
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 18785 10551 18843 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19150 10588 19156 10600
rect 19015 10560 19156 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 21082 10588 21088 10600
rect 20211 10560 21088 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 15988 10492 16160 10520
rect 16853 10523 16911 10529
rect 15988 10480 15994 10492
rect 16853 10489 16865 10523
rect 16899 10520 16911 10523
rect 19996 10520 20024 10551
rect 21082 10548 21088 10560
rect 21140 10548 21146 10600
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 20622 10520 20628 10532
rect 16899 10492 20628 10520
rect 16899 10489 16911 10492
rect 16853 10483 16911 10489
rect 20622 10480 20628 10492
rect 20680 10480 20686 10532
rect 12584 10424 12756 10452
rect 12584 10412 12590 10424
rect 12802 10412 12808 10464
rect 12860 10452 12866 10464
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12860 10424 12909 10452
rect 12860 10412 12866 10424
rect 12897 10421 12909 10424
rect 12943 10452 12955 10455
rect 14734 10452 14740 10464
rect 12943 10424 14740 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 15565 10455 15623 10461
rect 15565 10421 15577 10455
rect 15611 10452 15623 10455
rect 15672 10452 15700 10480
rect 15611 10424 15700 10452
rect 15611 10421 15623 10424
rect 15565 10415 15623 10421
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 17494 10452 17500 10464
rect 16724 10424 17500 10452
rect 16724 10412 16730 10424
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 17586 10412 17592 10464
rect 17644 10452 17650 10464
rect 21266 10452 21272 10464
rect 17644 10424 21272 10452
rect 17644 10412 17650 10424
rect 21266 10412 21272 10424
rect 21324 10412 21330 10464
rect 21376 10452 21404 10551
rect 21468 10520 21496 10628
rect 22002 10548 22008 10600
rect 22060 10548 22066 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22112 10560 22293 10588
rect 22112 10520 22140 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 23934 10548 23940 10600
rect 23992 10588 23998 10600
rect 24504 10588 24532 10696
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25409 10659 25467 10665
rect 25409 10656 25421 10659
rect 24627 10628 25421 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 25409 10625 25421 10628
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 25961 10659 26019 10665
rect 25961 10625 25973 10659
rect 26007 10656 26019 10659
rect 26694 10656 26700 10668
rect 26007 10628 26700 10656
rect 26007 10625 26019 10628
rect 25961 10619 26019 10625
rect 26694 10616 26700 10628
rect 26752 10616 26758 10668
rect 27264 10656 27292 10696
rect 27338 10684 27344 10736
rect 27396 10724 27402 10736
rect 28828 10733 28856 10764
rect 29914 10752 29920 10804
rect 29972 10792 29978 10804
rect 30561 10795 30619 10801
rect 30561 10792 30573 10795
rect 29972 10764 30573 10792
rect 29972 10752 29978 10764
rect 30561 10761 30573 10764
rect 30607 10761 30619 10795
rect 30561 10755 30619 10761
rect 31110 10752 31116 10804
rect 31168 10792 31174 10804
rect 31389 10795 31447 10801
rect 31389 10792 31401 10795
rect 31168 10764 31401 10792
rect 31168 10752 31174 10764
rect 31389 10761 31401 10764
rect 31435 10761 31447 10795
rect 31389 10755 31447 10761
rect 33045 10795 33103 10801
rect 33045 10761 33057 10795
rect 33091 10792 33103 10795
rect 33091 10764 36768 10792
rect 33091 10761 33103 10764
rect 33045 10755 33103 10761
rect 28815 10727 28873 10733
rect 27396 10696 28764 10724
rect 27396 10684 27402 10696
rect 28736 10656 28764 10696
rect 28815 10693 28827 10727
rect 28861 10693 28873 10727
rect 28815 10687 28873 10693
rect 29546 10684 29552 10736
rect 29604 10724 29610 10736
rect 30282 10724 30288 10736
rect 29604 10696 30288 10724
rect 29604 10684 29610 10696
rect 30282 10684 30288 10696
rect 30340 10684 30346 10736
rect 31478 10684 31484 10736
rect 31536 10724 31542 10736
rect 33318 10724 33324 10736
rect 31536 10696 33324 10724
rect 31536 10684 31542 10696
rect 33318 10684 33324 10696
rect 33376 10724 33382 10736
rect 35345 10727 35403 10733
rect 33376 10696 34178 10724
rect 33376 10684 33382 10696
rect 35345 10693 35357 10727
rect 35391 10724 35403 10727
rect 36630 10724 36636 10736
rect 35391 10696 36636 10724
rect 35391 10693 35403 10696
rect 35345 10687 35403 10693
rect 36630 10684 36636 10696
rect 36688 10684 36694 10736
rect 36740 10724 36768 10764
rect 36814 10752 36820 10804
rect 36872 10752 36878 10804
rect 37274 10724 37280 10736
rect 36740 10696 37280 10724
rect 37274 10684 37280 10696
rect 37332 10684 37338 10736
rect 49145 10727 49203 10733
rect 49145 10693 49157 10727
rect 49191 10724 49203 10727
rect 49234 10724 49240 10736
rect 49191 10696 49240 10724
rect 49191 10693 49203 10696
rect 49145 10687 49203 10693
rect 49234 10684 49240 10696
rect 49292 10684 49298 10736
rect 29730 10656 29736 10668
rect 27264 10628 28672 10656
rect 28736 10628 29736 10656
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 23992 10560 24685 10588
rect 23992 10548 23998 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 24857 10591 24915 10597
rect 24857 10557 24869 10591
rect 24903 10588 24915 10591
rect 26602 10588 26608 10600
rect 24903 10560 26608 10588
rect 24903 10557 24915 10560
rect 24857 10551 24915 10557
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 27338 10548 27344 10600
rect 27396 10548 27402 10600
rect 27433 10591 27491 10597
rect 27433 10557 27445 10591
rect 27479 10557 27491 10591
rect 28644 10588 28672 10628
rect 29730 10616 29736 10628
rect 29788 10656 29794 10668
rect 29788 10628 30604 10656
rect 29788 10616 29794 10628
rect 29454 10588 29460 10600
rect 28644 10560 29460 10588
rect 27433 10551 27491 10557
rect 21468 10492 22140 10520
rect 23566 10480 23572 10532
rect 23624 10520 23630 10532
rect 23753 10523 23811 10529
rect 23753 10520 23765 10523
rect 23624 10492 23765 10520
rect 23624 10480 23630 10492
rect 23753 10489 23765 10492
rect 23799 10520 23811 10523
rect 24762 10520 24768 10532
rect 23799 10492 24768 10520
rect 23799 10489 23811 10492
rect 23753 10483 23811 10489
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 27448 10520 27476 10551
rect 29454 10548 29460 10560
rect 29512 10548 29518 10600
rect 29546 10548 29552 10600
rect 29604 10548 29610 10600
rect 29822 10548 29828 10600
rect 29880 10588 29886 10600
rect 30377 10591 30435 10597
rect 30377 10588 30389 10591
rect 29880 10560 30389 10588
rect 29880 10548 29886 10560
rect 30377 10557 30389 10560
rect 30423 10557 30435 10591
rect 30377 10551 30435 10557
rect 30466 10548 30472 10600
rect 30524 10548 30530 10600
rect 30576 10588 30604 10628
rect 30650 10616 30656 10668
rect 30708 10656 30714 10668
rect 32677 10659 32735 10665
rect 32677 10656 32689 10659
rect 30708 10628 32689 10656
rect 30708 10616 30714 10628
rect 32677 10625 32689 10628
rect 32723 10625 32735 10659
rect 32677 10619 32735 10625
rect 35618 10616 35624 10668
rect 35676 10616 35682 10668
rect 36446 10616 36452 10668
rect 36504 10616 36510 10668
rect 39761 10659 39819 10665
rect 39761 10625 39773 10659
rect 39807 10656 39819 10659
rect 40221 10659 40279 10665
rect 40221 10656 40233 10659
rect 39807 10628 40233 10656
rect 39807 10625 39819 10628
rect 39761 10619 39819 10625
rect 40221 10625 40233 10628
rect 40267 10625 40279 10659
rect 40221 10619 40279 10625
rect 32214 10588 32220 10600
rect 30576 10560 32220 10588
rect 32214 10548 32220 10560
rect 32272 10548 32278 10600
rect 32306 10548 32312 10600
rect 32364 10588 32370 10600
rect 32401 10591 32459 10597
rect 32401 10588 32413 10591
rect 32364 10560 32413 10588
rect 32364 10548 32370 10560
rect 32401 10557 32413 10560
rect 32447 10557 32459 10591
rect 32401 10551 32459 10557
rect 32585 10591 32643 10597
rect 32585 10557 32597 10591
rect 32631 10557 32643 10591
rect 32585 10551 32643 10557
rect 26068 10492 27476 10520
rect 27893 10523 27951 10529
rect 26068 10464 26096 10492
rect 27893 10489 27905 10523
rect 27939 10520 27951 10523
rect 32600 10520 32628 10551
rect 34698 10548 34704 10600
rect 34756 10588 34762 10600
rect 36173 10591 36231 10597
rect 36173 10588 36185 10591
rect 34756 10560 36185 10588
rect 34756 10548 34762 10560
rect 36173 10557 36185 10560
rect 36219 10557 36231 10591
rect 36173 10551 36231 10557
rect 36354 10548 36360 10600
rect 36412 10548 36418 10600
rect 39776 10588 39804 10619
rect 47210 10616 47216 10668
rect 47268 10656 47274 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 47268 10628 47961 10656
rect 47268 10616 47274 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 36464 10560 39804 10588
rect 33873 10523 33931 10529
rect 33873 10520 33885 10523
rect 27939 10492 32628 10520
rect 32692 10492 33885 10520
rect 27939 10489 27951 10492
rect 27893 10483 27951 10489
rect 22094 10452 22100 10464
rect 21376 10424 22100 10452
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 26050 10412 26056 10464
rect 26108 10412 26114 10464
rect 26513 10455 26571 10461
rect 26513 10421 26525 10455
rect 26559 10452 26571 10455
rect 26694 10452 26700 10464
rect 26559 10424 26700 10452
rect 26559 10421 26571 10424
rect 26513 10415 26571 10421
rect 26694 10412 26700 10424
rect 26752 10412 26758 10464
rect 26789 10455 26847 10461
rect 26789 10421 26801 10455
rect 26835 10452 26847 10455
rect 27430 10452 27436 10464
rect 26835 10424 27436 10452
rect 26835 10421 26847 10424
rect 26789 10415 26847 10421
rect 27430 10412 27436 10424
rect 27488 10452 27494 10464
rect 30742 10452 30748 10464
rect 27488 10424 30748 10452
rect 27488 10412 27494 10424
rect 30742 10412 30748 10424
rect 30800 10412 30806 10464
rect 30929 10455 30987 10461
rect 30929 10421 30941 10455
rect 30975 10452 30987 10455
rect 31754 10452 31760 10464
rect 30975 10424 31760 10452
rect 30975 10421 30987 10424
rect 30929 10415 30987 10421
rect 31754 10412 31760 10424
rect 31812 10412 31818 10464
rect 31846 10412 31852 10464
rect 31904 10412 31910 10464
rect 32214 10412 32220 10464
rect 32272 10452 32278 10464
rect 32692 10452 32720 10492
rect 33873 10489 33885 10492
rect 33919 10489 33931 10523
rect 33873 10483 33931 10489
rect 35618 10480 35624 10532
rect 35676 10520 35682 10532
rect 36464 10520 36492 10560
rect 35676 10492 36492 10520
rect 35676 10480 35682 10492
rect 36538 10480 36544 10532
rect 36596 10520 36602 10532
rect 38930 10520 38936 10532
rect 36596 10492 38936 10520
rect 36596 10480 36602 10492
rect 38930 10480 38936 10492
rect 38988 10480 38994 10532
rect 39945 10523 40003 10529
rect 39945 10489 39957 10523
rect 39991 10520 40003 10523
rect 46934 10520 46940 10532
rect 39991 10492 46940 10520
rect 39991 10489 40003 10492
rect 39945 10483 40003 10489
rect 46934 10480 46940 10492
rect 46992 10480 46998 10532
rect 32272 10424 32720 10452
rect 32272 10412 32278 10424
rect 36906 10412 36912 10464
rect 36964 10452 36970 10464
rect 37277 10455 37335 10461
rect 37277 10452 37289 10455
rect 36964 10424 37289 10452
rect 36964 10412 36970 10424
rect 37277 10421 37289 10424
rect 37323 10452 37335 10455
rect 37461 10455 37519 10461
rect 37461 10452 37473 10455
rect 37323 10424 37473 10452
rect 37323 10421 37335 10424
rect 37277 10415 37335 10421
rect 37461 10421 37473 10424
rect 37507 10452 37519 10455
rect 38562 10452 38568 10464
rect 37507 10424 38568 10452
rect 37507 10421 37519 10424
rect 37461 10415 37519 10421
rect 38562 10412 38568 10424
rect 38620 10412 38626 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 1302 10208 1308 10260
rect 1360 10208 1366 10260
rect 2179 10251 2237 10257
rect 2179 10217 2191 10251
rect 2225 10248 2237 10251
rect 5442 10248 5448 10260
rect 2225 10220 5448 10248
rect 2225 10217 2237 10220
rect 2179 10211 2237 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 13449 10251 13507 10257
rect 13449 10217 13461 10251
rect 13495 10248 13507 10251
rect 16022 10248 16028 10260
rect 13495 10220 16028 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16666 10208 16672 10260
rect 16724 10208 16730 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 17276 10220 18153 10248
rect 17276 10208 17282 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 18322 10208 18328 10260
rect 18380 10248 18386 10260
rect 19150 10248 19156 10260
rect 18380 10220 19156 10248
rect 18380 10208 18386 10220
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 20254 10208 20260 10260
rect 20312 10208 20318 10260
rect 20364 10220 22094 10248
rect 1320 10180 1348 10208
rect 3789 10183 3847 10189
rect 3789 10180 3801 10183
rect 1320 10152 3801 10180
rect 3789 10149 3801 10152
rect 3835 10149 3847 10183
rect 14734 10180 14740 10192
rect 3789 10143 3847 10149
rect 12912 10152 14740 10180
rect 1302 10072 1308 10124
rect 1360 10112 1366 10124
rect 12912 10121 12940 10152
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 17310 10180 17316 10192
rect 15948 10152 17316 10180
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 1360 10084 2421 10112
rect 1360 10072 1366 10084
rect 2409 10081 2421 10084
rect 2455 10112 2467 10115
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 2455 10084 3985 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 15948 10112 15976 10152
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 17494 10140 17500 10192
rect 17552 10180 17558 10192
rect 19794 10180 19800 10192
rect 17552 10152 19800 10180
rect 17552 10140 17558 10152
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 13035 10084 15976 10112
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 16574 10072 16580 10124
rect 16632 10112 16638 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 16632 10084 17417 10112
rect 16632 10072 16638 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10112 17647 10115
rect 17862 10112 17868 10124
rect 17635 10084 17868 10112
rect 17635 10081 17647 10084
rect 17589 10075 17647 10081
rect 17862 10072 17868 10084
rect 17920 10112 17926 10124
rect 18322 10112 18328 10124
rect 17920 10084 18328 10112
rect 17920 10072 17926 10084
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 18598 10072 18604 10124
rect 18656 10072 18662 10124
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 19426 10112 19432 10124
rect 18831 10084 19432 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19668 10084 19717 10112
rect 19668 10072 19674 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3326 10044 3332 10056
rect 3191 10016 3332 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 13078 10044 13084 10056
rect 12492 10016 13084 10044
rect 12492 10004 12498 10016
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13596 10016 13829 10044
rect 13596 10004 13602 10016
rect 13817 10013 13829 10016
rect 13863 10044 13875 10047
rect 13863 10016 14674 10044
rect 13863 10013 13875 10016
rect 13817 10007 13875 10013
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10044 16543 10047
rect 18506 10044 18512 10056
rect 16531 10016 18512 10044
rect 16531 10013 16543 10016
rect 16485 10007 16543 10013
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 20364 10044 20392 10220
rect 22066 10180 22094 10220
rect 23750 10208 23756 10260
rect 23808 10208 23814 10260
rect 24302 10208 24308 10260
rect 24360 10248 24366 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 24360 10220 24593 10248
rect 24360 10208 24366 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 26326 10248 26332 10260
rect 24581 10211 24639 10217
rect 24688 10220 26332 10248
rect 24688 10180 24716 10220
rect 26326 10208 26332 10220
rect 26384 10208 26390 10260
rect 28721 10251 28779 10257
rect 28721 10217 28733 10251
rect 28767 10248 28779 10251
rect 29086 10248 29092 10260
rect 28767 10220 29092 10248
rect 28767 10217 28779 10220
rect 28721 10211 28779 10217
rect 29086 10208 29092 10220
rect 29144 10248 29150 10260
rect 29822 10248 29828 10260
rect 29144 10220 29828 10248
rect 29144 10208 29150 10220
rect 29822 10208 29828 10220
rect 29880 10208 29886 10260
rect 30374 10208 30380 10260
rect 30432 10208 30438 10260
rect 32030 10208 32036 10260
rect 32088 10248 32094 10260
rect 32088 10220 36400 10248
rect 32088 10208 32094 10220
rect 26602 10180 26608 10192
rect 22066 10152 24716 10180
rect 26252 10152 26608 10180
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21729 10115 21787 10121
rect 21729 10112 21741 10115
rect 21140 10084 21741 10112
rect 21140 10072 21146 10084
rect 21729 10081 21741 10084
rect 21775 10081 21787 10115
rect 21729 10075 21787 10081
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10112 26111 10115
rect 26252 10112 26280 10152
rect 26602 10140 26608 10152
rect 26660 10140 26666 10192
rect 28994 10140 29000 10192
rect 29052 10140 29058 10192
rect 29362 10140 29368 10192
rect 29420 10140 29426 10192
rect 30006 10140 30012 10192
rect 30064 10180 30070 10192
rect 34422 10180 34428 10192
rect 30064 10152 30788 10180
rect 30064 10140 30070 10152
rect 26099 10084 26280 10112
rect 26329 10115 26387 10121
rect 26099 10081 26111 10084
rect 26053 10075 26111 10081
rect 26329 10081 26341 10115
rect 26375 10112 26387 10115
rect 26878 10112 26884 10124
rect 26375 10084 26884 10112
rect 26375 10081 26387 10084
rect 26329 10075 26387 10081
rect 26878 10072 26884 10084
rect 26936 10112 26942 10124
rect 26973 10115 27031 10121
rect 26973 10112 26985 10115
rect 26936 10084 26985 10112
rect 26936 10072 26942 10084
rect 26973 10081 26985 10084
rect 27019 10112 27031 10115
rect 29546 10112 29552 10124
rect 27019 10084 29552 10112
rect 27019 10081 27031 10084
rect 26973 10075 27031 10081
rect 29546 10072 29552 10084
rect 29604 10072 29610 10124
rect 29917 10115 29975 10121
rect 29917 10081 29929 10115
rect 29963 10112 29975 10115
rect 30650 10112 30656 10124
rect 29963 10084 30656 10112
rect 29963 10081 29975 10084
rect 29917 10075 29975 10081
rect 30650 10072 30656 10084
rect 30708 10072 30714 10124
rect 30760 10112 30788 10152
rect 32048 10152 34428 10180
rect 32048 10112 32076 10152
rect 34422 10140 34428 10152
rect 34480 10140 34486 10192
rect 30760 10084 32076 10112
rect 32122 10072 32128 10124
rect 32180 10072 32186 10124
rect 32214 10072 32220 10124
rect 32272 10112 32278 10124
rect 32677 10115 32735 10121
rect 32677 10112 32689 10115
rect 32272 10084 32689 10112
rect 32272 10072 32278 10084
rect 32677 10081 32689 10084
rect 32723 10081 32735 10115
rect 32677 10075 32735 10081
rect 32766 10072 32772 10124
rect 32824 10112 32830 10124
rect 32861 10115 32919 10121
rect 32861 10112 32873 10115
rect 32824 10084 32873 10112
rect 32824 10072 32830 10084
rect 32861 10081 32873 10084
rect 32907 10081 32919 10115
rect 32861 10075 32919 10081
rect 34698 10072 34704 10124
rect 34756 10112 34762 10124
rect 35158 10112 35164 10124
rect 34756 10084 35164 10112
rect 34756 10072 34762 10084
rect 35158 10072 35164 10084
rect 35216 10072 35222 10124
rect 18616 10016 20392 10044
rect 14458 9976 14464 9988
rect 2976 9948 14464 9976
rect 2976 9917 3004 9948
rect 14458 9936 14464 9948
rect 14516 9936 14522 9988
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9945 15807 9979
rect 15749 9939 15807 9945
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9877 3019 9911
rect 2961 9871 3019 9877
rect 14274 9868 14280 9920
rect 14332 9868 14338 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 15010 9908 15016 9920
rect 14792 9880 15016 9908
rect 14792 9868 14798 9880
rect 15010 9868 15016 9880
rect 15068 9908 15074 9920
rect 15764 9908 15792 9939
rect 15838 9936 15844 9988
rect 15896 9976 15902 9988
rect 18616 9976 18644 10016
rect 22002 10004 22008 10056
rect 22060 10044 22066 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 22060 10016 23213 10044
rect 22060 10004 22066 10016
rect 23201 10013 23213 10016
rect 23247 10044 23259 10047
rect 24026 10044 24032 10056
rect 23247 10016 24032 10044
rect 23247 10013 23259 10016
rect 23201 10007 23259 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 30742 10004 30748 10056
rect 30800 10004 30806 10056
rect 32140 10044 32168 10072
rect 32490 10044 32496 10056
rect 32140 10016 32496 10044
rect 32490 10004 32496 10016
rect 32548 10004 32554 10056
rect 33502 10004 33508 10056
rect 33560 10044 33566 10056
rect 33560 10016 34284 10044
rect 33560 10004 33566 10016
rect 15896 9948 18644 9976
rect 15896 9936 15902 9948
rect 15068 9880 15792 9908
rect 15068 9868 15074 9880
rect 16942 9868 16948 9920
rect 17000 9868 17006 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 17313 9911 17371 9917
rect 17313 9908 17325 9911
rect 17276 9880 17325 9908
rect 17276 9868 17282 9880
rect 17313 9877 17325 9880
rect 17359 9877 17371 9911
rect 17313 9871 17371 9877
rect 18509 9911 18567 9917
rect 18509 9877 18521 9911
rect 18555 9908 18567 9911
rect 18616 9908 18644 9948
rect 19794 9936 19800 9988
rect 19852 9976 19858 9988
rect 20438 9976 20444 9988
rect 19852 9948 20444 9976
rect 19852 9936 19858 9948
rect 20438 9936 20444 9948
rect 20496 9976 20502 9988
rect 20496 9948 20562 9976
rect 20496 9936 20502 9948
rect 18555 9880 18644 9908
rect 18555 9877 18567 9880
rect 18509 9871 18567 9877
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 22020 9908 22048 10004
rect 34256 9988 34284 10016
rect 34882 10004 34888 10056
rect 34940 10004 34946 10056
rect 36372 10044 36400 10220
rect 36630 10208 36636 10260
rect 36688 10208 36694 10260
rect 38473 10115 38531 10121
rect 38473 10081 38485 10115
rect 38519 10112 38531 10115
rect 47118 10112 47124 10124
rect 38519 10084 47124 10112
rect 38519 10081 38531 10084
rect 38473 10075 38531 10081
rect 47118 10072 47124 10084
rect 47176 10072 47182 10124
rect 49142 10072 49148 10124
rect 49200 10072 49206 10124
rect 38289 10047 38347 10053
rect 38289 10044 38301 10047
rect 36372 10016 38301 10044
rect 38289 10013 38301 10016
rect 38335 10044 38347 10047
rect 38749 10047 38807 10053
rect 38749 10044 38761 10047
rect 38335 10016 38761 10044
rect 38335 10013 38347 10016
rect 38289 10007 38347 10013
rect 38749 10013 38761 10016
rect 38795 10013 38807 10047
rect 38749 10007 38807 10013
rect 38930 10004 38936 10056
rect 38988 10044 38994 10056
rect 40129 10047 40187 10053
rect 40129 10044 40141 10047
rect 38988 10016 40141 10044
rect 38988 10004 38994 10016
rect 40129 10013 40141 10016
rect 40175 10013 40187 10047
rect 40129 10007 40187 10013
rect 40313 10047 40371 10053
rect 40313 10013 40325 10047
rect 40359 10044 40371 10047
rect 45830 10044 45836 10056
rect 40359 10016 45836 10044
rect 40359 10013 40371 10016
rect 40313 10007 40371 10013
rect 22462 9936 22468 9988
rect 22520 9936 22526 9988
rect 23842 9936 23848 9988
rect 23900 9976 23906 9988
rect 23900 9948 24808 9976
rect 25622 9948 26004 9976
rect 23900 9936 23906 9948
rect 21508 9880 22048 9908
rect 21508 9868 21514 9880
rect 23934 9868 23940 9920
rect 23992 9908 23998 9920
rect 24029 9911 24087 9917
rect 24029 9908 24041 9911
rect 23992 9880 24041 9908
rect 23992 9868 23998 9880
rect 24029 9877 24041 9880
rect 24075 9877 24087 9911
rect 24780 9908 24808 9948
rect 25038 9908 25044 9920
rect 24780 9880 25044 9908
rect 24029 9871 24087 9877
rect 25038 9868 25044 9880
rect 25096 9908 25102 9920
rect 25700 9908 25728 9948
rect 25096 9880 25728 9908
rect 25976 9908 26004 9948
rect 26050 9936 26056 9988
rect 26108 9976 26114 9988
rect 26108 9948 26832 9976
rect 26108 9936 26114 9948
rect 26694 9908 26700 9920
rect 25976 9880 26700 9908
rect 25096 9868 25102 9880
rect 26694 9868 26700 9880
rect 26752 9868 26758 9920
rect 26804 9908 26832 9948
rect 27246 9936 27252 9988
rect 27304 9936 27310 9988
rect 28534 9976 28540 9988
rect 28474 9948 28540 9976
rect 28534 9936 28540 9948
rect 28592 9976 28598 9988
rect 28718 9976 28724 9988
rect 28592 9948 28724 9976
rect 28592 9936 28598 9948
rect 28718 9936 28724 9948
rect 28776 9936 28782 9988
rect 31849 9979 31907 9985
rect 28920 9948 29408 9976
rect 28920 9908 28948 9948
rect 26804 9880 28948 9908
rect 29380 9908 29408 9948
rect 31849 9945 31861 9979
rect 31895 9976 31907 9979
rect 31938 9976 31944 9988
rect 31895 9948 31944 9976
rect 31895 9945 31907 9948
rect 31849 9939 31907 9945
rect 31938 9936 31944 9948
rect 31996 9936 32002 9988
rect 32674 9936 32680 9988
rect 32732 9976 32738 9988
rect 33781 9979 33839 9985
rect 33781 9976 33793 9979
rect 32732 9948 33793 9976
rect 32732 9936 32738 9948
rect 33781 9945 33793 9948
rect 33827 9945 33839 9979
rect 33781 9939 33839 9945
rect 34238 9936 34244 9988
rect 34296 9976 34302 9988
rect 35434 9976 35440 9988
rect 34296 9948 35440 9976
rect 34296 9936 34302 9948
rect 35434 9936 35440 9948
rect 35492 9936 35498 9988
rect 35710 9936 35716 9988
rect 35768 9936 35774 9988
rect 40144 9976 40172 10007
rect 45830 10004 45836 10016
rect 45888 10004 45894 10056
rect 46106 10004 46112 10056
rect 46164 10004 46170 10056
rect 46658 10004 46664 10056
rect 46716 10044 46722 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46716 10016 47961 10044
rect 46716 10004 46722 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 40589 9979 40647 9985
rect 40589 9976 40601 9979
rect 40144 9948 40601 9976
rect 40589 9945 40601 9948
rect 40635 9945 40647 9979
rect 40589 9939 40647 9945
rect 44358 9936 44364 9988
rect 44416 9936 44422 9988
rect 44545 9979 44603 9985
rect 44545 9945 44557 9979
rect 44591 9976 44603 9979
rect 46750 9976 46756 9988
rect 44591 9948 46756 9976
rect 44591 9945 44603 9948
rect 44545 9939 44603 9945
rect 46750 9936 46756 9948
rect 46808 9936 46814 9988
rect 47302 9936 47308 9988
rect 47360 9936 47366 9988
rect 32030 9908 32036 9920
rect 29380 9880 32036 9908
rect 32030 9868 32036 9880
rect 32088 9868 32094 9920
rect 32398 9868 32404 9920
rect 32456 9908 32462 9920
rect 32953 9911 33011 9917
rect 32953 9908 32965 9911
rect 32456 9880 32965 9908
rect 32456 9868 32462 9880
rect 32953 9877 32965 9880
rect 32999 9877 33011 9911
rect 32953 9871 33011 9877
rect 33321 9911 33379 9917
rect 33321 9877 33333 9911
rect 33367 9908 33379 9911
rect 36814 9908 36820 9920
rect 33367 9880 36820 9908
rect 33367 9877 33379 9880
rect 33321 9871 33379 9877
rect 36814 9868 36820 9880
rect 36872 9868 36878 9920
rect 36906 9868 36912 9920
rect 36964 9868 36970 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 16666 9664 16672 9716
rect 16724 9704 16730 9716
rect 16724 9676 21036 9704
rect 16724 9664 16730 9676
rect 2225 9639 2283 9645
rect 2225 9605 2237 9639
rect 2271 9636 2283 9639
rect 3786 9636 3792 9648
rect 2271 9608 3792 9636
rect 2271 9605 2283 9608
rect 2225 9599 2283 9605
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12618 9636 12624 9648
rect 12483 9608 12624 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 13357 9639 13415 9645
rect 13357 9605 13369 9639
rect 13403 9636 13415 9639
rect 13722 9636 13728 9648
rect 13403 9608 13728 9636
rect 13403 9605 13415 9608
rect 13357 9599 13415 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 14642 9596 14648 9648
rect 14700 9596 14706 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 16022 9636 16028 9648
rect 15252 9608 16028 9636
rect 15252 9596 15258 9608
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2740 9540 2973 9568
rect 2740 9528 2746 9540
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 1596 9432 1624 9528
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 3528 9500 3556 9531
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 15396 9577 15424 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 16114 9596 16120 9648
rect 16172 9636 16178 9648
rect 16209 9639 16267 9645
rect 16209 9636 16221 9639
rect 16172 9608 16221 9636
rect 16172 9596 16178 9608
rect 16209 9605 16221 9608
rect 16255 9636 16267 9639
rect 16853 9639 16911 9645
rect 16853 9636 16865 9639
rect 16255 9608 16865 9636
rect 16255 9605 16267 9608
rect 16209 9599 16267 9605
rect 16853 9605 16865 9608
rect 16899 9605 16911 9639
rect 16853 9599 16911 9605
rect 19702 9596 19708 9648
rect 19760 9636 19766 9648
rect 21008 9636 21036 9676
rect 21082 9664 21088 9716
rect 21140 9664 21146 9716
rect 26050 9704 26056 9716
rect 21192 9676 26056 9704
rect 21192 9636 21220 9676
rect 26050 9664 26056 9676
rect 26108 9664 26114 9716
rect 26694 9664 26700 9716
rect 26752 9704 26758 9716
rect 28718 9704 28724 9716
rect 26752 9676 28724 9704
rect 26752 9664 26758 9676
rect 19760 9608 20102 9636
rect 21008 9608 21220 9636
rect 19760 9596 19766 9608
rect 21542 9596 21548 9648
rect 21600 9636 21606 9648
rect 22554 9636 22560 9648
rect 21600 9608 22560 9636
rect 21600 9596 21606 9608
rect 22554 9596 22560 9608
rect 22612 9636 22618 9648
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 22612 9608 22753 9636
rect 22612 9596 22618 9608
rect 22741 9605 22753 9608
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 24670 9596 24676 9648
rect 24728 9636 24734 9648
rect 27246 9636 27252 9648
rect 24728 9608 25268 9636
rect 24728 9596 24734 9608
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12400 9540 12541 9568
rect 12400 9528 12406 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9568 15807 9571
rect 15838 9568 15844 9580
rect 15795 9540 15844 9568
rect 15795 9537 15807 9540
rect 15749 9531 15807 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 16482 9528 16488 9580
rect 16540 9528 16546 9580
rect 17494 9528 17500 9580
rect 17552 9528 17558 9580
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9568 22707 9571
rect 23382 9568 23388 9580
rect 22695 9540 23388 9568
rect 22695 9537 22707 9540
rect 22649 9531 22707 9537
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23842 9528 23848 9580
rect 23900 9528 23906 9580
rect 25240 9577 25268 9608
rect 25884 9608 27252 9636
rect 25225 9571 25283 9577
rect 25225 9537 25237 9571
rect 25271 9537 25283 9571
rect 25225 9531 25283 9537
rect 2280 9472 3556 9500
rect 2280 9460 2286 9472
rect 3694 9460 3700 9512
rect 3752 9460 3758 9512
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11112 9472 12265 9500
rect 11112 9460 11118 9472
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 15102 9460 15108 9512
rect 15160 9460 15166 9512
rect 15933 9503 15991 9509
rect 15933 9469 15945 9503
rect 15979 9500 15991 9503
rect 17586 9500 17592 9512
rect 15979 9472 17592 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18598 9460 18604 9512
rect 18656 9460 18662 9512
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 19337 9503 19395 9509
rect 19337 9500 19349 9503
rect 18932 9472 19349 9500
rect 18932 9460 18938 9472
rect 19337 9469 19349 9472
rect 19383 9469 19395 9503
rect 19337 9463 19395 9469
rect 19610 9460 19616 9512
rect 19668 9460 19674 9512
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23750 9500 23756 9512
rect 22971 9472 23756 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23750 9460 23756 9472
rect 23808 9460 23814 9512
rect 3973 9435 4031 9441
rect 3973 9432 3985 9435
rect 1596 9404 3985 9432
rect 3973 9401 3985 9404
rect 4019 9401 4031 9435
rect 23860 9432 23888 9528
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 25884 9509 25912 9608
rect 27246 9596 27252 9608
rect 27304 9596 27310 9648
rect 27632 9636 27660 9676
rect 28718 9664 28724 9676
rect 28776 9664 28782 9716
rect 30190 9664 30196 9716
rect 30248 9704 30254 9716
rect 31570 9704 31576 9716
rect 30248 9676 31576 9704
rect 30248 9664 30254 9676
rect 31570 9664 31576 9676
rect 31628 9664 31634 9716
rect 31846 9704 31852 9716
rect 31726 9676 31852 9704
rect 28997 9639 29055 9645
rect 27632 9608 27830 9636
rect 28997 9605 29009 9639
rect 29043 9636 29055 9639
rect 30098 9636 30104 9648
rect 29043 9608 30104 9636
rect 29043 9605 29055 9608
rect 28997 9599 29055 9605
rect 30098 9596 30104 9608
rect 30156 9596 30162 9648
rect 30742 9596 30748 9648
rect 30800 9596 30806 9648
rect 31478 9596 31484 9648
rect 31536 9636 31542 9648
rect 31726 9636 31754 9676
rect 31846 9664 31852 9676
rect 31904 9704 31910 9716
rect 32030 9704 32036 9716
rect 31904 9676 32036 9704
rect 31904 9664 31910 9676
rect 32030 9664 32036 9676
rect 32088 9664 32094 9716
rect 32306 9664 32312 9716
rect 32364 9704 32370 9716
rect 32953 9707 33011 9713
rect 32953 9704 32965 9707
rect 32364 9676 32965 9704
rect 32364 9664 32370 9676
rect 32953 9673 32965 9676
rect 32999 9673 33011 9707
rect 34882 9704 34888 9716
rect 32953 9667 33011 9673
rect 34532 9676 34888 9704
rect 31536 9608 31754 9636
rect 31536 9596 31542 9608
rect 32490 9596 32496 9648
rect 32548 9636 32554 9648
rect 34532 9636 34560 9676
rect 34882 9664 34888 9676
rect 34940 9664 34946 9716
rect 35158 9664 35164 9716
rect 35216 9704 35222 9716
rect 35621 9707 35679 9713
rect 35621 9704 35633 9707
rect 35216 9676 35633 9704
rect 35216 9664 35222 9676
rect 35621 9673 35633 9676
rect 35667 9673 35679 9707
rect 35621 9667 35679 9673
rect 35710 9664 35716 9716
rect 35768 9704 35774 9716
rect 36173 9707 36231 9713
rect 36173 9704 36185 9707
rect 35768 9676 36185 9704
rect 35768 9664 35774 9676
rect 36173 9673 36185 9676
rect 36219 9704 36231 9707
rect 36906 9704 36912 9716
rect 36219 9676 36912 9704
rect 36219 9673 36231 9676
rect 36173 9667 36231 9673
rect 36078 9636 36084 9648
rect 32548 9608 34560 9636
rect 35374 9608 36084 9636
rect 32548 9596 32554 9608
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 24949 9503 25007 9509
rect 24949 9500 24961 9503
rect 24360 9472 24961 9500
rect 24360 9460 24366 9472
rect 24949 9469 24961 9472
rect 24995 9469 25007 9503
rect 24949 9463 25007 9469
rect 25869 9503 25927 9509
rect 25869 9469 25881 9503
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 25958 9460 25964 9512
rect 26016 9460 26022 9512
rect 3973 9395 4031 9401
rect 22066 9404 23888 9432
rect 22066 9376 22094 9404
rect 25774 9392 25780 9444
rect 25832 9432 25838 9444
rect 26068 9432 26096 9531
rect 31662 9528 31668 9580
rect 31720 9568 31726 9580
rect 33888 9577 33916 9608
rect 36078 9596 36084 9608
rect 36136 9636 36142 9648
rect 36188 9636 36216 9667
rect 36906 9664 36912 9676
rect 36964 9664 36970 9716
rect 36136 9608 36216 9636
rect 49145 9639 49203 9645
rect 36136 9596 36142 9608
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 49326 9636 49332 9648
rect 49191 9608 49332 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 49326 9596 49332 9608
rect 49384 9596 49390 9648
rect 32861 9571 32919 9577
rect 32861 9568 32873 9571
rect 31720 9540 32873 9568
rect 31720 9528 31726 9540
rect 32861 9537 32873 9540
rect 32907 9537 32919 9571
rect 32861 9531 32919 9537
rect 33873 9571 33931 9577
rect 33873 9537 33885 9571
rect 33919 9537 33931 9571
rect 33873 9531 33931 9537
rect 47394 9528 47400 9580
rect 47452 9568 47458 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 47452 9540 47961 9568
rect 47452 9528 47458 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 27154 9460 27160 9512
rect 27212 9500 27218 9512
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27212 9472 27537 9500
rect 27212 9460 27218 9472
rect 27525 9469 27537 9472
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 28000 9472 29224 9500
rect 25832 9404 26096 9432
rect 26421 9435 26479 9441
rect 25832 9392 25838 9404
rect 26421 9401 26433 9435
rect 26467 9432 26479 9435
rect 28000 9432 28028 9472
rect 26467 9404 28028 9432
rect 29196 9432 29224 9472
rect 29270 9460 29276 9512
rect 29328 9500 29334 9512
rect 29546 9500 29552 9512
rect 29328 9472 29552 9500
rect 29328 9460 29334 9472
rect 29546 9460 29552 9472
rect 29604 9500 29610 9512
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29604 9472 29745 9500
rect 29604 9460 29610 9472
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 30009 9503 30067 9509
rect 30009 9500 30021 9503
rect 29733 9463 29791 9469
rect 29840 9472 30021 9500
rect 29196 9404 29500 9432
rect 26467 9401 26479 9404
rect 26421 9395 26479 9401
rect 2774 9324 2780 9376
rect 2832 9324 2838 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 14918 9364 14924 9376
rect 12943 9336 14924 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 18782 9364 18788 9376
rect 16080 9336 18788 9364
rect 16080 9324 16086 9336
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 19794 9324 19800 9376
rect 19852 9364 19858 9376
rect 21361 9367 21419 9373
rect 21361 9364 21373 9367
rect 19852 9336 21373 9364
rect 19852 9324 19858 9336
rect 21361 9333 21373 9336
rect 21407 9364 21419 9367
rect 21913 9367 21971 9373
rect 21913 9364 21925 9367
rect 21407 9336 21925 9364
rect 21407 9333 21419 9336
rect 21361 9327 21419 9333
rect 21913 9333 21925 9336
rect 21959 9364 21971 9367
rect 22002 9364 22008 9376
rect 21959 9336 22008 9364
rect 21959 9333 21971 9336
rect 21913 9327 21971 9333
rect 22002 9324 22008 9336
rect 22060 9336 22094 9376
rect 22060 9324 22066 9336
rect 22278 9324 22284 9376
rect 22336 9324 22342 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23750 9364 23756 9376
rect 23523 9336 23756 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 28810 9324 28816 9376
rect 28868 9364 28874 9376
rect 29270 9364 29276 9376
rect 28868 9336 29276 9364
rect 28868 9324 28874 9336
rect 29270 9324 29276 9336
rect 29328 9324 29334 9376
rect 29472 9364 29500 9404
rect 29638 9392 29644 9444
rect 29696 9432 29702 9444
rect 29840 9432 29868 9472
rect 30009 9469 30021 9472
rect 30055 9469 30067 9503
rect 30009 9463 30067 9469
rect 30098 9460 30104 9512
rect 30156 9500 30162 9512
rect 31481 9503 31539 9509
rect 31481 9500 31493 9503
rect 30156 9472 31493 9500
rect 30156 9460 30162 9472
rect 31481 9469 31493 9472
rect 31527 9469 31539 9503
rect 31481 9463 31539 9469
rect 29696 9404 29868 9432
rect 31496 9432 31524 9463
rect 31754 9460 31760 9512
rect 31812 9460 31818 9512
rect 31938 9460 31944 9512
rect 31996 9500 32002 9512
rect 32677 9503 32735 9509
rect 32677 9500 32689 9503
rect 31996 9472 32689 9500
rect 31996 9460 32002 9472
rect 32677 9469 32689 9472
rect 32723 9469 32735 9503
rect 32677 9463 32735 9469
rect 32766 9460 32772 9512
rect 32824 9500 32830 9512
rect 34149 9503 34207 9509
rect 34149 9500 34161 9503
rect 32824 9472 34161 9500
rect 32824 9460 32830 9472
rect 34149 9469 34161 9472
rect 34195 9500 34207 9503
rect 35894 9500 35900 9512
rect 34195 9472 35900 9500
rect 34195 9469 34207 9472
rect 34149 9463 34207 9469
rect 35894 9460 35900 9472
rect 35952 9460 35958 9512
rect 32214 9432 32220 9444
rect 31496 9404 32220 9432
rect 29696 9392 29702 9404
rect 32214 9392 32220 9404
rect 32272 9392 32278 9444
rect 30466 9364 30472 9376
rect 29472 9336 30472 9364
rect 30466 9324 30472 9336
rect 30524 9324 30530 9376
rect 31754 9324 31760 9376
rect 31812 9364 31818 9376
rect 32125 9367 32183 9373
rect 32125 9364 32137 9367
rect 31812 9336 32137 9364
rect 31812 9324 31818 9336
rect 32125 9333 32137 9336
rect 32171 9364 32183 9367
rect 32582 9364 32588 9376
rect 32171 9336 32588 9364
rect 32171 9333 32183 9336
rect 32125 9327 32183 9333
rect 32582 9324 32588 9336
rect 32640 9364 32646 9376
rect 33226 9364 33232 9376
rect 32640 9336 33232 9364
rect 32640 9324 32646 9336
rect 33226 9324 33232 9336
rect 33284 9324 33290 9376
rect 33321 9367 33379 9373
rect 33321 9333 33333 9367
rect 33367 9364 33379 9367
rect 35526 9364 35532 9376
rect 33367 9336 35532 9364
rect 33367 9333 33379 9336
rect 33321 9327 33379 9333
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 2222 9120 2228 9172
rect 2280 9120 2286 9172
rect 2682 9120 2688 9172
rect 2740 9120 2746 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 13814 9160 13820 9172
rect 2832 9132 13820 9160
rect 2832 9120 2838 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 16393 9163 16451 9169
rect 16393 9160 16405 9163
rect 15804 9132 16405 9160
rect 15804 9120 15810 9132
rect 16393 9129 16405 9132
rect 16439 9160 16451 9163
rect 17126 9160 17132 9172
rect 16439 9132 17132 9160
rect 16439 9129 16451 9132
rect 16393 9123 16451 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 19429 9163 19487 9169
rect 19429 9160 19441 9163
rect 17460 9132 19441 9160
rect 17460 9120 17466 9132
rect 19429 9129 19441 9132
rect 19475 9160 19487 9163
rect 19610 9160 19616 9172
rect 19475 9132 19616 9160
rect 19475 9129 19487 9132
rect 19429 9123 19487 9129
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22152 9132 22293 9160
rect 22152 9120 22158 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 22520 9132 24409 9160
rect 22520 9120 22526 9132
rect 24397 9129 24409 9132
rect 24443 9129 24455 9163
rect 24397 9123 24455 9129
rect 24673 9163 24731 9169
rect 24673 9129 24685 9163
rect 24719 9160 24731 9163
rect 25038 9160 25044 9172
rect 24719 9132 25044 9160
rect 24719 9129 24731 9132
rect 24673 9123 24731 9129
rect 25038 9120 25044 9132
rect 25096 9160 25102 9172
rect 25317 9163 25375 9169
rect 25317 9160 25329 9163
rect 25096 9132 25329 9160
rect 25096 9120 25102 9132
rect 25317 9129 25329 9132
rect 25363 9129 25375 9163
rect 25317 9123 25375 9129
rect 28905 9163 28963 9169
rect 28905 9129 28917 9163
rect 28951 9160 28963 9163
rect 32398 9160 32404 9172
rect 28951 9132 32404 9160
rect 28951 9129 28963 9132
rect 28905 9123 28963 9129
rect 32398 9120 32404 9132
rect 32456 9120 32462 9172
rect 32582 9120 32588 9172
rect 32640 9160 32646 9172
rect 32769 9163 32827 9169
rect 32769 9160 32781 9163
rect 32640 9132 32781 9160
rect 32640 9120 32646 9132
rect 32769 9129 32781 9132
rect 32815 9160 32827 9163
rect 32953 9163 33011 9169
rect 32953 9160 32965 9163
rect 32815 9132 32965 9160
rect 32815 9129 32827 9132
rect 32769 9123 32827 9129
rect 32953 9129 32965 9132
rect 32999 9129 33011 9163
rect 32953 9123 33011 9129
rect 34057 9163 34115 9169
rect 34057 9129 34069 9163
rect 34103 9160 34115 9163
rect 36354 9160 36360 9172
rect 34103 9132 36360 9160
rect 34103 9129 34115 9132
rect 34057 9123 34115 9129
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 36725 9163 36783 9169
rect 36725 9129 36737 9163
rect 36771 9160 36783 9163
rect 43714 9160 43720 9172
rect 36771 9132 43720 9160
rect 36771 9129 36783 9132
rect 36725 9123 36783 9129
rect 43714 9120 43720 9132
rect 43772 9120 43778 9172
rect 14461 9095 14519 9101
rect 14461 9061 14473 9095
rect 14507 9092 14519 9095
rect 15838 9092 15844 9104
rect 14507 9064 15844 9092
rect 14507 9061 14519 9064
rect 14461 9055 14519 9061
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 15933 9095 15991 9101
rect 15933 9061 15945 9095
rect 15979 9092 15991 9095
rect 16850 9092 16856 9104
rect 15979 9064 16856 9092
rect 15979 9061 15991 9064
rect 15933 9055 15991 9061
rect 16850 9052 16856 9064
rect 16908 9052 16914 9104
rect 29638 9052 29644 9104
rect 29696 9092 29702 9104
rect 30745 9095 30803 9101
rect 30745 9092 30757 9095
rect 29696 9064 30757 9092
rect 29696 9052 29702 9064
rect 30745 9061 30757 9064
rect 30791 9061 30803 9095
rect 33318 9092 33324 9104
rect 30745 9055 30803 9061
rect 32416 9064 33324 9092
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 2746 8996 3985 9024
rect 1302 8916 1308 8968
rect 1360 8956 1366 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1360 8928 1593 8956
rect 1360 8916 1366 8928
rect 1581 8925 1593 8928
rect 1627 8956 1639 8959
rect 2746 8956 2774 8996
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 12526 9024 12532 9036
rect 4120 8996 12532 9024
rect 4120 8984 4126 8996
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15160 8996 15301 9024
rect 15160 8984 15166 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15470 8984 15476 9036
rect 15528 8984 15534 9036
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 18141 9027 18199 9033
rect 18141 9024 18153 9027
rect 16540 8996 18153 9024
rect 16540 8984 16546 8996
rect 18141 8993 18153 8996
rect 18187 9024 18199 9027
rect 18874 9024 18880 9036
rect 18187 8996 18880 9024
rect 18187 8993 18199 8996
rect 18141 8987 18199 8993
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 19484 8996 20913 9024
rect 19484 8984 19490 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 23750 8984 23756 9036
rect 23808 8984 23814 9036
rect 24026 8984 24032 9036
rect 24084 8984 24090 9036
rect 28353 9027 28411 9033
rect 28353 8993 28365 9027
rect 28399 9024 28411 9027
rect 29656 9024 29684 9052
rect 28399 8996 29684 9024
rect 28399 8993 28411 8996
rect 28353 8987 28411 8993
rect 30190 8984 30196 9036
rect 30248 9024 30254 9036
rect 31478 9024 31484 9036
rect 30248 8996 31484 9024
rect 30248 8984 30254 8996
rect 31478 8984 31484 8996
rect 31536 8984 31542 9036
rect 32217 9027 32275 9033
rect 32217 8993 32229 9027
rect 32263 9024 32275 9027
rect 32416 9024 32444 9064
rect 33318 9052 33324 9064
rect 33376 9052 33382 9104
rect 35986 9052 35992 9104
rect 36044 9092 36050 9104
rect 39853 9095 39911 9101
rect 39853 9092 39865 9095
rect 36044 9064 39865 9092
rect 36044 9052 36050 9064
rect 32263 8996 32444 9024
rect 32263 8993 32275 8996
rect 32217 8987 32275 8993
rect 32490 8984 32496 9036
rect 32548 8984 32554 9036
rect 32766 8984 32772 9036
rect 32824 9024 32830 9036
rect 33042 9024 33048 9036
rect 32824 8996 33048 9024
rect 32824 8984 32830 8996
rect 33042 8984 33048 8996
rect 33100 9024 33106 9036
rect 33413 9027 33471 9033
rect 33413 9024 33425 9027
rect 33100 8996 33425 9024
rect 33100 8984 33106 8996
rect 33413 8993 33425 8996
rect 33459 8993 33471 9027
rect 33413 8987 33471 8993
rect 34238 8984 34244 9036
rect 34296 9024 34302 9036
rect 34333 9027 34391 9033
rect 34333 9024 34345 9027
rect 34296 8996 34345 9024
rect 34296 8984 34302 8996
rect 34333 8993 34345 8996
rect 34379 8993 34391 9027
rect 34333 8987 34391 8993
rect 34974 8984 34980 9036
rect 35032 8984 35038 9036
rect 35066 8984 35072 9036
rect 35124 9024 35130 9036
rect 35161 9027 35219 9033
rect 35161 9024 35173 9027
rect 35124 8996 35173 9024
rect 35124 8984 35130 8996
rect 35161 8993 35173 8996
rect 35207 8993 35219 9027
rect 35161 8987 35219 8993
rect 35526 8984 35532 9036
rect 35584 9024 35590 9036
rect 35584 8996 37688 9024
rect 35584 8984 35590 8996
rect 1627 8928 2774 8956
rect 3329 8959 3387 8965
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 3344 8888 3372 8919
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 12216 8928 14289 8956
rect 12216 8916 12222 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 15654 8956 15660 8968
rect 15611 8928 15660 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 18690 8916 18696 8968
rect 18748 8916 18754 8968
rect 19794 8916 19800 8968
rect 19852 8916 19858 8968
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8956 21235 8959
rect 21450 8956 21456 8968
rect 21223 8928 21456 8956
rect 21223 8925 21235 8928
rect 21177 8919 21235 8925
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8956 25651 8959
rect 25958 8956 25964 8968
rect 25639 8928 25964 8956
rect 25639 8925 25651 8928
rect 25593 8919 25651 8925
rect 25958 8916 25964 8928
rect 26016 8956 26022 8968
rect 30926 8956 30932 8968
rect 26016 8928 30932 8956
rect 26016 8916 26022 8928
rect 30926 8916 30932 8928
rect 30984 8916 30990 8968
rect 33597 8959 33655 8965
rect 33597 8925 33609 8959
rect 33643 8956 33655 8959
rect 33870 8956 33876 8968
rect 33643 8928 33876 8956
rect 33643 8925 33655 8928
rect 33597 8919 33655 8925
rect 33870 8916 33876 8928
rect 33928 8916 33934 8968
rect 34514 8916 34520 8968
rect 34572 8956 34578 8968
rect 37660 8965 37688 8996
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 34572 8928 36553 8956
rect 34572 8916 34578 8928
rect 36541 8925 36553 8928
rect 36587 8925 36599 8959
rect 36541 8919 36599 8925
rect 37645 8959 37703 8965
rect 37645 8925 37657 8959
rect 37691 8925 37703 8959
rect 37645 8919 37703 8925
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 1268 8860 3801 8888
rect 1268 8848 1274 8860
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 15286 8888 15292 8900
rect 3789 8851 3847 8857
rect 12406 8860 15292 8888
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 12406 8820 12434 8860
rect 15286 8848 15292 8860
rect 15344 8848 15350 8900
rect 16574 8848 16580 8900
rect 16632 8888 16638 8900
rect 16632 8860 16698 8888
rect 16632 8848 16638 8860
rect 17862 8848 17868 8900
rect 17920 8848 17926 8900
rect 22002 8848 22008 8900
rect 22060 8888 22066 8900
rect 28537 8891 28595 8897
rect 22060 8860 22586 8888
rect 23400 8860 24900 8888
rect 22060 8848 22066 8860
rect 2648 8792 12434 8820
rect 2648 8780 2654 8792
rect 14642 8780 14648 8832
rect 14700 8820 14706 8832
rect 14921 8823 14979 8829
rect 14921 8820 14933 8823
rect 14700 8792 14933 8820
rect 14700 8780 14706 8792
rect 14921 8789 14933 8792
rect 14967 8820 14979 8823
rect 16592 8820 16620 8848
rect 23400 8832 23428 8860
rect 24872 8832 24900 8860
rect 28537 8857 28549 8891
rect 28583 8888 28595 8891
rect 29733 8891 29791 8897
rect 29733 8888 29745 8891
rect 28583 8860 29745 8888
rect 28583 8857 28595 8860
rect 28537 8851 28595 8857
rect 29733 8857 29745 8860
rect 29779 8857 29791 8891
rect 29733 8851 29791 8857
rect 31754 8848 31760 8900
rect 31812 8848 31818 8900
rect 36446 8888 36452 8900
rect 32600 8860 36452 8888
rect 14967 8792 16620 8820
rect 21821 8823 21879 8829
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 21821 8789 21833 8823
rect 21867 8820 21879 8823
rect 22186 8820 22192 8832
rect 21867 8792 22192 8820
rect 21867 8789 21879 8792
rect 21821 8783 21879 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 23382 8780 23388 8832
rect 23440 8780 23446 8832
rect 24854 8780 24860 8832
rect 24912 8780 24918 8832
rect 25774 8780 25780 8832
rect 25832 8780 25838 8832
rect 27798 8780 27804 8832
rect 27856 8820 27862 8832
rect 28445 8823 28503 8829
rect 28445 8820 28457 8823
rect 27856 8792 28457 8820
rect 27856 8780 27862 8792
rect 28445 8789 28457 8792
rect 28491 8820 28503 8823
rect 30190 8820 30196 8832
rect 28491 8792 30196 8820
rect 28491 8789 28503 8792
rect 28445 8783 28503 8789
rect 30190 8780 30196 8792
rect 30248 8780 30254 8832
rect 30285 8823 30343 8829
rect 30285 8789 30297 8823
rect 30331 8820 30343 8823
rect 30742 8820 30748 8832
rect 30331 8792 30748 8820
rect 30331 8789 30343 8792
rect 30285 8783 30343 8789
rect 30742 8780 30748 8792
rect 30800 8780 30806 8832
rect 32122 8780 32128 8832
rect 32180 8820 32186 8832
rect 32600 8820 32628 8860
rect 36446 8848 36452 8860
rect 36504 8848 36510 8900
rect 39316 8897 39344 9064
rect 39853 9061 39865 9064
rect 39899 9061 39911 9095
rect 39853 9055 39911 9061
rect 49145 9027 49203 9033
rect 49145 8993 49157 9027
rect 49191 9024 49203 9027
rect 49234 9024 49240 9036
rect 49191 8996 49240 9024
rect 49191 8993 49203 8996
rect 49145 8987 49203 8993
rect 49234 8984 49240 8996
rect 49292 8984 49298 9036
rect 39390 8916 39396 8968
rect 39448 8956 39454 8968
rect 46474 8956 46480 8968
rect 39448 8928 46480 8956
rect 39448 8916 39454 8928
rect 46474 8916 46480 8928
rect 46532 8916 46538 8968
rect 47026 8916 47032 8968
rect 47084 8956 47090 8968
rect 47949 8959 48007 8965
rect 47949 8956 47961 8959
rect 47084 8928 47961 8956
rect 47084 8916 47090 8928
rect 47949 8925 47961 8928
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 39301 8891 39359 8897
rect 39301 8857 39313 8891
rect 39347 8857 39359 8891
rect 39301 8851 39359 8857
rect 39485 8891 39543 8897
rect 39485 8857 39497 8891
rect 39531 8888 39543 8891
rect 47578 8888 47584 8900
rect 39531 8860 47584 8888
rect 39531 8857 39543 8860
rect 39485 8851 39543 8857
rect 47578 8848 47584 8860
rect 47636 8848 47642 8900
rect 32180 8792 32628 8820
rect 33689 8823 33747 8829
rect 32180 8780 32186 8792
rect 33689 8789 33701 8823
rect 33735 8820 33747 8823
rect 34238 8820 34244 8832
rect 33735 8792 34244 8820
rect 33735 8789 33747 8792
rect 33689 8783 33747 8789
rect 34238 8780 34244 8792
rect 34296 8780 34302 8832
rect 35250 8780 35256 8832
rect 35308 8780 35314 8832
rect 35618 8780 35624 8832
rect 35676 8780 35682 8832
rect 37826 8780 37832 8832
rect 37884 8780 37890 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 3053 8619 3111 8625
rect 3053 8585 3065 8619
rect 3099 8616 3111 8619
rect 3099 8588 6914 8616
rect 3099 8585 3111 8588
rect 3053 8579 3111 8585
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2590 8480 2596 8492
rect 2179 8452 2596 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 2832 8452 2973 8480
rect 2832 8440 2838 8452
rect 2961 8449 2973 8452
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 2464 8384 3433 8412
rect 2464 8372 2470 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 6886 8412 6914 8588
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 15194 8616 15200 8628
rect 12768 8588 15200 8616
rect 12768 8576 12774 8588
rect 13648 8489 13676 8588
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 17494 8616 17500 8628
rect 16592 8588 17500 8616
rect 16592 8560 16620 8588
rect 17494 8576 17500 8588
rect 17552 8616 17558 8628
rect 17862 8616 17868 8628
rect 17552 8588 17868 8616
rect 17552 8576 17558 8588
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 19058 8576 19064 8628
rect 19116 8576 19122 8628
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 19886 8616 19892 8628
rect 19751 8588 19892 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21192 8588 22017 8616
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8548 13967 8551
rect 14182 8548 14188 8560
rect 13955 8520 14188 8548
rect 13955 8517 13967 8520
rect 13909 8511 13967 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 15749 8551 15807 8557
rect 15749 8548 15761 8551
rect 15134 8520 15761 8548
rect 15749 8517 15761 8520
rect 15795 8548 15807 8551
rect 16209 8551 16267 8557
rect 16209 8548 16221 8551
rect 15795 8520 16221 8548
rect 15795 8517 15807 8520
rect 15749 8511 15807 8517
rect 16209 8517 16221 8520
rect 16255 8548 16267 8551
rect 16574 8548 16580 8560
rect 16255 8520 16580 8548
rect 16255 8517 16267 8520
rect 16209 8511 16267 8517
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17126 8548 17132 8560
rect 16816 8520 17132 8548
rect 16816 8508 16822 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17512 8548 17540 8576
rect 17512 8520 17618 8548
rect 19794 8508 19800 8560
rect 19852 8548 19858 8560
rect 21192 8557 21220 8588
rect 21177 8551 21235 8557
rect 19852 8520 20010 8548
rect 19852 8508 19858 8520
rect 21177 8517 21189 8551
rect 21223 8517 21235 8551
rect 21177 8511 21235 8517
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 16482 8480 16488 8492
rect 15252 8452 16488 8480
rect 15252 8440 15258 8452
rect 16482 8440 16488 8452
rect 16540 8480 16546 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16540 8452 16865 8480
rect 16540 8440 16546 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 6886 8384 15056 8412
rect 3421 8375 3479 8381
rect 15028 8344 15056 8384
rect 15102 8372 15108 8424
rect 15160 8412 15166 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15160 8384 15393 8412
rect 15160 8372 15166 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 17218 8412 17224 8424
rect 16448 8384 17224 8412
rect 16448 8372 16454 8384
rect 17218 8372 17224 8384
rect 17276 8412 17282 8424
rect 21174 8412 21180 8424
rect 17276 8384 21180 8412
rect 17276 8372 17282 8384
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 21450 8372 21456 8424
rect 21508 8372 21514 8424
rect 16666 8344 16672 8356
rect 15028 8316 16672 8344
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 21928 8344 21956 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 22388 8588 23152 8616
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 22388 8480 22416 8588
rect 23124 8548 23152 8588
rect 30466 8576 30472 8628
rect 30524 8616 30530 8628
rect 31297 8619 31355 8625
rect 31297 8616 31309 8619
rect 30524 8588 31309 8616
rect 30524 8576 30530 8588
rect 31297 8585 31309 8588
rect 31343 8585 31355 8619
rect 31297 8579 31355 8585
rect 31757 8619 31815 8625
rect 31757 8585 31769 8619
rect 31803 8616 31815 8619
rect 32122 8616 32128 8628
rect 31803 8588 32128 8616
rect 31803 8585 31815 8588
rect 31757 8579 31815 8585
rect 32122 8576 32128 8588
rect 32180 8576 32186 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32548 8588 32996 8616
rect 32548 8576 32554 8588
rect 24121 8551 24179 8557
rect 24121 8548 24133 8551
rect 23046 8520 24133 8548
rect 24121 8517 24133 8520
rect 24167 8517 24179 8551
rect 24121 8511 24179 8517
rect 29086 8508 29092 8560
rect 29144 8508 29150 8560
rect 30742 8548 30748 8560
rect 30314 8520 30748 8548
rect 30742 8508 30748 8520
rect 30800 8508 30806 8560
rect 32582 8548 32588 8560
rect 30852 8520 32588 8548
rect 22060 8466 22416 8480
rect 23753 8483 23811 8489
rect 22060 8452 22402 8466
rect 22060 8440 22066 8452
rect 23753 8449 23765 8483
rect 23799 8480 23811 8483
rect 24026 8480 24032 8492
rect 23799 8452 24032 8480
rect 23799 8449 23811 8452
rect 23753 8443 23811 8449
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 23477 8415 23535 8421
rect 23477 8412 23489 8415
rect 22152 8384 23489 8412
rect 22152 8372 22158 8384
rect 23477 8381 23489 8384
rect 23523 8381 23535 8415
rect 23477 8375 23535 8381
rect 28810 8372 28816 8424
rect 28868 8372 28874 8424
rect 30852 8412 30880 8520
rect 32582 8508 32588 8520
rect 32640 8508 32646 8560
rect 32968 8548 32996 8588
rect 33318 8576 33324 8628
rect 33376 8616 33382 8628
rect 34057 8619 34115 8625
rect 34057 8616 34069 8619
rect 33376 8588 34069 8616
rect 33376 8576 33382 8588
rect 34057 8585 34069 8588
rect 34103 8616 34115 8619
rect 34974 8616 34980 8628
rect 34103 8588 34980 8616
rect 34103 8585 34115 8588
rect 34057 8579 34115 8585
rect 34974 8576 34980 8588
rect 35032 8576 35038 8628
rect 37645 8619 37703 8625
rect 37645 8585 37657 8619
rect 37691 8616 37703 8619
rect 40034 8616 40040 8628
rect 37691 8588 40040 8616
rect 37691 8585 37703 8588
rect 37645 8579 37703 8585
rect 40034 8576 40040 8588
rect 40092 8576 40098 8628
rect 32968 8520 33074 8548
rect 33870 8508 33876 8560
rect 33928 8548 33934 8560
rect 34330 8548 34336 8560
rect 33928 8520 34336 8548
rect 33928 8508 33934 8520
rect 34330 8508 34336 8520
rect 34388 8548 34394 8560
rect 34388 8520 34468 8548
rect 34388 8508 34394 8520
rect 31110 8440 31116 8492
rect 31168 8480 31174 8492
rect 31389 8483 31447 8489
rect 31389 8480 31401 8483
rect 31168 8452 31401 8480
rect 31168 8440 31174 8452
rect 31389 8449 31401 8452
rect 31435 8449 31447 8483
rect 31389 8443 31447 8449
rect 32306 8440 32312 8492
rect 32364 8440 32370 8492
rect 28920 8384 30880 8412
rect 31205 8415 31263 8421
rect 22462 8344 22468 8356
rect 21928 8316 22468 8344
rect 22462 8304 22468 8316
rect 22520 8304 22526 8356
rect 24854 8304 24860 8356
rect 24912 8344 24918 8356
rect 28920 8344 28948 8384
rect 31205 8381 31217 8415
rect 31251 8412 31263 8415
rect 31846 8412 31852 8424
rect 31251 8384 31852 8412
rect 31251 8381 31263 8384
rect 31205 8375 31263 8381
rect 31846 8372 31852 8384
rect 31904 8372 31910 8424
rect 32214 8372 32220 8424
rect 32272 8412 32278 8424
rect 32585 8415 32643 8421
rect 32585 8412 32597 8415
rect 32272 8384 32597 8412
rect 32272 8372 32278 8384
rect 32585 8381 32597 8384
rect 32631 8412 32643 8415
rect 32950 8412 32956 8424
rect 32631 8384 32956 8412
rect 32631 8381 32643 8384
rect 32585 8375 32643 8381
rect 32950 8372 32956 8384
rect 33008 8372 33014 8424
rect 33042 8372 33048 8424
rect 33100 8412 33106 8424
rect 34333 8415 34391 8421
rect 34333 8412 34345 8415
rect 33100 8384 34345 8412
rect 33100 8372 33106 8384
rect 34333 8381 34345 8384
rect 34379 8381 34391 8415
rect 34440 8412 34468 8520
rect 35618 8508 35624 8560
rect 35676 8548 35682 8560
rect 35676 8520 37596 8548
rect 35676 8508 35682 8520
rect 34793 8483 34851 8489
rect 34793 8449 34805 8483
rect 34839 8480 34851 8483
rect 36078 8480 36084 8492
rect 34839 8452 36084 8480
rect 34839 8449 34851 8452
rect 34793 8443 34851 8449
rect 36078 8440 36084 8452
rect 36136 8440 36142 8492
rect 36814 8440 36820 8492
rect 36872 8480 36878 8492
rect 37461 8483 37519 8489
rect 37461 8480 37473 8483
rect 36872 8452 37473 8480
rect 36872 8440 36878 8452
rect 37461 8449 37473 8452
rect 37507 8449 37519 8483
rect 37568 8480 37596 8520
rect 37826 8508 37832 8560
rect 37884 8548 37890 8560
rect 44177 8551 44235 8557
rect 44177 8548 44189 8551
rect 37884 8520 44189 8548
rect 37884 8508 37890 8520
rect 44177 8517 44189 8520
rect 44223 8517 44235 8551
rect 44177 8511 44235 8517
rect 44361 8551 44419 8557
rect 44361 8517 44373 8551
rect 44407 8548 44419 8551
rect 47762 8548 47768 8560
rect 44407 8520 47768 8548
rect 44407 8517 44419 8520
rect 44361 8511 44419 8517
rect 47762 8508 47768 8520
rect 47820 8508 47826 8560
rect 49142 8508 49148 8560
rect 49200 8508 49206 8560
rect 38933 8483 38991 8489
rect 38933 8480 38945 8483
rect 37568 8452 38945 8480
rect 37461 8443 37519 8449
rect 38933 8449 38945 8452
rect 38979 8449 38991 8483
rect 38933 8443 38991 8449
rect 40310 8440 40316 8492
rect 40368 8480 40374 8492
rect 40773 8483 40831 8489
rect 40773 8480 40785 8483
rect 40368 8452 40785 8480
rect 40368 8440 40374 8452
rect 40773 8449 40785 8452
rect 40819 8449 40831 8483
rect 40773 8443 40831 8449
rect 45830 8440 45836 8492
rect 45888 8440 45894 8492
rect 46750 8440 46756 8492
rect 46808 8480 46814 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46808 8452 47961 8480
rect 46808 8440 46814 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 34609 8415 34667 8421
rect 34609 8412 34621 8415
rect 34440 8384 34621 8412
rect 34333 8375 34391 8381
rect 34609 8381 34621 8384
rect 34655 8412 34667 8415
rect 39390 8412 39396 8424
rect 34655 8384 39396 8412
rect 34655 8381 34667 8384
rect 34609 8375 34667 8381
rect 39390 8372 39396 8384
rect 39448 8372 39454 8424
rect 40497 8415 40555 8421
rect 40497 8381 40509 8415
rect 40543 8412 40555 8415
rect 40543 8384 45554 8412
rect 40543 8381 40555 8384
rect 40497 8375 40555 8381
rect 24912 8316 28948 8344
rect 30561 8347 30619 8353
rect 24912 8304 24918 8316
rect 30561 8313 30573 8347
rect 30607 8344 30619 8347
rect 31938 8344 31944 8356
rect 30607 8316 31944 8344
rect 30607 8313 30619 8316
rect 30561 8307 30619 8313
rect 31938 8304 31944 8316
rect 31996 8304 32002 8356
rect 38746 8344 38752 8356
rect 38626 8316 38752 8344
rect 32030 8236 32036 8288
rect 32088 8276 32094 8288
rect 38626 8276 38654 8316
rect 38746 8304 38752 8316
rect 38804 8304 38810 8356
rect 39117 8347 39175 8353
rect 39117 8313 39129 8347
rect 39163 8344 39175 8347
rect 44910 8344 44916 8356
rect 39163 8316 44916 8344
rect 39163 8313 39175 8316
rect 39117 8307 39175 8313
rect 44910 8304 44916 8316
rect 44968 8304 44974 8356
rect 45526 8344 45554 8384
rect 46842 8372 46848 8424
rect 46900 8372 46906 8424
rect 47670 8344 47676 8356
rect 45526 8316 47676 8344
rect 47670 8304 47676 8316
rect 47728 8304 47734 8356
rect 32088 8248 38654 8276
rect 32088 8236 32094 8248
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 2225 8075 2283 8081
rect 2225 8041 2237 8075
rect 2271 8072 2283 8075
rect 2774 8072 2780 8084
rect 2271 8044 2780 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 18564 8044 18981 8072
rect 18564 8032 18570 8044
rect 18969 8041 18981 8044
rect 19015 8041 19027 8075
rect 18969 8035 19027 8041
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22005 8075 22063 8081
rect 22005 8072 22017 8075
rect 21968 8044 22017 8072
rect 21968 8032 21974 8044
rect 22005 8041 22017 8044
rect 22051 8041 22063 8075
rect 22005 8035 22063 8041
rect 30377 8075 30435 8081
rect 30377 8041 30389 8075
rect 30423 8072 30435 8075
rect 30558 8072 30564 8084
rect 30423 8044 30564 8072
rect 30423 8041 30435 8044
rect 30377 8035 30435 8041
rect 30558 8032 30564 8044
rect 30616 8032 30622 8084
rect 31757 8075 31815 8081
rect 31757 8041 31769 8075
rect 31803 8072 31815 8075
rect 35250 8072 35256 8084
rect 31803 8044 35256 8072
rect 31803 8041 31815 8044
rect 31757 8035 31815 8041
rect 35250 8032 35256 8044
rect 35308 8032 35314 8084
rect 15749 8007 15807 8013
rect 15749 7973 15761 8007
rect 15795 8004 15807 8007
rect 18874 8004 18880 8016
rect 15795 7976 18880 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 18874 7964 18880 7976
rect 18932 7964 18938 8016
rect 27522 7964 27528 8016
rect 27580 8004 27586 8016
rect 37553 8007 37611 8013
rect 37553 8004 37565 8007
rect 27580 7976 37565 8004
rect 27580 7964 27586 7976
rect 37553 7973 37565 7976
rect 37599 7973 37611 8007
rect 37553 7967 37611 7973
rect 3237 7939 3295 7945
rect 3237 7936 3249 7939
rect 1596 7908 3249 7936
rect 1596 7880 1624 7908
rect 3237 7905 3249 7908
rect 3283 7905 3295 7939
rect 3237 7899 3295 7905
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 16390 7936 16396 7948
rect 3568 7908 16396 7936
rect 3568 7896 3574 7908
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16758 7896 16764 7948
rect 16816 7896 16822 7948
rect 16942 7896 16948 7948
rect 17000 7896 17006 7948
rect 18049 7939 18107 7945
rect 18049 7905 18061 7939
rect 18095 7936 18107 7939
rect 18598 7936 18604 7948
rect 18095 7908 18604 7936
rect 18095 7905 18107 7908
rect 18049 7899 18107 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 19944 7908 20913 7936
rect 19944 7896 19950 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7936 22707 7939
rect 23566 7936 23572 7948
rect 22695 7908 23572 7936
rect 22695 7905 22707 7908
rect 22649 7899 22707 7905
rect 23566 7896 23572 7908
rect 23624 7896 23630 7948
rect 29914 7896 29920 7948
rect 29972 7896 29978 7948
rect 31205 7939 31263 7945
rect 31205 7905 31217 7939
rect 31251 7936 31263 7939
rect 32214 7936 32220 7948
rect 31251 7908 32220 7936
rect 31251 7905 31263 7908
rect 31205 7899 31263 7905
rect 32214 7896 32220 7908
rect 32272 7896 32278 7948
rect 32493 7939 32551 7945
rect 32493 7905 32505 7939
rect 32539 7936 32551 7939
rect 33413 7939 33471 7945
rect 33413 7936 33425 7939
rect 32539 7908 33425 7936
rect 32539 7905 32551 7908
rect 32493 7899 32551 7905
rect 33413 7905 33425 7908
rect 33459 7936 33471 7939
rect 34606 7936 34612 7948
rect 33459 7908 34612 7936
rect 33459 7905 33471 7908
rect 33413 7899 33471 7905
rect 34606 7896 34612 7908
rect 34664 7896 34670 7948
rect 1578 7828 1584 7880
rect 1636 7828 1642 7880
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2280 7840 2697 7868
rect 2280 7828 2286 7840
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 14976 7840 15577 7868
rect 14976 7828 14982 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7868 17095 7871
rect 18322 7868 18328 7880
rect 17083 7840 18328 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 19794 7828 19800 7880
rect 19852 7828 19858 7880
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 21450 7868 21456 7880
rect 21223 7840 21456 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 14366 7800 14372 7812
rect 2884 7772 14372 7800
rect 2884 7741 2912 7772
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 17420 7772 18245 7800
rect 17420 7741 17448 7772
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 19610 7800 19616 7812
rect 18233 7763 18291 7769
rect 18616 7772 19616 7800
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 17405 7735 17463 7741
rect 17405 7701 17417 7735
rect 17451 7701 17463 7735
rect 17405 7695 17463 7701
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18414 7732 18420 7744
rect 18187 7704 18420 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 18616 7741 18644 7772
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 20990 7760 20996 7812
rect 21048 7800 21054 7812
rect 21192 7800 21220 7831
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22244 7840 22385 7868
rect 22244 7828 22250 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 30558 7828 30564 7880
rect 30616 7868 30622 7880
rect 31297 7871 31355 7877
rect 31297 7868 31309 7871
rect 30616 7840 31309 7868
rect 30616 7828 30622 7840
rect 31297 7837 31309 7840
rect 31343 7837 31355 7871
rect 31297 7831 31355 7837
rect 32674 7828 32680 7880
rect 32732 7828 32738 7880
rect 37568 7868 37596 7967
rect 49145 7939 49203 7945
rect 49145 7905 49157 7939
rect 49191 7936 49203 7939
rect 49326 7936 49332 7948
rect 49191 7908 49332 7936
rect 49191 7905 49203 7908
rect 49145 7899 49203 7905
rect 49326 7896 49332 7908
rect 49384 7896 49390 7948
rect 38013 7871 38071 7877
rect 38013 7868 38025 7871
rect 37568 7840 38025 7868
rect 38013 7837 38025 7840
rect 38059 7837 38071 7871
rect 39022 7868 39028 7880
rect 38013 7831 38071 7837
rect 38120 7840 39028 7868
rect 21048 7772 21220 7800
rect 21048 7760 21054 7772
rect 21266 7760 21272 7812
rect 21324 7800 21330 7812
rect 21324 7772 22094 7800
rect 21324 7760 21330 7772
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7701 18659 7735
rect 18601 7695 18659 7701
rect 21450 7692 21456 7744
rect 21508 7732 21514 7744
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21508 7704 21649 7732
rect 21508 7692 21514 7704
rect 21637 7701 21649 7704
rect 21683 7701 21695 7735
rect 22066 7732 22094 7772
rect 30742 7760 30748 7812
rect 30800 7800 30806 7812
rect 31662 7800 31668 7812
rect 30800 7772 31668 7800
rect 30800 7760 30806 7772
rect 31662 7760 31668 7772
rect 31720 7800 31726 7812
rect 31754 7800 31760 7812
rect 31720 7772 31760 7800
rect 31720 7760 31726 7772
rect 31754 7760 31760 7772
rect 31812 7760 31818 7812
rect 38120 7800 38148 7840
rect 39022 7828 39028 7840
rect 39080 7828 39086 7880
rect 46934 7828 46940 7880
rect 46992 7868 46998 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 46992 7840 47961 7868
rect 46992 7828 46998 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 33060 7772 38148 7800
rect 22465 7735 22523 7741
rect 22465 7732 22477 7735
rect 22066 7704 22477 7732
rect 21637 7695 21695 7701
rect 22465 7701 22477 7704
rect 22511 7732 22523 7735
rect 23109 7735 23167 7741
rect 23109 7732 23121 7735
rect 22511 7704 23121 7732
rect 22511 7701 22523 7704
rect 22465 7695 22523 7701
rect 23109 7701 23121 7704
rect 23155 7732 23167 7735
rect 25774 7732 25780 7744
rect 23155 7704 25780 7732
rect 23155 7701 23167 7704
rect 23109 7695 23167 7701
rect 25774 7692 25780 7704
rect 25832 7692 25838 7744
rect 30466 7692 30472 7744
rect 30524 7692 30530 7744
rect 31386 7692 31392 7744
rect 31444 7692 31450 7744
rect 32582 7692 32588 7744
rect 32640 7692 32646 7744
rect 33060 7741 33088 7772
rect 38746 7760 38752 7812
rect 38804 7760 38810 7812
rect 38933 7803 38991 7809
rect 38933 7769 38945 7803
rect 38979 7800 38991 7803
rect 40586 7800 40592 7812
rect 38979 7772 40592 7800
rect 38979 7769 38991 7772
rect 38933 7763 38991 7769
rect 40586 7760 40592 7772
rect 40644 7760 40650 7812
rect 33045 7735 33103 7741
rect 33045 7701 33057 7735
rect 33091 7701 33103 7735
rect 33045 7695 33103 7701
rect 38105 7735 38163 7741
rect 38105 7701 38117 7735
rect 38151 7732 38163 7735
rect 38654 7732 38660 7744
rect 38151 7704 38660 7732
rect 38151 7701 38163 7704
rect 38105 7695 38163 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 38764 7732 38792 7760
rect 39209 7735 39267 7741
rect 39209 7732 39221 7735
rect 38764 7704 39221 7732
rect 39209 7701 39221 7704
rect 39255 7701 39267 7735
rect 39209 7695 39267 7701
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 2222 7488 2228 7540
rect 2280 7488 2286 7540
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 21266 7528 21272 7540
rect 3660 7500 21272 7528
rect 3660 7488 3666 7500
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 22278 7488 22284 7540
rect 22336 7528 22342 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22336 7500 22477 7528
rect 22336 7488 22342 7500
rect 22465 7497 22477 7500
rect 22511 7528 22523 7531
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22511 7500 23029 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 31110 7488 31116 7540
rect 31168 7488 31174 7540
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 32309 7531 32367 7537
rect 32309 7528 32321 7531
rect 31444 7500 32321 7528
rect 31444 7488 31450 7500
rect 32309 7497 32321 7500
rect 32355 7497 32367 7531
rect 39025 7531 39083 7537
rect 39025 7528 39037 7531
rect 32309 7491 32367 7497
rect 38580 7500 39037 7528
rect 3789 7463 3847 7469
rect 3789 7460 3801 7463
rect 2746 7432 3801 7460
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1360 7364 1593 7392
rect 1360 7352 1366 7364
rect 1581 7361 1593 7364
rect 1627 7392 1639 7395
rect 2746 7392 2774 7432
rect 3789 7429 3801 7432
rect 3835 7429 3847 7463
rect 3789 7423 3847 7429
rect 21174 7420 21180 7472
rect 21232 7460 21238 7472
rect 21361 7463 21419 7469
rect 21361 7460 21373 7463
rect 21232 7432 21373 7460
rect 21232 7420 21238 7432
rect 21361 7429 21373 7432
rect 21407 7429 21419 7463
rect 21361 7423 21419 7429
rect 1627 7364 2774 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 3326 7352 3332 7404
rect 3384 7392 3390 7404
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 3384 7364 3617 7392
rect 3384 7352 3390 7364
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 18012 7364 18245 7392
rect 18012 7352 18018 7364
rect 18233 7361 18245 7364
rect 18279 7392 18291 7395
rect 18693 7395 18751 7401
rect 18693 7392 18705 7395
rect 18279 7364 18705 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18693 7361 18705 7364
rect 18739 7392 18751 7395
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18739 7364 18981 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 18969 7361 18981 7364
rect 19015 7392 19027 7395
rect 19794 7392 19800 7404
rect 19015 7364 19800 7392
rect 19015 7361 19027 7364
rect 18969 7355 19027 7361
rect 19794 7352 19800 7364
rect 19852 7392 19858 7404
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 19852 7364 21281 7392
rect 19852 7352 19858 7364
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21376 7392 21404 7423
rect 31846 7420 31852 7472
rect 31904 7460 31910 7472
rect 32766 7460 32772 7472
rect 31904 7432 32772 7460
rect 31904 7420 31910 7432
rect 32766 7420 32772 7432
rect 32824 7420 32830 7472
rect 34422 7420 34428 7472
rect 34480 7460 34486 7472
rect 38580 7469 38608 7500
rect 39025 7497 39037 7500
rect 39071 7497 39083 7531
rect 39025 7491 39083 7497
rect 38565 7463 38623 7469
rect 38565 7460 38577 7463
rect 34480 7432 38577 7460
rect 34480 7420 34486 7432
rect 38565 7429 38577 7432
rect 38611 7429 38623 7463
rect 38565 7423 38623 7429
rect 38654 7420 38660 7472
rect 38712 7460 38718 7472
rect 46934 7460 46940 7472
rect 38712 7432 46940 7460
rect 38712 7420 38718 7432
rect 46934 7420 46940 7432
rect 46992 7420 46998 7472
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 49234 7460 49240 7472
rect 49191 7432 49240 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 49234 7420 49240 7432
rect 49292 7420 49298 7472
rect 22373 7395 22431 7401
rect 22373 7392 22385 7395
rect 21376 7364 22385 7392
rect 21269 7355 21327 7361
rect 22373 7361 22385 7364
rect 22419 7392 22431 7395
rect 30466 7392 30472 7404
rect 22419 7364 30472 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 21284 7324 21312 7355
rect 30466 7352 30472 7364
rect 30524 7352 30530 7404
rect 37829 7395 37887 7401
rect 37829 7392 37841 7395
rect 37384 7364 37841 7392
rect 21450 7324 21456 7336
rect 21284 7296 21456 7324
rect 21450 7284 21456 7296
rect 21508 7324 21514 7336
rect 21545 7327 21603 7333
rect 21545 7324 21557 7327
rect 21508 7296 21557 7324
rect 21508 7284 21514 7296
rect 21545 7293 21557 7296
rect 21591 7293 21603 7327
rect 21545 7287 21603 7293
rect 22554 7284 22560 7336
rect 22612 7284 22618 7336
rect 20714 7216 20720 7268
rect 20772 7256 20778 7268
rect 22005 7259 22063 7265
rect 22005 7256 22017 7259
rect 20772 7228 22017 7256
rect 20772 7216 20778 7228
rect 22005 7225 22017 7228
rect 22051 7225 22063 7259
rect 22005 7219 22063 7225
rect 28626 7216 28632 7268
rect 28684 7256 28690 7268
rect 37384 7265 37412 7364
rect 37829 7361 37841 7364
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 44910 7352 44916 7404
rect 44968 7352 44974 7404
rect 47118 7352 47124 7404
rect 47176 7392 47182 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 47176 7364 47961 7392
rect 47176 7352 47182 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 37369 7259 37427 7265
rect 37369 7256 37381 7259
rect 28684 7228 37381 7256
rect 28684 7216 28690 7228
rect 37369 7225 37381 7228
rect 37415 7225 37427 7259
rect 37369 7219 37427 7225
rect 38749 7259 38807 7265
rect 38749 7225 38761 7259
rect 38795 7256 38807 7259
rect 45097 7259 45155 7265
rect 38795 7228 42104 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 2774 7188 2780 7200
rect 2731 7160 2780 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 32582 7148 32588 7200
rect 32640 7188 32646 7200
rect 32861 7191 32919 7197
rect 32861 7188 32873 7191
rect 32640 7160 32873 7188
rect 32640 7148 32646 7160
rect 32861 7157 32873 7160
rect 32907 7188 32919 7191
rect 37274 7188 37280 7200
rect 32907 7160 37280 7188
rect 32907 7157 32919 7160
rect 32861 7151 32919 7157
rect 37274 7148 37280 7160
rect 37332 7148 37338 7200
rect 37918 7148 37924 7200
rect 37976 7148 37982 7200
rect 42076 7188 42104 7228
rect 45097 7225 45109 7259
rect 45143 7256 45155 7259
rect 47854 7256 47860 7268
rect 45143 7228 47860 7256
rect 45143 7225 45155 7228
rect 45097 7219 45155 7225
rect 47854 7216 47860 7228
rect 47912 7216 47918 7268
rect 45738 7188 45744 7200
rect 42076 7160 45744 7188
rect 45738 7148 45744 7160
rect 45796 7148 45802 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 30466 6944 30472 6996
rect 30524 6984 30530 6996
rect 38470 6984 38476 6996
rect 30524 6956 38476 6984
rect 30524 6944 30530 6956
rect 38470 6944 38476 6956
rect 38528 6944 38534 6996
rect 37918 6876 37924 6928
rect 37976 6916 37982 6928
rect 47026 6916 47032 6928
rect 37976 6888 47032 6916
rect 37976 6876 37982 6888
rect 47026 6876 47032 6888
rect 47084 6876 47090 6928
rect 3237 6851 3295 6857
rect 3237 6848 3249 6851
rect 1596 6820 3249 6848
rect 1596 6792 1624 6820
rect 3237 6817 3249 6820
rect 3283 6817 3295 6851
rect 3237 6811 3295 6817
rect 49142 6808 49148 6860
rect 49200 6808 49206 6860
rect 1578 6740 1584 6792
rect 1636 6740 1642 6792
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2271 6752 2697 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 2685 6743 2743 6749
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6780 4031 6783
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 4019 6752 4445 6780
rect 4019 6749 4031 6752
rect 3973 6743 4031 6749
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 3988 6712 4016 6743
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 16908 6752 17693 6780
rect 16908 6740 16914 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 40586 6740 40592 6792
rect 40644 6780 40650 6792
rect 46109 6783 46167 6789
rect 46109 6780 46121 6783
rect 40644 6752 46121 6780
rect 40644 6740 40650 6752
rect 46109 6749 46121 6752
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 47762 6740 47768 6792
rect 47820 6780 47826 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47820 6752 47961 6780
rect 47820 6740 47826 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 10594 6712 10600 6724
rect 1360 6684 4016 6712
rect 4172 6684 10600 6712
rect 1360 6672 1366 6684
rect 2866 6604 2872 6656
rect 2924 6604 2930 6656
rect 4172 6653 4200 6684
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 47305 6715 47363 6721
rect 47305 6681 47317 6715
rect 47351 6712 47363 6715
rect 48682 6712 48688 6724
rect 47351 6684 48688 6712
rect 47351 6681 47363 6684
rect 47305 6675 47363 6681
rect 48682 6672 48688 6684
rect 48740 6672 48746 6724
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6613 4215 6647
rect 4157 6607 4215 6613
rect 17865 6647 17923 6653
rect 17865 6613 17877 6647
rect 17911 6644 17923 6647
rect 19242 6644 19248 6656
rect 17911 6616 19248 6644
rect 17911 6613 17923 6616
rect 17865 6607 17923 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19797 6647 19855 6653
rect 19797 6613 19809 6647
rect 19843 6644 19855 6647
rect 21910 6644 21916 6656
rect 19843 6616 21916 6644
rect 19843 6613 19855 6616
rect 19797 6607 19855 6613
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 2774 6332 2780 6384
rect 2832 6332 2838 6384
rect 2961 6375 3019 6381
rect 2961 6341 2973 6375
rect 3007 6372 3019 6375
rect 27798 6372 27804 6384
rect 3007 6344 27804 6372
rect 3007 6341 3019 6344
rect 2961 6335 3019 6341
rect 27798 6332 27804 6344
rect 27856 6332 27862 6384
rect 30834 6332 30840 6384
rect 30892 6372 30898 6384
rect 37553 6375 37611 6381
rect 37553 6372 37565 6375
rect 30892 6344 37565 6372
rect 30892 6332 30898 6344
rect 37553 6341 37565 6344
rect 37599 6372 37611 6375
rect 38013 6375 38071 6381
rect 38013 6372 38025 6375
rect 37599 6344 38025 6372
rect 37599 6341 37611 6344
rect 37553 6335 37611 6341
rect 38013 6341 38025 6344
rect 38059 6341 38071 6375
rect 38013 6335 38071 6341
rect 40034 6332 40040 6384
rect 40092 6372 40098 6384
rect 43993 6375 44051 6381
rect 43993 6372 44005 6375
rect 40092 6344 44005 6372
rect 40092 6332 40098 6344
rect 43993 6341 44005 6344
rect 44039 6341 44051 6375
rect 43993 6335 44051 6341
rect 49145 6375 49203 6381
rect 49145 6341 49157 6375
rect 49191 6372 49203 6375
rect 49326 6372 49332 6384
rect 49191 6344 49332 6372
rect 49191 6341 49203 6344
rect 49145 6335 49203 6341
rect 49326 6332 49332 6344
rect 49384 6332 49390 6384
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6304 2283 6307
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 2271 6276 3433 6304
rect 2271 6273 2283 6276
rect 2225 6267 2283 6273
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 1596 6236 1624 6267
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 23934 6304 23940 6316
rect 11020 6276 23940 6304
rect 11020 6264 11026 6276
rect 23934 6264 23940 6276
rect 23992 6264 23998 6316
rect 27062 6264 27068 6316
rect 27120 6304 27126 6316
rect 36814 6304 36820 6316
rect 27120 6276 36820 6304
rect 27120 6264 27126 6276
rect 36814 6264 36820 6276
rect 36872 6264 36878 6316
rect 36998 6264 37004 6316
rect 37056 6304 37062 6316
rect 47210 6304 47216 6316
rect 37056 6276 47216 6304
rect 37056 6264 37062 6276
rect 47210 6264 47216 6276
rect 47268 6264 47274 6316
rect 47578 6264 47584 6316
rect 47636 6304 47642 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 47636 6276 47961 6304
rect 47636 6264 47642 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 1596 6208 3985 6236
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 15838 6196 15844 6248
rect 15896 6236 15902 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 15896 6208 18061 6236
rect 15896 6196 15902 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18322 6236 18328 6248
rect 18279 6208 18328 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 26970 6196 26976 6248
rect 27028 6236 27034 6248
rect 37734 6236 37740 6248
rect 27028 6208 37740 6236
rect 27028 6196 27034 6208
rect 37734 6196 37740 6208
rect 37792 6196 37798 6248
rect 3605 6171 3663 6177
rect 3605 6137 3617 6171
rect 3651 6168 3663 6171
rect 11698 6168 11704 6180
rect 3651 6140 11704 6168
rect 3651 6137 3663 6140
rect 3605 6131 3663 6137
rect 11698 6128 11704 6140
rect 11756 6128 11762 6180
rect 28350 6128 28356 6180
rect 28408 6168 28414 6180
rect 39206 6168 39212 6180
rect 28408 6140 39212 6168
rect 28408 6128 28414 6140
rect 39206 6128 39212 6140
rect 39264 6128 39270 6180
rect 44177 6171 44235 6177
rect 44177 6137 44189 6171
rect 44223 6168 44235 6171
rect 47118 6168 47124 6180
rect 44223 6140 47124 6168
rect 44223 6137 44235 6140
rect 44177 6131 44235 6137
rect 47118 6128 47124 6140
rect 47176 6128 47182 6180
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 12434 6100 12440 6112
rect 2188 6072 12440 6100
rect 2188 6060 2194 6072
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19426 6100 19432 6112
rect 18739 6072 19432 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 37642 6060 37648 6112
rect 37700 6060 37706 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 47394 5896 47400 5908
rect 37700 5868 47400 5896
rect 37700 5856 37706 5868
rect 47394 5856 47400 5868
rect 47452 5856 47458 5908
rect 49145 5763 49203 5769
rect 49145 5729 49157 5763
rect 49191 5760 49203 5763
rect 49234 5760 49240 5772
rect 49191 5732 49240 5760
rect 49191 5729 49203 5732
rect 49145 5723 49203 5729
rect 49234 5720 49240 5732
rect 49292 5720 49298 5772
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1452 5664 1593 5692
rect 1452 5652 1458 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5692 2743 5695
rect 3329 5695 3387 5701
rect 2731 5664 2765 5692
rect 2731 5661 2743 5664
rect 2685 5655 2743 5661
rect 3329 5661 3341 5695
rect 3375 5692 3387 5695
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3375 5664 3985 5692
rect 3375 5661 3387 5664
rect 3329 5655 3387 5661
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 1302 5584 1308 5636
rect 1360 5624 1366 5636
rect 2700 5624 2728 5655
rect 43714 5652 43720 5704
rect 43772 5652 43778 5704
rect 47670 5652 47676 5704
rect 47728 5692 47734 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 47728 5664 47961 5692
rect 47728 5652 47734 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 3418 5624 3424 5636
rect 1360 5596 3424 5624
rect 1360 5584 1366 5596
rect 3418 5584 3424 5596
rect 3476 5584 3482 5636
rect 43901 5627 43959 5633
rect 43901 5593 43913 5627
rect 43947 5624 43959 5627
rect 45646 5624 45652 5636
rect 43947 5596 45652 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 45646 5584 45652 5596
rect 45704 5584 45710 5636
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5556 2283 5559
rect 2866 5556 2872 5568
rect 2271 5528 2872 5556
rect 2271 5525 2283 5528
rect 2225 5519 2283 5525
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 16022 5556 16028 5568
rect 4203 5528 16028 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 3418 5312 3424 5364
rect 3476 5312 3482 5364
rect 11882 5284 11888 5296
rect 2746 5256 11888 5284
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2746 5216 2774 5256
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 37274 5244 37280 5296
rect 37332 5284 37338 5296
rect 37369 5287 37427 5293
rect 37369 5284 37381 5287
rect 37332 5256 37381 5284
rect 37332 5244 37338 5256
rect 37369 5253 37381 5256
rect 37415 5284 37427 5287
rect 37737 5287 37795 5293
rect 37737 5284 37749 5287
rect 37415 5256 37749 5284
rect 37415 5253 37427 5256
rect 37369 5247 37427 5253
rect 37737 5253 37749 5256
rect 37783 5253 37795 5287
rect 37737 5247 37795 5253
rect 38470 5244 38476 5296
rect 38528 5284 38534 5296
rect 38933 5287 38991 5293
rect 38933 5284 38945 5287
rect 38528 5256 38945 5284
rect 38528 5244 38534 5256
rect 38933 5253 38945 5256
rect 38979 5253 38991 5287
rect 38933 5247 38991 5253
rect 49142 5244 49148 5296
rect 49200 5244 49206 5296
rect 2179 5188 2774 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 18874 5176 18880 5228
rect 18932 5176 18938 5228
rect 45738 5176 45744 5228
rect 45796 5216 45802 5228
rect 45833 5219 45891 5225
rect 45833 5216 45845 5219
rect 45796 5188 45845 5216
rect 45796 5176 45802 5188
rect 45833 5185 45845 5188
rect 45879 5185 45891 5219
rect 45833 5179 45891 5185
rect 47854 5176 47860 5228
rect 47912 5216 47918 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47912 5188 47961 5216
rect 47912 5176 47918 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 1360 5120 2421 5148
rect 1360 5108 1366 5120
rect 2409 5117 2421 5120
rect 2455 5148 2467 5151
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 2455 5120 3801 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 3789 5117 3801 5120
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 19058 5108 19064 5160
rect 19116 5108 19122 5160
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48314 5148 48320 5160
rect 46891 5120 48320 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 13354 5080 13360 5092
rect 3099 5052 13360 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 13354 5040 13360 5052
rect 13412 5040 13418 5092
rect 38657 5083 38715 5089
rect 38657 5049 38669 5083
rect 38703 5080 38715 5083
rect 40034 5080 40040 5092
rect 38703 5052 40040 5080
rect 38703 5049 38715 5052
rect 38657 5043 38715 5049
rect 40034 5040 40040 5052
rect 40092 5040 40098 5092
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 3605 5015 3663 5021
rect 3605 5012 3617 5015
rect 1452 4984 3617 5012
rect 1452 4972 1458 4984
rect 3605 4981 3617 4984
rect 3651 4981 3663 5015
rect 3605 4975 3663 4981
rect 19521 5015 19579 5021
rect 19521 4981 19533 5015
rect 19567 5012 19579 5015
rect 20622 5012 20628 5024
rect 19567 4984 20628 5012
rect 19567 4981 19579 4984
rect 19521 4975 19579 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 37826 4972 37832 5024
rect 37884 4972 37890 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 3510 4808 3516 4820
rect 2915 4780 3516 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 23382 4808 23388 4820
rect 5592 4780 23388 4808
rect 5592 4768 5598 4780
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 25774 4768 25780 4820
rect 25832 4808 25838 4820
rect 36446 4808 36452 4820
rect 25832 4780 36452 4808
rect 25832 4768 25838 4780
rect 36446 4768 36452 4780
rect 36504 4768 36510 4820
rect 36814 4768 36820 4820
rect 36872 4768 36878 4820
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 47302 4808 47308 4820
rect 37884 4780 47308 4808
rect 37884 4768 37890 4780
rect 47302 4768 47308 4780
rect 47360 4768 47366 4820
rect 19058 4700 19064 4752
rect 19116 4740 19122 4752
rect 22557 4743 22615 4749
rect 19116 4712 22094 4740
rect 19116 4700 19122 4712
rect 3237 4675 3295 4681
rect 3237 4672 3249 4675
rect 1596 4644 3249 4672
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1596 4613 1624 4644
rect 3237 4641 3249 4644
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 19242 4632 19248 4684
rect 19300 4672 19306 4684
rect 20441 4675 20499 4681
rect 20441 4672 20453 4675
rect 19300 4644 20453 4672
rect 19300 4632 19306 4644
rect 20441 4641 20453 4644
rect 20487 4641 20499 4675
rect 20441 4635 20499 4641
rect 21910 4632 21916 4684
rect 21968 4632 21974 4684
rect 22066 4672 22094 4712
rect 22557 4709 22569 4743
rect 22603 4740 22615 4743
rect 26142 4740 26148 4752
rect 22603 4712 26148 4740
rect 22603 4709 22615 4712
rect 22557 4703 22615 4709
rect 26142 4700 26148 4712
rect 26200 4700 26206 4752
rect 46474 4700 46480 4752
rect 46532 4700 46538 4752
rect 47210 4700 47216 4752
rect 47268 4700 47274 4752
rect 23566 4672 23572 4684
rect 22066 4644 23572 4672
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 2682 4564 2688 4616
rect 2740 4564 2746 4616
rect 19978 4564 19984 4616
rect 20036 4604 20042 4616
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 20036 4576 20637 4604
rect 20036 4564 20042 4576
rect 20625 4573 20637 4576
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 23124 4613 23152 4644
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 49145 4675 49203 4681
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49418 4672 49424 4684
rect 49191 4644 49424 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 23084 4607 23152 4613
rect 23084 4573 23096 4607
rect 23130 4576 23152 4607
rect 23130 4573 23142 4576
rect 23084 4567 23142 4573
rect 23198 4564 23204 4616
rect 23256 4604 23262 4616
rect 23256 4576 26004 4604
rect 23256 4564 23262 4576
rect 2225 4539 2283 4545
rect 2225 4505 2237 4539
rect 2271 4536 2283 4539
rect 4065 4539 4123 4545
rect 4065 4536 4077 4539
rect 2271 4508 4077 4536
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 4065 4505 4077 4508
rect 4111 4505 4123 4539
rect 4065 4499 4123 4505
rect 15838 4496 15844 4548
rect 15896 4536 15902 4548
rect 25869 4539 25927 4545
rect 25869 4536 25881 4539
rect 15896 4508 25881 4536
rect 15896 4496 15902 4508
rect 25869 4505 25881 4508
rect 25915 4505 25927 4539
rect 25976 4536 26004 4576
rect 36814 4564 36820 4616
rect 36872 4604 36878 4616
rect 37277 4607 37335 4613
rect 37277 4604 37289 4607
rect 36872 4576 37289 4604
rect 36872 4564 36878 4576
rect 37277 4573 37289 4576
rect 37323 4573 37335 4607
rect 37277 4567 37335 4573
rect 37734 4564 37740 4616
rect 37792 4604 37798 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 37792 4576 38025 4604
rect 37792 4564 37798 4576
rect 38013 4573 38025 4576
rect 38059 4604 38071 4607
rect 38473 4607 38531 4613
rect 38473 4604 38485 4607
rect 38059 4576 38485 4604
rect 38059 4573 38071 4576
rect 38013 4567 38071 4573
rect 38473 4573 38485 4576
rect 38519 4573 38531 4607
rect 38473 4567 38531 4573
rect 46934 4564 46940 4616
rect 46992 4604 46998 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 46992 4576 47961 4604
rect 46992 4564 46998 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 26789 4539 26847 4545
rect 26789 4536 26801 4539
rect 25976 4508 26801 4536
rect 25869 4499 25927 4505
rect 26789 4505 26801 4508
rect 26835 4505 26847 4539
rect 26789 4499 26847 4505
rect 26881 4539 26939 4545
rect 26881 4505 26893 4539
rect 26927 4536 26939 4539
rect 28718 4536 28724 4548
rect 26927 4508 28724 4536
rect 26927 4505 26939 4508
rect 26881 4499 26939 4505
rect 28718 4496 28724 4508
rect 28776 4496 28782 4548
rect 38197 4539 38255 4545
rect 38197 4505 38209 4539
rect 38243 4536 38255 4539
rect 39758 4536 39764 4548
rect 38243 4508 39764 4536
rect 38243 4505 38255 4508
rect 38197 4499 38255 4505
rect 39758 4496 39764 4508
rect 39816 4496 39822 4548
rect 46661 4539 46719 4545
rect 46661 4505 46673 4539
rect 46707 4505 46719 4539
rect 46661 4499 46719 4505
rect 47397 4539 47455 4545
rect 47397 4505 47409 4539
rect 47443 4536 47455 4539
rect 47670 4536 47676 4548
rect 47443 4508 47676 4536
rect 47443 4505 47455 4508
rect 47397 4499 47455 4505
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 10962 4468 10968 4480
rect 4203 4440 10968 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21266 4468 21272 4480
rect 21131 4440 21272 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 23155 4471 23213 4477
rect 23155 4437 23167 4471
rect 23201 4468 23213 4471
rect 24762 4468 24768 4480
rect 23201 4440 24768 4468
rect 23201 4437 23213 4440
rect 23155 4431 23213 4437
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 37366 4428 37372 4480
rect 37424 4428 37430 4480
rect 46201 4471 46259 4477
rect 46201 4437 46213 4471
rect 46247 4468 46259 4471
rect 46676 4468 46704 4499
rect 47670 4496 47676 4508
rect 47728 4496 47734 4548
rect 49786 4468 49792 4480
rect 46247 4440 49792 4468
rect 46247 4437 46259 4440
rect 46201 4431 46259 4437
rect 49786 4428 49792 4440
rect 49844 4428 49850 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 2682 4264 2688 4276
rect 2271 4236 2688 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 2682 4224 2688 4236
rect 2740 4224 2746 4276
rect 37366 4224 37372 4276
rect 37424 4264 37430 4276
rect 45830 4264 45836 4276
rect 37424 4236 45836 4264
rect 37424 4224 37430 4236
rect 45830 4224 45836 4236
rect 45888 4224 45894 4276
rect 17037 4199 17095 4205
rect 3252 4168 3464 4196
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1268 4100 1593 4128
rect 1268 4088 1274 4100
rect 1581 4097 1593 4100
rect 1627 4128 1639 4131
rect 3252 4128 3280 4168
rect 1627 4100 3280 4128
rect 3329 4131 3387 4137
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3436 4128 3464 4168
rect 17037 4165 17049 4199
rect 17083 4196 17095 4199
rect 18322 4196 18328 4208
rect 17083 4168 18328 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 18322 4156 18328 4168
rect 18380 4196 18386 4208
rect 18380 4168 19104 4196
rect 18380 4156 18386 4168
rect 3789 4131 3847 4137
rect 3789 4128 3801 4131
rect 3436 4100 3801 4128
rect 3329 4091 3387 4097
rect 3789 4097 3801 4100
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 3344 4060 3372 4091
rect 15746 4088 15752 4140
rect 15804 4088 15810 4140
rect 19076 4128 19104 4168
rect 22094 4156 22100 4208
rect 22152 4196 22158 4208
rect 22152 4168 23336 4196
rect 22152 4156 22158 4168
rect 22348 4131 22406 4137
rect 22348 4128 22360 4131
rect 19076 4100 22360 4128
rect 22348 4097 22360 4100
rect 22394 4128 22406 4131
rect 22960 4131 23018 4137
rect 22960 4128 22972 4131
rect 22394 4100 22876 4128
rect 22394 4097 22406 4100
rect 22348 4091 22406 4097
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 1360 4032 3617 4060
rect 1360 4020 1366 4032
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 14550 4020 14556 4072
rect 14608 4020 14614 4072
rect 1118 3952 1124 4004
rect 1176 3992 1182 4004
rect 14568 3992 14596 4020
rect 1176 3964 14596 3992
rect 22848 3992 22876 4100
rect 22940 4097 22972 4128
rect 23006 4097 23018 4131
rect 22940 4091 23018 4097
rect 23063 4131 23121 4137
rect 23063 4097 23075 4131
rect 23109 4128 23121 4131
rect 23198 4128 23204 4140
rect 23109 4100 23204 4128
rect 23109 4097 23121 4100
rect 23063 4091 23121 4097
rect 22940 4060 22968 4091
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23308 4128 23336 4168
rect 24762 4156 24768 4208
rect 24820 4196 24826 4208
rect 25869 4199 25927 4205
rect 25869 4196 25881 4199
rect 24820 4168 25881 4196
rect 24820 4156 24826 4168
rect 25869 4165 25881 4168
rect 25915 4165 25927 4199
rect 28813 4199 28871 4205
rect 28813 4196 28825 4199
rect 25869 4159 25927 4165
rect 28092 4168 28825 4196
rect 23604 4131 23662 4137
rect 23604 4128 23616 4131
rect 23308 4100 23616 4128
rect 23604 4097 23616 4100
rect 23650 4097 23662 4131
rect 23604 4091 23662 4097
rect 23290 4060 23296 4072
rect 22940 4032 23296 4060
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 24854 4020 24860 4072
rect 24912 4060 24918 4072
rect 24949 4063 25007 4069
rect 24949 4060 24961 4063
rect 24912 4032 24961 4060
rect 24912 4020 24918 4032
rect 24949 4029 24961 4032
rect 24995 4029 25007 4063
rect 24949 4023 25007 4029
rect 25961 4063 26019 4069
rect 25961 4029 25973 4063
rect 26007 4060 26019 4063
rect 27798 4060 27804 4072
rect 26007 4032 27804 4060
rect 26007 4029 26019 4032
rect 25961 4023 26019 4029
rect 27798 4020 27804 4032
rect 27856 4020 27862 4072
rect 27890 4020 27896 4072
rect 27948 4020 27954 4072
rect 23707 3995 23765 4001
rect 22848 3964 22968 3992
rect 1176 3952 1182 3964
rect 2682 3884 2688 3936
rect 2740 3884 2746 3936
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 13412 3896 16957 3924
rect 13412 3884 13418 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 16945 3887 17003 3893
rect 22419 3927 22477 3933
rect 22419 3893 22431 3927
rect 22465 3924 22477 3927
rect 22830 3924 22836 3936
rect 22465 3896 22836 3924
rect 22465 3893 22477 3896
rect 22419 3887 22477 3893
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 22940 3924 22968 3964
rect 23707 3961 23719 3995
rect 23753 3992 23765 3995
rect 28092 3992 28120 4168
rect 28813 4165 28825 4168
rect 28859 4165 28871 4199
rect 28813 4159 28871 4165
rect 36538 4088 36544 4140
rect 36596 4128 36602 4140
rect 45833 4131 45891 4137
rect 45833 4128 45845 4131
rect 36596 4100 45845 4128
rect 36596 4088 36602 4100
rect 45833 4097 45845 4100
rect 45879 4097 45891 4131
rect 45833 4091 45891 4097
rect 47026 4088 47032 4140
rect 47084 4128 47090 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 47084 4100 47961 4128
rect 47084 4088 47090 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4128 49203 4131
rect 49326 4128 49332 4140
rect 49191 4100 49332 4128
rect 49191 4097 49203 4100
rect 49145 4091 49203 4097
rect 49326 4088 49332 4100
rect 49384 4088 49390 4140
rect 28905 4063 28963 4069
rect 28905 4029 28917 4063
rect 28951 4060 28963 4063
rect 35066 4060 35072 4072
rect 28951 4032 35072 4060
rect 28951 4029 28963 4032
rect 28905 4023 28963 4029
rect 35066 4020 35072 4032
rect 35124 4020 35130 4072
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 23753 3964 28120 3992
rect 23753 3961 23765 3964
rect 23707 3955 23765 3961
rect 27522 3924 27528 3936
rect 22940 3896 27528 3924
rect 27522 3884 27528 3896
rect 27580 3884 27586 3936
rect 47670 3884 47676 3936
rect 47728 3884 47734 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7524 3692 12434 3720
rect 7524 3680 7530 3692
rect 3145 3655 3203 3661
rect 3145 3621 3157 3655
rect 3191 3652 3203 3655
rect 5534 3652 5540 3664
rect 3191 3624 5540 3652
rect 3191 3621 3203 3624
rect 3145 3615 3203 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 12406 3652 12434 3692
rect 19978 3680 19984 3732
rect 20036 3720 20042 3732
rect 23290 3720 23296 3732
rect 20036 3692 23296 3720
rect 20036 3680 20042 3692
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 23566 3680 23572 3732
rect 23624 3680 23630 3732
rect 23937 3723 23995 3729
rect 23937 3689 23949 3723
rect 23983 3720 23995 3723
rect 25958 3720 25964 3732
rect 23983 3692 25964 3720
rect 23983 3689 23995 3692
rect 23937 3683 23995 3689
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 36538 3680 36544 3732
rect 36596 3680 36602 3732
rect 17678 3652 17684 3664
rect 12406 3624 17684 3652
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 1360 3556 2421 3584
rect 1360 3544 1366 3556
rect 2409 3553 2421 3556
rect 2455 3584 2467 3587
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 2455 3556 3433 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 15286 3584 15292 3596
rect 5408 3556 15292 3584
rect 5408 3544 5414 3556
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 16592 3593 16620 3624
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 16577 3587 16635 3593
rect 16577 3553 16589 3587
rect 16623 3553 16635 3587
rect 25317 3587 25375 3593
rect 25317 3584 25329 3587
rect 16577 3547 16635 3553
rect 17604 3556 25329 3584
rect 2130 3476 2136 3528
rect 2188 3476 2194 3528
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 2961 3519 3019 3525
rect 2961 3516 2973 3519
rect 2740 3488 2973 3516
rect 2740 3476 2746 3488
rect 2961 3485 2973 3488
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 10318 3516 10324 3528
rect 9723 3488 10324 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 11149 3519 11207 3525
rect 11149 3516 11161 3519
rect 10468 3488 11161 3516
rect 10468 3476 10474 3488
rect 11149 3485 11161 3488
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 12345 3519 12403 3525
rect 12345 3516 12357 3519
rect 11839 3488 12357 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 12345 3485 12357 3488
rect 12391 3485 12403 3519
rect 12345 3479 12403 3485
rect 15749 3519 15807 3525
rect 15749 3485 15761 3519
rect 15795 3516 15807 3519
rect 15838 3516 15844 3528
rect 15795 3488 15844 3516
rect 15795 3485 15807 3488
rect 15749 3479 15807 3485
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 17604 3525 17632 3556
rect 25317 3553 25329 3556
rect 25363 3553 25375 3587
rect 28350 3584 28356 3596
rect 25317 3547 25375 3553
rect 25516 3556 28356 3584
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 20990 3476 20996 3528
rect 21048 3476 21054 3528
rect 22830 3476 22836 3528
rect 22888 3516 22894 3528
rect 22888 3488 23704 3516
rect 22888 3476 22894 3488
rect 3326 3408 3332 3460
rect 3384 3448 3390 3460
rect 14737 3451 14795 3457
rect 14737 3448 14749 3451
rect 3384 3420 14749 3448
rect 3384 3408 3390 3420
rect 14737 3417 14749 3420
rect 14783 3448 14795 3451
rect 18966 3448 18972 3460
rect 14783 3420 18972 3448
rect 14783 3417 14795 3420
rect 14737 3411 14795 3417
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 21269 3451 21327 3457
rect 21269 3448 21281 3451
rect 19392 3420 21281 3448
rect 19392 3408 19398 3420
rect 21269 3417 21281 3420
rect 21315 3417 21327 3451
rect 23676 3448 23704 3488
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 24029 3519 24087 3525
rect 24029 3516 24041 3519
rect 23808 3488 24041 3516
rect 23808 3476 23814 3488
rect 24029 3485 24041 3488
rect 24075 3516 24087 3519
rect 25516 3516 25544 3556
rect 28350 3544 28356 3556
rect 28408 3544 28414 3596
rect 33962 3544 33968 3596
rect 34020 3584 34026 3596
rect 45373 3587 45431 3593
rect 45373 3584 45385 3587
rect 34020 3556 45385 3584
rect 34020 3544 34026 3556
rect 45373 3553 45385 3556
rect 45419 3553 45431 3587
rect 45373 3547 45431 3553
rect 49142 3544 49148 3596
rect 49200 3544 49206 3596
rect 24075 3488 25544 3516
rect 24075 3485 24087 3488
rect 24029 3479 24087 3485
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 31754 3516 31760 3528
rect 26568 3488 31760 3516
rect 26568 3476 26574 3488
rect 31754 3476 31760 3488
rect 31812 3476 31818 3528
rect 36446 3476 36452 3528
rect 36504 3516 36510 3528
rect 36909 3519 36967 3525
rect 36909 3516 36921 3519
rect 36504 3488 36921 3516
rect 36504 3476 36510 3488
rect 36909 3485 36921 3488
rect 36955 3485 36967 3519
rect 36909 3479 36967 3485
rect 40034 3476 40040 3528
rect 40092 3516 40098 3528
rect 46109 3519 46167 3525
rect 46109 3516 46121 3519
rect 40092 3488 46121 3516
rect 40092 3476 40098 3488
rect 46109 3485 46121 3488
rect 46155 3485 46167 3519
rect 46109 3479 46167 3485
rect 47118 3476 47124 3528
rect 47176 3516 47182 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 47176 3488 47961 3516
rect 47176 3476 47182 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 26237 3451 26295 3457
rect 26237 3448 26249 3451
rect 22494 3420 23152 3448
rect 23676 3420 26249 3448
rect 21269 3411 21327 3417
rect 3786 3340 3792 3392
rect 3844 3340 3850 3392
rect 10321 3383 10379 3389
rect 10321 3349 10333 3383
rect 10367 3380 10379 3383
rect 10686 3380 10692 3392
rect 10367 3352 10692 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 12989 3383 13047 3389
rect 12989 3349 13001 3383
rect 13035 3380 13047 3383
rect 14826 3380 14832 3392
rect 13035 3352 14832 3380
rect 13035 3349 13047 3352
rect 12989 3343 13047 3349
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 21284 3380 21312 3411
rect 22278 3380 22284 3392
rect 21284 3352 22284 3380
rect 22278 3340 22284 3352
rect 22336 3340 22342 3392
rect 22738 3340 22744 3392
rect 22796 3340 22802 3392
rect 23124 3389 23152 3420
rect 26237 3417 26249 3420
rect 26283 3417 26295 3451
rect 26237 3411 26295 3417
rect 26329 3451 26387 3457
rect 26329 3417 26341 3451
rect 26375 3448 26387 3451
rect 28994 3448 29000 3460
rect 26375 3420 29000 3448
rect 26375 3417 26387 3420
rect 26329 3411 26387 3417
rect 28994 3408 29000 3420
rect 29052 3408 29058 3460
rect 31294 3448 31300 3460
rect 29104 3420 31300 3448
rect 23109 3383 23167 3389
rect 23109 3349 23121 3383
rect 23155 3380 23167 3383
rect 26510 3380 26516 3392
rect 23155 3352 26516 3380
rect 23155 3349 23167 3352
rect 23109 3343 23167 3349
rect 26510 3340 26516 3352
rect 26568 3340 26574 3392
rect 28350 3340 28356 3392
rect 28408 3380 28414 3392
rect 29104 3380 29132 3420
rect 31294 3408 31300 3420
rect 31352 3408 31358 3460
rect 45097 3451 45155 3457
rect 45097 3417 45109 3451
rect 45143 3448 45155 3451
rect 45554 3448 45560 3460
rect 45143 3420 45560 3448
rect 45143 3417 45155 3420
rect 45097 3411 45155 3417
rect 45554 3408 45560 3420
rect 45612 3448 45618 3460
rect 47305 3451 47363 3457
rect 45612 3420 45657 3448
rect 45612 3408 45618 3420
rect 47305 3417 47317 3451
rect 47351 3448 47363 3451
rect 48682 3448 48688 3460
rect 47351 3420 48688 3448
rect 47351 3417 47363 3420
rect 47305 3411 47363 3417
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 28408 3352 29132 3380
rect 28408 3340 28414 3352
rect 29546 3340 29552 3392
rect 29604 3340 29610 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 3605 3179 3663 3185
rect 3605 3145 3617 3179
rect 3651 3176 3663 3179
rect 4062 3176 4068 3188
rect 3651 3148 4068 3176
rect 3651 3145 3663 3148
rect 3605 3139 3663 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 15194 3176 15200 3188
rect 14568 3148 15200 3176
rect 4157 3111 4215 3117
rect 4157 3108 4169 3111
rect 1596 3080 4169 3108
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1596 3049 1624 3080
rect 4157 3077 4169 3080
rect 4203 3077 4215 3111
rect 4157 3071 4215 3077
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 3436 2972 3464 3003
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9640 3012 9689 3040
rect 9640 3000 9646 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13354 3040 13360 3052
rect 13219 3012 13360 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 14568 3049 14596 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 19334 3176 19340 3188
rect 16347 3148 19340 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19981 3179 20039 3185
rect 19981 3176 19993 3179
rect 19536 3148 19993 3176
rect 14826 3068 14832 3120
rect 14884 3068 14890 3120
rect 16574 3108 16580 3120
rect 16054 3080 16580 3108
rect 16574 3068 16580 3080
rect 16632 3108 16638 3120
rect 16669 3111 16727 3117
rect 16669 3108 16681 3111
rect 16632 3080 16681 3108
rect 16632 3068 16638 3080
rect 16669 3077 16681 3080
rect 16715 3077 16727 3111
rect 16669 3071 16727 3077
rect 17497 3111 17555 3117
rect 17497 3077 17509 3111
rect 17543 3108 17555 3111
rect 19058 3108 19064 3120
rect 17543 3080 19064 3108
rect 17543 3077 17555 3080
rect 17497 3071 17555 3077
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19536 3049 19564 3148
rect 19981 3145 19993 3148
rect 20027 3145 20039 3179
rect 19981 3139 20039 3145
rect 21453 3179 21511 3185
rect 21453 3145 21465 3179
rect 21499 3176 21511 3179
rect 24578 3176 24584 3188
rect 21499 3148 24584 3176
rect 21499 3145 21511 3148
rect 21453 3139 21511 3145
rect 24578 3136 24584 3148
rect 24636 3136 24642 3188
rect 25958 3136 25964 3188
rect 26016 3136 26022 3188
rect 27522 3136 27528 3188
rect 27580 3136 27586 3188
rect 27798 3136 27804 3188
rect 27856 3176 27862 3188
rect 31205 3179 31263 3185
rect 31205 3176 31217 3179
rect 27856 3148 31217 3176
rect 27856 3136 27862 3148
rect 31205 3145 31217 3148
rect 31251 3145 31263 3179
rect 31205 3139 31263 3145
rect 31294 3136 31300 3188
rect 31352 3176 31358 3188
rect 31352 3148 38056 3176
rect 31352 3136 31358 3148
rect 25976 3108 26004 3136
rect 29181 3111 29239 3117
rect 29181 3108 29193 3111
rect 25976 3080 29193 3108
rect 29181 3077 29193 3080
rect 29227 3077 29239 3111
rect 31754 3108 31760 3120
rect 30406 3080 31760 3108
rect 29181 3071 29239 3077
rect 31754 3068 31760 3080
rect 31812 3108 31818 3120
rect 31812 3080 31857 3108
rect 31812 3068 31818 3080
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 2271 2944 3464 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11756 2944 11989 2972
rect 11756 2932 11762 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 14516 2944 17325 2972
rect 14516 2932 14522 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 2961 2907 3019 2913
rect 2961 2873 2973 2907
rect 3007 2904 3019 2907
rect 3602 2904 3608 2916
rect 3007 2876 3608 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 3602 2864 3608 2876
rect 3660 2864 3666 2916
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 3973 2839 4031 2845
rect 3973 2836 3985 2839
rect 3936 2808 3985 2836
rect 3936 2796 3942 2808
rect 3973 2805 3985 2808
rect 4019 2805 4031 2839
rect 3973 2799 4031 2805
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 9582 2836 9588 2848
rect 9447 2808 9588 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 20180 2836 20208 3003
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 21266 3000 21272 3052
rect 21324 3000 21330 3052
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3040 22707 3043
rect 23750 3040 23756 3052
rect 22695 3012 23756 3040
rect 22695 3009 22707 3012
rect 22649 3003 22707 3009
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 21048 2944 24225 2972
rect 21048 2932 21054 2944
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24489 2975 24547 2981
rect 24489 2972 24501 2975
rect 24213 2935 24271 2941
rect 24320 2944 24501 2972
rect 20809 2907 20867 2913
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 22094 2904 22100 2916
rect 20855 2876 22100 2904
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 22186 2864 22192 2916
rect 22244 2864 22250 2916
rect 22738 2864 22744 2916
rect 22796 2904 22802 2916
rect 24320 2904 24348 2944
rect 24489 2941 24501 2944
rect 24535 2941 24547 2975
rect 25608 2972 25636 3026
rect 26142 3000 26148 3052
rect 26200 3040 26206 3052
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 26200 3012 26433 3040
rect 26200 3000 26206 3012
rect 26421 3009 26433 3012
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 27985 3043 28043 3049
rect 27985 3009 27997 3043
rect 28031 3040 28043 3043
rect 28350 3040 28356 3052
rect 28031 3012 28356 3040
rect 28031 3009 28043 3012
rect 27985 3003 28043 3009
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28868 3012 28917 3040
rect 28868 3000 28874 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 31386 3000 31392 3052
rect 31444 3000 31450 3052
rect 33137 3043 33195 3049
rect 33137 3009 33149 3043
rect 33183 3040 33195 3043
rect 33686 3040 33692 3052
rect 33183 3012 33692 3040
rect 33183 3009 33195 3012
rect 33137 3003 33195 3009
rect 33686 3000 33692 3012
rect 33744 3000 33750 3052
rect 35250 3000 35256 3052
rect 35308 3000 35314 3052
rect 38028 3049 38056 3148
rect 49145 3111 49203 3117
rect 49145 3077 49157 3111
rect 49191 3108 49203 3111
rect 49234 3108 49240 3120
rect 49191 3080 49240 3108
rect 49191 3077 49203 3080
rect 49145 3071 49203 3077
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 38013 3043 38071 3049
rect 38013 3009 38025 3043
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 39816 3012 44005 3040
rect 39816 3000 39822 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 45646 3000 45652 3052
rect 45704 3040 45710 3052
rect 45833 3043 45891 3049
rect 45833 3040 45845 3043
rect 45704 3012 45845 3040
rect 45704 3000 45710 3012
rect 45833 3009 45845 3012
rect 45879 3009 45891 3043
rect 45833 3003 45891 3009
rect 47394 3000 47400 3052
rect 47452 3040 47458 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47452 3012 47961 3040
rect 47452 3000 47458 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 26326 2972 26332 2984
rect 25608 2944 26332 2972
rect 24489 2935 24547 2941
rect 26326 2932 26332 2944
rect 26384 2972 26390 2984
rect 26510 2972 26516 2984
rect 26384 2944 26516 2972
rect 26384 2932 26390 2944
rect 26510 2932 26516 2944
rect 26568 2932 26574 2984
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 28776 2944 31754 2972
rect 28776 2932 28782 2944
rect 31726 2904 31754 2944
rect 38286 2932 38292 2984
rect 38344 2932 38350 2984
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 46750 2972 46756 2984
rect 45235 2944 46756 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 46842 2932 46848 2984
rect 46900 2932 46906 2984
rect 32953 2907 33011 2913
rect 32953 2904 32965 2907
rect 22796 2876 24348 2904
rect 30668 2876 31340 2904
rect 31726 2876 32965 2904
rect 22796 2864 22802 2876
rect 22204 2836 22232 2864
rect 20180 2808 22232 2836
rect 22278 2796 22284 2848
rect 22336 2836 22342 2848
rect 22373 2839 22431 2845
rect 22373 2836 22385 2839
rect 22336 2808 22385 2836
rect 22336 2796 22342 2808
rect 22373 2805 22385 2808
rect 22419 2805 22431 2839
rect 22373 2799 22431 2805
rect 23290 2796 23296 2848
rect 23348 2796 23354 2848
rect 23492 2845 23520 2876
rect 23477 2839 23535 2845
rect 23477 2805 23489 2839
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 26605 2839 26663 2845
rect 26605 2805 26617 2839
rect 26651 2836 26663 2839
rect 27154 2836 27160 2848
rect 26651 2808 27160 2836
rect 26651 2805 26663 2808
rect 26605 2799 26663 2805
rect 27154 2796 27160 2808
rect 27212 2796 27218 2848
rect 30668 2845 30696 2876
rect 27893 2839 27951 2845
rect 27893 2805 27905 2839
rect 27939 2836 27951 2839
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 27939 2808 30665 2836
rect 27939 2805 27951 2808
rect 27893 2799 27951 2805
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 31312 2836 31340 2876
rect 32953 2873 32965 2876
rect 32999 2873 33011 2907
rect 40678 2904 40684 2916
rect 32953 2867 33011 2873
rect 34992 2876 40684 2904
rect 34992 2836 35020 2876
rect 40678 2864 40684 2876
rect 40736 2864 40742 2916
rect 31312 2808 35020 2836
rect 30653 2799 30711 2805
rect 35066 2796 35072 2848
rect 35124 2796 35130 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2225 2635 2283 2641
rect 2225 2601 2237 2635
rect 2271 2632 2283 2635
rect 2774 2632 2780 2644
rect 2271 2604 2780 2632
rect 2271 2601 2283 2604
rect 2225 2595 2283 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 10410 2632 10416 2644
rect 9631 2604 10416 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 26326 2592 26332 2644
rect 26384 2592 26390 2644
rect 28994 2592 29000 2644
rect 29052 2592 29058 2644
rect 31386 2592 31392 2644
rect 31444 2632 31450 2644
rect 31573 2635 31631 2641
rect 31573 2632 31585 2635
rect 31444 2604 31585 2632
rect 31444 2592 31450 2604
rect 31573 2601 31585 2604
rect 31619 2601 31631 2635
rect 31573 2595 31631 2601
rect 33686 2592 33692 2644
rect 33744 2592 33750 2644
rect 35250 2592 35256 2644
rect 35308 2632 35314 2644
rect 35805 2635 35863 2641
rect 35805 2632 35817 2635
rect 35308 2604 35817 2632
rect 35308 2592 35314 2604
rect 35805 2601 35817 2604
rect 35851 2601 35863 2635
rect 35805 2595 35863 2601
rect 38105 2635 38163 2641
rect 38105 2601 38117 2635
rect 38151 2632 38163 2635
rect 38286 2632 38292 2644
rect 38151 2604 38292 2632
rect 38151 2601 38163 2604
rect 38105 2595 38163 2601
rect 38286 2592 38292 2604
rect 38344 2592 38350 2644
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 12802 2564 12808 2576
rect 4203 2536 12808 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 12802 2524 12808 2536
rect 12860 2524 12866 2576
rect 24854 2564 24860 2576
rect 16546 2536 24860 2564
rect 3786 2496 3792 2508
rect 1596 2468 3792 2496
rect 1210 2388 1216 2440
rect 1268 2428 1274 2440
rect 1596 2437 1624 2468
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 13265 2499 13323 2505
rect 13265 2465 13277 2499
rect 13311 2496 13323 2499
rect 13814 2496 13820 2508
rect 13311 2468 13820 2496
rect 13311 2465 13323 2468
rect 13265 2459 13323 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 15286 2456 15292 2508
rect 15344 2456 15350 2508
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1268 2400 1593 2428
rect 1268 2388 1274 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2428 3387 2431
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3375 2400 3985 2428
rect 3375 2397 3387 2400
rect 3329 2391 3387 2397
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 2700 2360 2728 2391
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4120 2400 4721 2428
rect 4120 2388 4126 2400
rect 4709 2397 4721 2400
rect 4755 2428 4767 2431
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 4755 2400 5181 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5169 2397 5181 2400
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2428 9459 2431
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 9447 2400 10057 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 10686 2388 10692 2440
rect 10744 2388 10750 2440
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 14458 2428 14464 2440
rect 13771 2400 14464 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16546 2428 16574 2536
rect 24854 2524 24860 2536
rect 24912 2524 24918 2576
rect 34146 2524 34152 2576
rect 34204 2564 34210 2576
rect 34204 2536 43852 2564
rect 34204 2524 34210 2536
rect 19978 2496 19984 2508
rect 18892 2468 19984 2496
rect 18892 2437 18920 2468
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22336 2468 22845 2496
rect 22336 2456 22342 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 24394 2456 24400 2508
rect 24452 2496 24458 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24452 2468 25053 2496
rect 24452 2456 24458 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 28994 2456 29000 2508
rect 29052 2496 29058 2508
rect 29546 2496 29552 2508
rect 29052 2468 29552 2496
rect 29052 2456 29058 2468
rect 29546 2456 29552 2468
rect 29604 2496 29610 2508
rect 29604 2468 29776 2496
rect 29604 2456 29610 2468
rect 16347 2400 16574 2428
rect 18233 2431 18291 2437
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18877 2431 18935 2437
rect 18279 2400 18736 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 3878 2360 3884 2372
rect 1360 2332 3884 2360
rect 1360 2320 1366 2332
rect 3878 2320 3884 2332
rect 3936 2320 3942 2372
rect 12066 2360 12072 2372
rect 4908 2332 12072 2360
rect 4908 2301 4936 2332
rect 12066 2320 12072 2332
rect 12124 2320 12130 2372
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 17037 2363 17095 2369
rect 17037 2360 17049 2363
rect 15988 2332 17049 2360
rect 15988 2320 15994 2332
rect 17037 2329 17049 2332
rect 17083 2329 17095 2363
rect 17037 2323 17095 2329
rect 18708 2301 18736 2400
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 19628 2400 20085 2428
rect 19628 2301 19656 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22152 2400 22385 2428
rect 22152 2388 22158 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 29748 2437 29776 2468
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 43824 2505 43852 2536
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 41380 2468 41429 2496
rect 41380 2456 41386 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 41417 2459 41475 2465
rect 43809 2499 43867 2505
rect 43809 2465 43821 2499
rect 43855 2465 43867 2499
rect 43809 2459 43867 2465
rect 49142 2456 49148 2508
rect 49200 2456 49206 2508
rect 29181 2431 29239 2437
rect 29181 2397 29193 2431
rect 29227 2397 29239 2431
rect 29181 2391 29239 2397
rect 29733 2431 29791 2437
rect 29733 2397 29745 2431
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 29196 2360 29224 2391
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30800 2400 30941 2428
rect 30800 2388 30806 2400
rect 30929 2397 30941 2400
rect 30975 2428 30987 2431
rect 31849 2431 31907 2437
rect 31849 2428 31861 2431
rect 30975 2400 31861 2428
rect 30975 2397 30987 2400
rect 30929 2391 30987 2397
rect 31849 2397 31861 2400
rect 31895 2397 31907 2431
rect 33045 2431 33103 2437
rect 33045 2428 33057 2431
rect 31849 2391 31907 2397
rect 32876 2400 33057 2428
rect 30377 2363 30435 2369
rect 30377 2360 30389 2363
rect 29196 2332 30389 2360
rect 30377 2329 30389 2332
rect 30423 2329 30435 2363
rect 30377 2323 30435 2329
rect 32876 2304 32904 2400
rect 33045 2397 33057 2400
rect 33091 2397 33103 2431
rect 35161 2431 35219 2437
rect 35161 2428 35173 2431
rect 33045 2391 33103 2397
rect 34992 2400 35173 2428
rect 34992 2304 35020 2400
rect 35161 2397 35173 2400
rect 35207 2397 35219 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35161 2391 35219 2397
rect 37108 2400 37473 2428
rect 37108 2304 37136 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 40678 2388 40684 2440
rect 40736 2388 40742 2440
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 43456 2400 43545 2428
rect 43456 2304 43484 2400
rect 43533 2397 43545 2400
rect 43579 2397 43591 2431
rect 43533 2391 43591 2397
rect 45830 2388 45836 2440
rect 45888 2388 45894 2440
rect 47302 2388 47308 2440
rect 47360 2428 47366 2440
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 47360 2400 47961 2428
rect 47360 2388 47366 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2360 47087 2363
rect 48498 2360 48504 2372
rect 47075 2332 48504 2360
rect 47075 2329 47087 2332
rect 47029 2323 47087 2329
rect 48498 2320 48504 2332
rect 48556 2320 48562 2372
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2261 4951 2295
rect 4893 2255 4951 2261
rect 18693 2295 18751 2301
rect 18693 2261 18705 2295
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 32769 2295 32827 2301
rect 32769 2261 32781 2295
rect 32815 2292 32827 2295
rect 32858 2292 32864 2304
rect 32815 2264 32864 2292
rect 32815 2261 32827 2264
rect 32769 2255 32827 2261
rect 32858 2252 32864 2264
rect 32916 2252 32922 2304
rect 34885 2295 34943 2301
rect 34885 2261 34897 2295
rect 34931 2292 34943 2295
rect 34974 2292 34980 2304
rect 34931 2264 34980 2292
rect 34931 2261 34943 2264
rect 34885 2255 34943 2261
rect 34974 2252 34980 2264
rect 35032 2252 35038 2304
rect 37090 2252 37096 2304
rect 37148 2252 37154 2304
rect 43257 2295 43315 2301
rect 43257 2261 43269 2295
rect 43303 2292 43315 2295
rect 43438 2292 43444 2304
rect 43303 2264 43444 2292
rect 43303 2261 43315 2264
rect 43257 2255 43315 2261
rect 43438 2252 43444 2264
rect 43496 2252 43502 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 34060 26324 34112 26376
rect 43352 26324 43404 26376
rect 4068 25168 4120 25220
rect 9772 25168 9824 25220
rect 21548 24828 21600 24880
rect 25964 24828 26016 24880
rect 16028 24760 16080 24812
rect 24492 24760 24544 24812
rect 18880 24692 18932 24744
rect 26332 24760 26384 24812
rect 26424 24760 26476 24812
rect 35164 24760 35216 24812
rect 29552 24692 29604 24744
rect 32864 24692 32916 24744
rect 34980 24692 35032 24744
rect 40592 24760 40644 24812
rect 35532 24692 35584 24744
rect 24768 24624 24820 24676
rect 30380 24624 30432 24676
rect 30564 24624 30616 24676
rect 38844 24624 38896 24676
rect 39212 24692 39264 24744
rect 43904 24692 43956 24744
rect 39396 24624 39448 24676
rect 39580 24624 39632 24676
rect 44364 24624 44416 24676
rect 45560 24624 45612 24676
rect 46756 24624 46808 24676
rect 3608 24556 3660 24608
rect 6552 24556 6604 24608
rect 20812 24556 20864 24608
rect 29736 24556 29788 24608
rect 31852 24556 31904 24608
rect 39488 24556 39540 24608
rect 40408 24556 40460 24608
rect 47124 24556 47176 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 19064 24352 19116 24404
rect 3516 24216 3568 24268
rect 3884 24148 3936 24200
rect 9864 24284 9916 24336
rect 6736 24216 6788 24268
rect 8668 24216 8720 24268
rect 11888 24284 11940 24336
rect 2320 24080 2372 24132
rect 7104 24148 7156 24200
rect 7472 24148 7524 24200
rect 12348 24216 12400 24268
rect 13820 24216 13872 24268
rect 17684 24216 17736 24268
rect 19616 24284 19668 24336
rect 20260 24284 20312 24336
rect 9588 24080 9640 24132
rect 13636 24148 13688 24200
rect 13728 24191 13780 24200
rect 13728 24157 13737 24191
rect 13737 24157 13771 24191
rect 13771 24157 13780 24191
rect 13728 24148 13780 24157
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 20628 24216 20680 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 24492 24284 24544 24336
rect 26424 24395 26476 24404
rect 26424 24361 26433 24395
rect 26433 24361 26467 24395
rect 26467 24361 26476 24395
rect 26424 24352 26476 24361
rect 29736 24395 29788 24404
rect 29736 24361 29745 24395
rect 29745 24361 29779 24395
rect 29779 24361 29788 24395
rect 29736 24352 29788 24361
rect 30196 24352 30248 24404
rect 35900 24352 35952 24404
rect 37556 24352 37608 24404
rect 39396 24352 39448 24404
rect 25780 24327 25832 24336
rect 25780 24293 25789 24327
rect 25789 24293 25823 24327
rect 25823 24293 25832 24327
rect 25780 24284 25832 24293
rect 26332 24284 26384 24336
rect 28632 24284 28684 24336
rect 26608 24259 26660 24268
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 20812 24148 20864 24200
rect 15568 24080 15620 24132
rect 17224 24080 17276 24132
rect 21456 24148 21508 24200
rect 25412 24148 25464 24200
rect 6644 24012 6696 24064
rect 7472 24012 7524 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 11152 24012 11204 24064
rect 11796 24012 11848 24064
rect 18604 24012 18656 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 22652 24080 22704 24132
rect 25320 24080 25372 24132
rect 23940 24012 23992 24064
rect 24860 24012 24912 24064
rect 26608 24225 26617 24259
rect 26617 24225 26651 24259
rect 26651 24225 26660 24259
rect 26608 24216 26660 24225
rect 27344 24216 27396 24268
rect 26056 24148 26108 24200
rect 26424 24080 26476 24132
rect 27252 24080 27304 24132
rect 27344 24123 27396 24132
rect 27344 24089 27353 24123
rect 27353 24089 27387 24123
rect 27387 24089 27396 24123
rect 27344 24080 27396 24089
rect 30380 24191 30432 24200
rect 30380 24157 30389 24191
rect 30389 24157 30423 24191
rect 30423 24157 30432 24191
rect 30380 24148 30432 24157
rect 30564 24284 30616 24336
rect 31300 24284 31352 24336
rect 33048 24284 33100 24336
rect 36452 24284 36504 24336
rect 31576 24216 31628 24268
rect 32772 24216 32824 24268
rect 34336 24216 34388 24268
rect 34980 24259 35032 24268
rect 34980 24225 34989 24259
rect 34989 24225 35023 24259
rect 35023 24225 35032 24259
rect 34980 24216 35032 24225
rect 35164 24259 35216 24268
rect 35164 24225 35173 24259
rect 35173 24225 35207 24259
rect 35207 24225 35216 24259
rect 35164 24216 35216 24225
rect 36728 24259 36780 24268
rect 36728 24225 36737 24259
rect 36737 24225 36771 24259
rect 36771 24225 36780 24259
rect 36728 24216 36780 24225
rect 37464 24216 37516 24268
rect 38660 24284 38712 24336
rect 32864 24148 32916 24200
rect 33324 24148 33376 24200
rect 33876 24148 33928 24200
rect 26976 24012 27028 24064
rect 27804 24012 27856 24064
rect 28356 24012 28408 24064
rect 28632 24012 28684 24064
rect 30564 24055 30616 24064
rect 30564 24021 30573 24055
rect 30573 24021 30607 24055
rect 30607 24021 30616 24055
rect 30564 24012 30616 24021
rect 31116 24012 31168 24064
rect 32312 24055 32364 24064
rect 32312 24021 32321 24055
rect 32321 24021 32355 24055
rect 32355 24021 32364 24055
rect 32312 24012 32364 24021
rect 34428 24080 34480 24132
rect 40132 24216 40184 24268
rect 40592 24259 40644 24268
rect 40592 24225 40601 24259
rect 40601 24225 40635 24259
rect 40635 24225 40644 24259
rect 40592 24216 40644 24225
rect 38844 24191 38896 24200
rect 38844 24157 38853 24191
rect 38853 24157 38887 24191
rect 38887 24157 38896 24191
rect 38844 24148 38896 24157
rect 39488 24191 39540 24200
rect 39488 24157 39497 24191
rect 39497 24157 39531 24191
rect 39531 24157 39540 24191
rect 39488 24148 39540 24157
rect 40408 24191 40460 24200
rect 40408 24157 40417 24191
rect 40417 24157 40451 24191
rect 40451 24157 40460 24191
rect 40408 24148 40460 24157
rect 42892 24284 42944 24336
rect 42156 24216 42208 24268
rect 44272 24352 44324 24404
rect 46296 24352 46348 24404
rect 47860 24352 47912 24404
rect 43536 24284 43588 24336
rect 43352 24148 43404 24200
rect 43536 24148 43588 24200
rect 46756 24284 46808 24336
rect 44456 24148 44508 24200
rect 42156 24080 42208 24132
rect 44732 24080 44784 24132
rect 47676 24148 47728 24200
rect 34060 24055 34112 24064
rect 34060 24021 34069 24055
rect 34069 24021 34103 24055
rect 34103 24021 34112 24055
rect 34060 24012 34112 24021
rect 35256 24055 35308 24064
rect 35256 24021 35265 24055
rect 35265 24021 35299 24055
rect 35299 24021 35308 24055
rect 35256 24012 35308 24021
rect 35624 24055 35676 24064
rect 35624 24021 35633 24055
rect 35633 24021 35667 24055
rect 35667 24021 35676 24055
rect 35624 24012 35676 24021
rect 36084 24055 36136 24064
rect 36084 24021 36093 24055
rect 36093 24021 36127 24055
rect 36127 24021 36136 24055
rect 36084 24012 36136 24021
rect 36820 24012 36872 24064
rect 37832 24055 37884 24064
rect 37832 24021 37841 24055
rect 37841 24021 37875 24055
rect 37875 24021 37884 24055
rect 37832 24012 37884 24021
rect 38384 24012 38436 24064
rect 40040 24055 40092 24064
rect 40040 24021 40049 24055
rect 40049 24021 40083 24055
rect 40083 24021 40092 24055
rect 40040 24012 40092 24021
rect 40960 24012 41012 24064
rect 42616 24012 42668 24064
rect 42800 24012 42852 24064
rect 44180 24055 44232 24064
rect 44180 24021 44189 24055
rect 44189 24021 44223 24055
rect 44223 24021 44232 24055
rect 44180 24012 44232 24021
rect 44640 24055 44692 24064
rect 44640 24021 44649 24055
rect 44649 24021 44683 24055
rect 44683 24021 44692 24055
rect 44640 24012 44692 24021
rect 45376 24012 45428 24064
rect 48044 24055 48096 24064
rect 48044 24021 48053 24055
rect 48053 24021 48087 24055
rect 48087 24021 48096 24055
rect 48044 24012 48096 24021
rect 48780 24055 48832 24064
rect 48780 24021 48789 24055
rect 48789 24021 48823 24055
rect 48823 24021 48832 24055
rect 48780 24012 48832 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 2320 23851 2372 23860
rect 2320 23817 2329 23851
rect 2329 23817 2363 23851
rect 2363 23817 2372 23851
rect 2320 23808 2372 23817
rect 4068 23715 4120 23724
rect 4068 23681 4077 23715
rect 4077 23681 4111 23715
rect 4111 23681 4120 23715
rect 4068 23672 4120 23681
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 4712 23672 4764 23681
rect 4160 23604 4212 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 3976 23536 4028 23588
rect 5816 23536 5868 23588
rect 8576 23672 8628 23724
rect 11796 23740 11848 23792
rect 12164 23672 12216 23724
rect 14372 23740 14424 23792
rect 19616 23808 19668 23860
rect 21456 23851 21508 23860
rect 21456 23817 21465 23851
rect 21465 23817 21499 23851
rect 21499 23817 21508 23851
rect 21456 23808 21508 23817
rect 19248 23740 19300 23792
rect 20352 23740 20404 23792
rect 8392 23604 8444 23656
rect 9220 23604 9272 23656
rect 10600 23647 10652 23656
rect 10600 23613 10609 23647
rect 10609 23613 10643 23647
rect 10643 23613 10652 23647
rect 10600 23604 10652 23613
rect 10324 23536 10376 23588
rect 12624 23647 12676 23656
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 16396 23604 16448 23656
rect 18328 23604 18380 23656
rect 17224 23536 17276 23588
rect 2780 23468 2832 23520
rect 5724 23468 5776 23520
rect 6000 23468 6052 23520
rect 18788 23511 18840 23520
rect 18788 23477 18797 23511
rect 18797 23477 18831 23511
rect 18831 23477 18840 23511
rect 18788 23468 18840 23477
rect 23480 23740 23532 23792
rect 25872 23740 25924 23792
rect 27712 23740 27764 23792
rect 23572 23672 23624 23724
rect 24952 23672 25004 23724
rect 21732 23604 21784 23656
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 23756 23647 23808 23656
rect 23756 23613 23765 23647
rect 23765 23613 23799 23647
rect 23799 23613 23808 23647
rect 23756 23604 23808 23613
rect 22744 23536 22796 23588
rect 23664 23536 23716 23588
rect 24860 23604 24912 23656
rect 25596 23604 25648 23656
rect 26608 23647 26660 23656
rect 26608 23613 26617 23647
rect 26617 23613 26651 23647
rect 26651 23613 26660 23647
rect 26608 23604 26660 23613
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 28540 23672 28592 23724
rect 40040 23808 40092 23860
rect 31024 23740 31076 23792
rect 31392 23740 31444 23792
rect 32496 23740 32548 23792
rect 33048 23740 33100 23792
rect 35624 23740 35676 23792
rect 39212 23783 39264 23792
rect 39212 23749 39221 23783
rect 39221 23749 39255 23783
rect 39255 23749 39264 23783
rect 39212 23740 39264 23749
rect 41696 23808 41748 23860
rect 42524 23808 42576 23860
rect 28448 23604 28500 23656
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 32772 23672 32824 23724
rect 29184 23604 29236 23656
rect 31024 23604 31076 23656
rect 31760 23647 31812 23656
rect 31760 23613 31769 23647
rect 31769 23613 31803 23647
rect 31803 23613 31812 23647
rect 31760 23604 31812 23613
rect 20812 23468 20864 23520
rect 20996 23468 21048 23520
rect 23848 23468 23900 23520
rect 24860 23511 24912 23520
rect 24860 23477 24869 23511
rect 24869 23477 24903 23511
rect 24903 23477 24912 23511
rect 24860 23468 24912 23477
rect 29736 23536 29788 23588
rect 29828 23536 29880 23588
rect 27804 23468 27856 23520
rect 29276 23511 29328 23520
rect 29276 23477 29285 23511
rect 29285 23477 29319 23511
rect 29319 23477 29328 23511
rect 29276 23468 29328 23477
rect 30288 23468 30340 23520
rect 32312 23468 32364 23520
rect 34980 23604 35032 23656
rect 35900 23579 35952 23588
rect 35900 23545 35909 23579
rect 35909 23545 35943 23579
rect 35943 23545 35952 23579
rect 35900 23536 35952 23545
rect 36176 23604 36228 23656
rect 36452 23647 36504 23656
rect 36452 23613 36461 23647
rect 36461 23613 36495 23647
rect 36495 23613 36504 23647
rect 36452 23604 36504 23613
rect 36544 23604 36596 23656
rect 38844 23672 38896 23724
rect 47308 23808 47360 23860
rect 49148 23851 49200 23860
rect 49148 23817 49157 23851
rect 49157 23817 49191 23851
rect 49191 23817 49200 23851
rect 49148 23808 49200 23817
rect 49516 23851 49568 23860
rect 49516 23817 49525 23851
rect 49525 23817 49559 23851
rect 49559 23817 49568 23851
rect 49516 23808 49568 23817
rect 42984 23740 43036 23792
rect 44824 23715 44876 23724
rect 44824 23681 44833 23715
rect 44833 23681 44867 23715
rect 44867 23681 44876 23715
rect 44824 23672 44876 23681
rect 34520 23468 34572 23520
rect 35440 23468 35492 23520
rect 36544 23468 36596 23520
rect 39764 23604 39816 23656
rect 41052 23604 41104 23656
rect 39488 23536 39540 23588
rect 46388 23715 46440 23724
rect 46388 23681 46397 23715
rect 46397 23681 46431 23715
rect 46431 23681 46440 23715
rect 46388 23672 46440 23681
rect 46848 23672 46900 23724
rect 48228 23672 48280 23724
rect 38568 23511 38620 23520
rect 38568 23477 38577 23511
rect 38577 23477 38611 23511
rect 38611 23477 38620 23511
rect 38568 23468 38620 23477
rect 39396 23468 39448 23520
rect 41512 23536 41564 23588
rect 43536 23579 43588 23588
rect 43536 23545 43545 23579
rect 43545 23545 43579 23579
rect 43579 23545 43588 23579
rect 43536 23536 43588 23545
rect 43996 23579 44048 23588
rect 43996 23545 44005 23579
rect 44005 23545 44039 23579
rect 44039 23545 44048 23579
rect 43996 23536 44048 23545
rect 46020 23536 46072 23588
rect 42432 23468 42484 23520
rect 42892 23511 42944 23520
rect 42892 23477 42901 23511
rect 42901 23477 42935 23511
rect 42935 23477 42944 23511
rect 42892 23468 42944 23477
rect 43628 23468 43680 23520
rect 44732 23468 44784 23520
rect 48044 23468 48096 23520
rect 49332 23511 49384 23520
rect 49332 23477 49341 23511
rect 49341 23477 49375 23511
rect 49375 23477 49384 23511
rect 49332 23468 49384 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 4712 23307 4764 23316
rect 4712 23273 4721 23307
rect 4721 23273 4755 23307
rect 4755 23273 4764 23307
rect 4712 23264 4764 23273
rect 23664 23264 23716 23316
rect 23756 23264 23808 23316
rect 28540 23264 28592 23316
rect 29184 23307 29236 23316
rect 29184 23273 29193 23307
rect 29193 23273 29227 23307
rect 29227 23273 29236 23307
rect 29184 23264 29236 23273
rect 29736 23307 29788 23316
rect 29736 23273 29745 23307
rect 29745 23273 29779 23307
rect 29779 23273 29788 23307
rect 29736 23264 29788 23273
rect 29920 23264 29972 23316
rect 33324 23264 33376 23316
rect 35072 23264 35124 23316
rect 36636 23264 36688 23316
rect 5632 23196 5684 23248
rect 4436 23060 4488 23112
rect 1768 23035 1820 23044
rect 1768 23001 1777 23035
rect 1777 23001 1811 23035
rect 1811 23001 1820 23035
rect 1768 22992 1820 23001
rect 3608 22992 3660 23044
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 15844 23196 15896 23248
rect 19616 23239 19668 23248
rect 19616 23205 19625 23239
rect 19625 23205 19659 23239
rect 19659 23205 19668 23239
rect 19616 23196 19668 23205
rect 20352 23239 20404 23248
rect 20352 23205 20361 23239
rect 20361 23205 20395 23239
rect 20395 23205 20404 23239
rect 20352 23196 20404 23205
rect 22744 23196 22796 23248
rect 25412 23196 25464 23248
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 13360 23128 13412 23180
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 6644 23060 6696 23112
rect 9128 23060 9180 23112
rect 11888 23103 11940 23112
rect 11888 23069 11897 23103
rect 11897 23069 11931 23103
rect 11931 23069 11940 23103
rect 11888 23060 11940 23069
rect 13912 23060 13964 23112
rect 17592 23128 17644 23180
rect 18236 23128 18288 23180
rect 19064 23128 19116 23180
rect 19248 23128 19300 23180
rect 20812 23128 20864 23180
rect 21732 23128 21784 23180
rect 24860 23128 24912 23180
rect 26332 23128 26384 23180
rect 7840 22992 7892 23044
rect 4620 22924 4672 22976
rect 5448 22924 5500 22976
rect 14188 22967 14240 22976
rect 14188 22933 14197 22967
rect 14197 22933 14231 22967
rect 14231 22933 14240 22967
rect 14188 22924 14240 22933
rect 14372 22967 14424 22976
rect 14372 22933 14381 22967
rect 14381 22933 14415 22967
rect 14415 22933 14424 22967
rect 14372 22924 14424 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 17224 22924 17276 22976
rect 18880 23103 18932 23112
rect 18880 23069 18889 23103
rect 18889 23069 18923 23103
rect 18923 23069 18932 23103
rect 18880 23060 18932 23069
rect 18512 22992 18564 23044
rect 19524 22992 19576 23044
rect 19800 23035 19852 23044
rect 19800 23001 19809 23035
rect 19809 23001 19843 23035
rect 19843 23001 19852 23035
rect 19800 22992 19852 23001
rect 21548 22992 21600 23044
rect 21824 23035 21876 23044
rect 21824 23001 21833 23035
rect 21833 23001 21867 23035
rect 21867 23001 21876 23035
rect 21824 22992 21876 23001
rect 21916 22992 21968 23044
rect 24676 22992 24728 23044
rect 24768 23035 24820 23044
rect 24768 23001 24777 23035
rect 24777 23001 24811 23035
rect 24811 23001 24820 23035
rect 24768 22992 24820 23001
rect 18788 22924 18840 22976
rect 22008 22924 22060 22976
rect 23296 22967 23348 22976
rect 23296 22933 23305 22967
rect 23305 22933 23339 22967
rect 23339 22933 23348 22967
rect 23296 22924 23348 22933
rect 23664 22967 23716 22976
rect 23664 22933 23673 22967
rect 23673 22933 23707 22967
rect 23707 22933 23716 22967
rect 23664 22924 23716 22933
rect 25320 22967 25372 22976
rect 25320 22933 25329 22967
rect 25329 22933 25363 22967
rect 25363 22933 25372 22967
rect 25320 22924 25372 22933
rect 25688 23103 25740 23112
rect 25688 23069 25697 23103
rect 25697 23069 25731 23103
rect 25731 23069 25740 23103
rect 25688 23060 25740 23069
rect 31300 23196 31352 23248
rect 32864 23196 32916 23248
rect 30196 23171 30248 23180
rect 30196 23137 30205 23171
rect 30205 23137 30239 23171
rect 30239 23137 30248 23171
rect 30196 23128 30248 23137
rect 30288 23171 30340 23180
rect 30288 23137 30297 23171
rect 30297 23137 30331 23171
rect 30331 23137 30340 23171
rect 30288 23128 30340 23137
rect 31024 23128 31076 23180
rect 31668 23128 31720 23180
rect 31760 23128 31812 23180
rect 33324 23128 33376 23180
rect 33784 23128 33836 23180
rect 34520 23128 34572 23180
rect 35716 23128 35768 23180
rect 39028 23264 39080 23316
rect 39304 23307 39356 23316
rect 39304 23273 39313 23307
rect 39313 23273 39347 23307
rect 39347 23273 39356 23307
rect 39304 23264 39356 23273
rect 41604 23264 41656 23316
rect 43536 23264 43588 23316
rect 43628 23264 43680 23316
rect 44548 23264 44600 23316
rect 44824 23264 44876 23316
rect 48228 23307 48280 23316
rect 48228 23273 48237 23307
rect 48237 23273 48271 23307
rect 48271 23273 48280 23307
rect 48228 23264 48280 23273
rect 38660 23128 38712 23180
rect 39212 23128 39264 23180
rect 27252 22992 27304 23044
rect 27620 22992 27672 23044
rect 32772 23060 32824 23112
rect 27436 22967 27488 22976
rect 27436 22933 27445 22967
rect 27445 22933 27479 22967
rect 27479 22933 27488 22967
rect 27436 22924 27488 22933
rect 29368 22967 29420 22976
rect 29368 22933 29377 22967
rect 29377 22933 29411 22967
rect 29411 22933 29420 22967
rect 29368 22924 29420 22933
rect 30104 22967 30156 22976
rect 30104 22933 30113 22967
rect 30113 22933 30147 22967
rect 30147 22933 30156 22967
rect 30104 22924 30156 22933
rect 30748 22924 30800 22976
rect 31208 22924 31260 22976
rect 34244 23060 34296 23112
rect 34980 23060 35032 23112
rect 33232 22992 33284 23044
rect 33784 22924 33836 22976
rect 34336 22992 34388 23044
rect 35624 22992 35676 23044
rect 35992 22992 36044 23044
rect 34520 22924 34572 22976
rect 34612 22924 34664 22976
rect 34796 22924 34848 22976
rect 37372 23060 37424 23112
rect 41052 23171 41104 23180
rect 41052 23137 41061 23171
rect 41061 23137 41095 23171
rect 41095 23137 41104 23171
rect 41052 23128 41104 23137
rect 42248 23196 42300 23248
rect 44272 23196 44324 23248
rect 47032 23196 47084 23248
rect 48596 23196 48648 23248
rect 37004 22992 37056 23044
rect 36912 22924 36964 22976
rect 38660 22992 38712 23044
rect 41512 23103 41564 23112
rect 41512 23069 41521 23103
rect 41521 23069 41555 23103
rect 41555 23069 41564 23103
rect 41512 23060 41564 23069
rect 42156 23060 42208 23112
rect 44180 23060 44232 23112
rect 44548 23060 44600 23112
rect 45376 23103 45428 23112
rect 45376 23069 45385 23103
rect 45385 23069 45419 23103
rect 45419 23069 45428 23103
rect 45376 23060 45428 23069
rect 48044 23128 48096 23180
rect 47584 23103 47636 23112
rect 47584 23069 47593 23103
rect 47593 23069 47627 23103
rect 47627 23069 47636 23103
rect 47584 23060 47636 23069
rect 49332 23103 49384 23112
rect 49332 23069 49341 23103
rect 49341 23069 49375 23103
rect 49375 23069 49384 23103
rect 49332 23060 49384 23069
rect 41236 22992 41288 23044
rect 39764 22924 39816 22976
rect 39948 22924 40000 22976
rect 40500 22967 40552 22976
rect 40500 22933 40509 22967
rect 40509 22933 40543 22967
rect 40543 22933 40552 22967
rect 40500 22924 40552 22933
rect 41052 22924 41104 22976
rect 44732 22992 44784 23044
rect 43352 22924 43404 22976
rect 46756 22924 46808 22976
rect 48320 22924 48372 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 1584 22720 1636 22772
rect 3424 22720 3476 22772
rect 4804 22695 4856 22704
rect 4804 22661 4813 22695
rect 4813 22661 4847 22695
rect 4847 22661 4856 22695
rect 4804 22652 4856 22661
rect 7564 22652 7616 22704
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 7196 22584 7248 22636
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 7104 22559 7156 22568
rect 7104 22525 7113 22559
rect 7113 22525 7147 22559
rect 7147 22525 7156 22559
rect 7104 22516 7156 22525
rect 7380 22516 7432 22568
rect 12624 22720 12676 22772
rect 13544 22720 13596 22772
rect 14188 22720 14240 22772
rect 14556 22763 14608 22772
rect 14556 22729 14565 22763
rect 14565 22729 14599 22763
rect 14599 22729 14608 22763
rect 14556 22720 14608 22729
rect 9956 22695 10008 22704
rect 9956 22661 9965 22695
rect 9965 22661 9999 22695
rect 9999 22661 10008 22695
rect 9956 22652 10008 22661
rect 12808 22695 12860 22704
rect 12808 22661 12817 22695
rect 12817 22661 12851 22695
rect 12851 22661 12860 22695
rect 12808 22652 12860 22661
rect 15108 22695 15160 22704
rect 15108 22661 15117 22695
rect 15117 22661 15151 22695
rect 15151 22661 15160 22695
rect 15108 22652 15160 22661
rect 11152 22627 11204 22636
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 11428 22584 11480 22636
rect 14648 22584 14700 22636
rect 18880 22720 18932 22772
rect 19340 22720 19392 22772
rect 21180 22763 21232 22772
rect 21180 22729 21189 22763
rect 21189 22729 21223 22763
rect 21223 22729 21232 22763
rect 21180 22720 21232 22729
rect 21824 22720 21876 22772
rect 22008 22720 22060 22772
rect 18512 22652 18564 22704
rect 19248 22652 19300 22704
rect 23940 22652 23992 22704
rect 2780 22448 2832 22500
rect 6460 22448 6512 22500
rect 9128 22448 9180 22500
rect 3792 22380 3844 22432
rect 6000 22380 6052 22432
rect 7748 22380 7800 22432
rect 15384 22448 15436 22500
rect 11980 22380 12032 22432
rect 12256 22423 12308 22432
rect 12256 22389 12265 22423
rect 12265 22389 12299 22423
rect 12299 22389 12308 22423
rect 12256 22380 12308 22389
rect 14372 22380 14424 22432
rect 16212 22380 16264 22432
rect 19340 22584 19392 22636
rect 20812 22584 20864 22636
rect 21548 22584 21600 22636
rect 21732 22584 21784 22636
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 23756 22584 23808 22636
rect 24952 22584 25004 22636
rect 25872 22652 25924 22704
rect 27252 22720 27304 22772
rect 27344 22763 27396 22772
rect 27344 22729 27353 22763
rect 27353 22729 27387 22763
rect 27387 22729 27396 22763
rect 27344 22720 27396 22729
rect 27436 22720 27488 22772
rect 29460 22652 29512 22704
rect 30012 22652 30064 22704
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 27252 22584 27304 22636
rect 28264 22584 28316 22636
rect 17132 22559 17184 22568
rect 17132 22525 17141 22559
rect 17141 22525 17175 22559
rect 17175 22525 17184 22559
rect 17132 22516 17184 22525
rect 18420 22516 18472 22568
rect 18328 22380 18380 22432
rect 23296 22516 23348 22568
rect 23664 22516 23716 22568
rect 21824 22448 21876 22500
rect 21640 22423 21692 22432
rect 21640 22389 21649 22423
rect 21649 22389 21683 22423
rect 21683 22389 21692 22423
rect 21640 22380 21692 22389
rect 23388 22448 23440 22500
rect 24860 22491 24912 22500
rect 24860 22457 24869 22491
rect 24869 22457 24903 22491
rect 24903 22457 24912 22491
rect 24860 22448 24912 22457
rect 26608 22559 26660 22568
rect 26608 22525 26617 22559
rect 26617 22525 26651 22559
rect 26651 22525 26660 22559
rect 26608 22516 26660 22525
rect 27528 22448 27580 22500
rect 27712 22448 27764 22500
rect 28080 22491 28132 22500
rect 28080 22457 28089 22491
rect 28089 22457 28123 22491
rect 28123 22457 28132 22491
rect 28080 22448 28132 22457
rect 23480 22380 23532 22432
rect 24032 22380 24084 22432
rect 24584 22423 24636 22432
rect 24584 22389 24593 22423
rect 24593 22389 24627 22423
rect 24627 22389 24636 22423
rect 24584 22380 24636 22389
rect 25136 22380 25188 22432
rect 26332 22380 26384 22432
rect 28908 22516 28960 22568
rect 30380 22516 30432 22568
rect 30840 22720 30892 22772
rect 33232 22720 33284 22772
rect 30656 22627 30708 22636
rect 30656 22593 30665 22627
rect 30665 22593 30699 22627
rect 30699 22593 30708 22627
rect 30656 22584 30708 22593
rect 30748 22627 30800 22636
rect 30748 22593 30757 22627
rect 30757 22593 30791 22627
rect 30791 22593 30800 22627
rect 30748 22584 30800 22593
rect 33600 22652 33652 22704
rect 34980 22720 35032 22772
rect 35440 22763 35492 22772
rect 35440 22729 35449 22763
rect 35449 22729 35483 22763
rect 35483 22729 35492 22763
rect 35440 22720 35492 22729
rect 35900 22720 35952 22772
rect 33876 22652 33928 22704
rect 34612 22652 34664 22704
rect 36360 22652 36412 22704
rect 37280 22652 37332 22704
rect 30012 22448 30064 22500
rect 31208 22448 31260 22500
rect 35532 22584 35584 22636
rect 34428 22516 34480 22568
rect 30196 22380 30248 22432
rect 30472 22380 30524 22432
rect 30840 22380 30892 22432
rect 31484 22423 31536 22432
rect 31484 22389 31493 22423
rect 31493 22389 31527 22423
rect 31527 22389 31536 22423
rect 31484 22380 31536 22389
rect 33692 22448 33744 22500
rect 38660 22720 38712 22772
rect 38936 22720 38988 22772
rect 38844 22652 38896 22704
rect 44456 22720 44508 22772
rect 47584 22720 47636 22772
rect 37832 22584 37884 22636
rect 39212 22627 39264 22636
rect 39212 22593 39221 22627
rect 39221 22593 39255 22627
rect 39255 22593 39264 22627
rect 39212 22584 39264 22593
rect 39764 22627 39816 22636
rect 39764 22593 39773 22627
rect 39773 22593 39807 22627
rect 39807 22593 39816 22627
rect 39764 22584 39816 22593
rect 40408 22627 40460 22636
rect 40408 22593 40417 22627
rect 40417 22593 40451 22627
rect 40451 22593 40460 22627
rect 40408 22584 40460 22593
rect 41144 22584 41196 22636
rect 41604 22584 41656 22636
rect 42616 22627 42668 22636
rect 42616 22593 42625 22627
rect 42625 22593 42659 22627
rect 42659 22593 42668 22627
rect 42616 22584 42668 22593
rect 44088 22652 44140 22704
rect 44732 22652 44784 22704
rect 45744 22695 45796 22704
rect 45744 22661 45753 22695
rect 45753 22661 45787 22695
rect 45787 22661 45796 22695
rect 45744 22652 45796 22661
rect 47308 22652 47360 22704
rect 47860 22652 47912 22704
rect 44180 22584 44232 22636
rect 49148 22584 49200 22636
rect 49240 22584 49292 22636
rect 37648 22516 37700 22568
rect 38844 22516 38896 22568
rect 33968 22380 34020 22432
rect 34520 22380 34572 22432
rect 36452 22448 36504 22500
rect 35808 22380 35860 22432
rect 37556 22448 37608 22500
rect 39304 22448 39356 22500
rect 36912 22380 36964 22432
rect 40684 22516 40736 22568
rect 39488 22448 39540 22500
rect 43996 22559 44048 22568
rect 43996 22525 44005 22559
rect 44005 22525 44039 22559
rect 44039 22525 44048 22559
rect 43996 22516 44048 22525
rect 46664 22516 46716 22568
rect 47584 22516 47636 22568
rect 47860 22516 47912 22568
rect 44548 22448 44600 22500
rect 45008 22491 45060 22500
rect 45008 22457 45017 22491
rect 45017 22457 45051 22491
rect 45051 22457 45060 22491
rect 45008 22448 45060 22457
rect 40040 22423 40092 22432
rect 40040 22389 40049 22423
rect 40049 22389 40083 22423
rect 40083 22389 40092 22423
rect 40040 22380 40092 22389
rect 40316 22380 40368 22432
rect 45284 22380 45336 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 4252 22176 4304 22228
rect 11888 22176 11940 22228
rect 3976 22108 4028 22160
rect 3516 22040 3568 22092
rect 3792 22040 3844 22092
rect 1032 21904 1084 21956
rect 5356 22015 5408 22024
rect 5356 21981 5365 22015
rect 5365 21981 5399 22015
rect 5399 21981 5408 22015
rect 5356 21972 5408 21981
rect 9680 22040 9732 22092
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 11980 22040 12032 22092
rect 17132 22176 17184 22228
rect 19800 22176 19852 22228
rect 27068 22176 27120 22228
rect 27620 22176 27672 22228
rect 14372 22108 14424 22160
rect 17040 22108 17092 22160
rect 19708 22108 19760 22160
rect 18972 22040 19024 22092
rect 23480 22108 23532 22160
rect 22652 22040 22704 22092
rect 23388 22040 23440 22092
rect 24860 22108 24912 22160
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 26608 22108 26660 22160
rect 27160 22108 27212 22160
rect 30656 22176 30708 22228
rect 31484 22176 31536 22228
rect 31668 22176 31720 22228
rect 34244 22219 34296 22228
rect 34244 22185 34253 22219
rect 34253 22185 34287 22219
rect 34287 22185 34296 22219
rect 34244 22176 34296 22185
rect 29736 22151 29788 22160
rect 29736 22117 29745 22151
rect 29745 22117 29779 22151
rect 29779 22117 29788 22151
rect 29736 22108 29788 22117
rect 28080 22040 28132 22092
rect 28908 22083 28960 22092
rect 28908 22049 28917 22083
rect 28917 22049 28951 22083
rect 28951 22049 28960 22083
rect 28908 22040 28960 22049
rect 3516 21904 3568 21956
rect 5632 21904 5684 21956
rect 8484 21904 8536 21956
rect 8300 21836 8352 21888
rect 8392 21879 8444 21888
rect 8392 21845 8401 21879
rect 8401 21845 8435 21879
rect 8435 21845 8444 21879
rect 8392 21836 8444 21845
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 13728 21972 13780 22024
rect 16948 22015 17000 22024
rect 16948 21981 16957 22015
rect 16957 21981 16991 22015
rect 16991 21981 17000 22015
rect 16948 21972 17000 21981
rect 11428 21904 11480 21956
rect 12716 21904 12768 21956
rect 14648 21947 14700 21956
rect 14648 21913 14657 21947
rect 14657 21913 14691 21947
rect 14691 21913 14700 21947
rect 14648 21904 14700 21913
rect 16212 21904 16264 21956
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 15292 21836 15344 21888
rect 16672 21947 16724 21956
rect 16672 21913 16681 21947
rect 16681 21913 16715 21947
rect 16715 21913 16724 21947
rect 16672 21904 16724 21913
rect 18512 21972 18564 22024
rect 17224 21904 17276 21956
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 22284 21972 22336 22024
rect 22928 21972 22980 22024
rect 23940 21972 23992 22024
rect 24860 21972 24912 22024
rect 25596 21972 25648 22024
rect 21732 21904 21784 21956
rect 18972 21836 19024 21888
rect 21456 21879 21508 21888
rect 21456 21845 21465 21879
rect 21465 21845 21499 21879
rect 21499 21845 21508 21879
rect 21456 21836 21508 21845
rect 23480 21904 23532 21956
rect 23572 21904 23624 21956
rect 22468 21836 22520 21888
rect 22560 21836 22612 21888
rect 22928 21836 22980 21888
rect 23664 21836 23716 21888
rect 26056 21904 26108 21956
rect 30196 22040 30248 22092
rect 31576 22040 31628 22092
rect 32772 22040 32824 22092
rect 35440 22108 35492 22160
rect 33968 22040 34020 22092
rect 35900 22040 35952 22092
rect 39120 22176 39172 22228
rect 39212 22176 39264 22228
rect 39580 22219 39632 22228
rect 36820 22151 36872 22160
rect 36820 22117 36829 22151
rect 36829 22117 36863 22151
rect 36863 22117 36872 22151
rect 36820 22108 36872 22117
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 30380 21972 30432 22024
rect 30840 22015 30892 22024
rect 30840 21981 30849 22015
rect 30849 21981 30883 22015
rect 30883 21981 30892 22015
rect 30840 21972 30892 21981
rect 32220 21972 32272 22024
rect 37096 22040 37148 22092
rect 37648 22040 37700 22092
rect 26884 21904 26936 21956
rect 27804 21904 27856 21956
rect 28540 21904 28592 21956
rect 28724 21947 28776 21956
rect 28724 21913 28733 21947
rect 28733 21913 28767 21947
rect 28767 21913 28776 21947
rect 28724 21904 28776 21913
rect 30472 21904 30524 21956
rect 31208 21904 31260 21956
rect 24768 21836 24820 21888
rect 25320 21836 25372 21888
rect 25780 21836 25832 21888
rect 26700 21836 26752 21888
rect 29644 21836 29696 21888
rect 30380 21879 30432 21888
rect 30380 21845 30389 21879
rect 30389 21845 30423 21879
rect 30423 21845 30432 21879
rect 30380 21836 30432 21845
rect 30748 21836 30800 21888
rect 33692 21904 33744 21956
rect 37832 22040 37884 22092
rect 39580 22185 39589 22219
rect 39589 22185 39623 22219
rect 39623 22185 39632 22219
rect 39580 22176 39632 22185
rect 40500 22176 40552 22228
rect 44732 22219 44784 22228
rect 44732 22185 44741 22219
rect 44741 22185 44775 22219
rect 44775 22185 44784 22219
rect 44732 22176 44784 22185
rect 47032 22176 47084 22228
rect 39856 22151 39908 22160
rect 39856 22117 39865 22151
rect 39865 22117 39899 22151
rect 39899 22117 39908 22151
rect 39856 22108 39908 22117
rect 34612 21904 34664 21956
rect 36544 21904 36596 21956
rect 32496 21836 32548 21888
rect 32680 21836 32732 21888
rect 33416 21879 33468 21888
rect 33416 21845 33425 21879
rect 33425 21845 33459 21879
rect 33459 21845 33468 21879
rect 33416 21836 33468 21845
rect 35164 21879 35216 21888
rect 35164 21845 35173 21879
rect 35173 21845 35207 21879
rect 35207 21845 35216 21879
rect 35164 21836 35216 21845
rect 35256 21879 35308 21888
rect 35256 21845 35265 21879
rect 35265 21845 35299 21879
rect 35299 21845 35308 21879
rect 35256 21836 35308 21845
rect 36176 21836 36228 21888
rect 36360 21879 36412 21888
rect 36360 21845 36369 21879
rect 36369 21845 36403 21879
rect 36403 21845 36412 21879
rect 36360 21836 36412 21845
rect 37372 21879 37424 21888
rect 37372 21845 37381 21879
rect 37381 21845 37415 21879
rect 37415 21845 37424 21879
rect 37372 21836 37424 21845
rect 38844 21947 38896 21956
rect 38844 21913 38853 21947
rect 38853 21913 38887 21947
rect 38887 21913 38896 21947
rect 38844 21904 38896 21913
rect 39304 21836 39356 21888
rect 40316 22040 40368 22092
rect 40684 22083 40736 22092
rect 40684 22049 40693 22083
rect 40693 22049 40727 22083
rect 40727 22049 40736 22083
rect 40684 22040 40736 22049
rect 41972 22040 42024 22092
rect 42156 22040 42208 22092
rect 45284 22108 45336 22160
rect 42800 22040 42852 22092
rect 44548 22083 44600 22092
rect 44548 22049 44557 22083
rect 44557 22049 44591 22083
rect 44591 22049 44600 22083
rect 44548 22040 44600 22049
rect 45192 22083 45244 22092
rect 45192 22049 45201 22083
rect 45201 22049 45235 22083
rect 45235 22049 45244 22083
rect 45192 22040 45244 22049
rect 46848 22040 46900 22092
rect 47676 22040 47728 22092
rect 40684 21904 40736 21956
rect 42616 21904 42668 21956
rect 40592 21879 40644 21888
rect 40592 21845 40601 21879
rect 40601 21845 40635 21879
rect 40635 21845 40644 21879
rect 40592 21836 40644 21845
rect 41236 21836 41288 21888
rect 41696 21836 41748 21888
rect 43444 21972 43496 22024
rect 44180 22015 44232 22024
rect 44180 21981 44189 22015
rect 44189 21981 44223 22015
rect 44223 21981 44232 22015
rect 44180 21972 44232 21981
rect 45468 22015 45520 22024
rect 45468 21981 45477 22015
rect 45477 21981 45511 22015
rect 45511 21981 45520 22015
rect 45468 21972 45520 21981
rect 46756 22015 46808 22024
rect 46756 21981 46765 22015
rect 46765 21981 46799 22015
rect 46799 21981 46808 22015
rect 46756 21972 46808 21981
rect 49516 22040 49568 22092
rect 49332 22015 49384 22024
rect 42800 21904 42852 21956
rect 45836 21904 45888 21956
rect 47492 21904 47544 21956
rect 49332 21981 49341 22015
rect 49341 21981 49375 22015
rect 49375 21981 49384 22015
rect 49332 21972 49384 21981
rect 45008 21836 45060 21888
rect 46572 21879 46624 21888
rect 46572 21845 46581 21879
rect 46581 21845 46615 21879
rect 46615 21845 46624 21879
rect 46572 21836 46624 21845
rect 48688 21879 48740 21888
rect 48688 21845 48697 21879
rect 48697 21845 48731 21879
rect 48731 21845 48740 21879
rect 48688 21836 48740 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 5356 21632 5408 21684
rect 3332 21564 3384 21616
rect 3700 21564 3752 21616
rect 9588 21632 9640 21684
rect 11520 21632 11572 21684
rect 12624 21632 12676 21684
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 14004 21632 14056 21684
rect 20996 21632 21048 21684
rect 1768 21471 1820 21480
rect 1768 21437 1777 21471
rect 1777 21437 1811 21471
rect 1811 21437 1820 21471
rect 1768 21428 1820 21437
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 6368 21496 6420 21548
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 5816 21428 5868 21480
rect 12256 21496 12308 21548
rect 12808 21564 12860 21616
rect 12624 21496 12676 21548
rect 11428 21428 11480 21480
rect 12440 21428 12492 21480
rect 13912 21496 13964 21548
rect 14280 21564 14332 21616
rect 16212 21564 16264 21616
rect 17224 21564 17276 21616
rect 11796 21360 11848 21412
rect 12348 21360 12400 21412
rect 7656 21292 7708 21344
rect 11704 21292 11756 21344
rect 11980 21292 12032 21344
rect 14004 21360 14056 21412
rect 13728 21292 13780 21344
rect 18328 21496 18380 21548
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 15292 21428 15344 21480
rect 16764 21428 16816 21480
rect 18788 21564 18840 21616
rect 19432 21564 19484 21616
rect 20628 21564 20680 21616
rect 22836 21632 22888 21684
rect 21548 21564 21600 21616
rect 25412 21632 25464 21684
rect 24124 21564 24176 21616
rect 27620 21632 27672 21684
rect 28724 21632 28776 21684
rect 30564 21632 30616 21684
rect 17040 21360 17092 21412
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 18972 21428 19024 21480
rect 15936 21292 15988 21344
rect 16580 21292 16632 21344
rect 17500 21292 17552 21344
rect 21364 21360 21416 21412
rect 22192 21428 22244 21480
rect 22836 21428 22888 21480
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25136 21496 25188 21505
rect 24584 21428 24636 21480
rect 25228 21471 25280 21480
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 19340 21292 19392 21344
rect 19432 21292 19484 21344
rect 21640 21292 21692 21344
rect 22192 21335 22244 21344
rect 22192 21301 22201 21335
rect 22201 21301 22235 21335
rect 22235 21301 22244 21335
rect 22192 21292 22244 21301
rect 22468 21292 22520 21344
rect 26976 21496 27028 21548
rect 29828 21564 29880 21616
rect 31208 21632 31260 21684
rect 33416 21632 33468 21684
rect 33600 21675 33652 21684
rect 33600 21641 33609 21675
rect 33609 21641 33643 21675
rect 33643 21641 33652 21675
rect 33600 21632 33652 21641
rect 34796 21675 34848 21684
rect 34796 21641 34805 21675
rect 34805 21641 34839 21675
rect 34839 21641 34848 21675
rect 34796 21632 34848 21641
rect 35072 21632 35124 21684
rect 32588 21564 32640 21616
rect 35624 21564 35676 21616
rect 40040 21632 40092 21684
rect 40960 21632 41012 21684
rect 41328 21632 41380 21684
rect 25412 21471 25464 21480
rect 25412 21437 25421 21471
rect 25421 21437 25455 21471
rect 25455 21437 25464 21471
rect 25412 21428 25464 21437
rect 26056 21471 26108 21480
rect 26056 21437 26065 21471
rect 26065 21437 26099 21471
rect 26099 21437 26108 21471
rect 26056 21428 26108 21437
rect 27344 21428 27396 21480
rect 27896 21496 27948 21548
rect 28816 21471 28868 21480
rect 28816 21437 28825 21471
rect 28825 21437 28859 21471
rect 28859 21437 28868 21471
rect 28816 21428 28868 21437
rect 28908 21471 28960 21480
rect 28908 21437 28917 21471
rect 28917 21437 28951 21471
rect 28951 21437 28960 21471
rect 28908 21428 28960 21437
rect 29460 21360 29512 21412
rect 30932 21496 30984 21548
rect 33508 21539 33560 21548
rect 33508 21505 33517 21539
rect 33517 21505 33551 21539
rect 33551 21505 33560 21539
rect 33508 21496 33560 21505
rect 33692 21496 33744 21548
rect 37280 21607 37332 21616
rect 37280 21573 37289 21607
rect 37289 21573 37323 21607
rect 37323 21573 37332 21607
rect 37280 21564 37332 21573
rect 37832 21564 37884 21616
rect 38568 21564 38620 21616
rect 39764 21564 39816 21616
rect 42616 21675 42668 21684
rect 42616 21641 42625 21675
rect 42625 21641 42659 21675
rect 42659 21641 42668 21675
rect 42616 21632 42668 21641
rect 44456 21632 44508 21684
rect 49240 21632 49292 21684
rect 44640 21564 44692 21616
rect 47032 21564 47084 21616
rect 48688 21564 48740 21616
rect 37556 21539 37608 21548
rect 30288 21428 30340 21480
rect 30748 21428 30800 21480
rect 30564 21360 30616 21412
rect 25136 21292 25188 21344
rect 25872 21335 25924 21344
rect 25872 21301 25881 21335
rect 25881 21301 25915 21335
rect 25915 21301 25924 21335
rect 25872 21292 25924 21301
rect 26056 21292 26108 21344
rect 27252 21292 27304 21344
rect 30196 21292 30248 21344
rect 35992 21428 36044 21480
rect 36176 21471 36228 21480
rect 36176 21437 36185 21471
rect 36185 21437 36219 21471
rect 36219 21437 36228 21471
rect 36176 21428 36228 21437
rect 36268 21471 36320 21480
rect 36268 21437 36277 21471
rect 36277 21437 36311 21471
rect 36311 21437 36320 21471
rect 36268 21428 36320 21437
rect 37556 21505 37565 21539
rect 37565 21505 37599 21539
rect 37599 21505 37608 21539
rect 37556 21496 37608 21505
rect 40224 21496 40276 21548
rect 42432 21496 42484 21548
rect 43352 21496 43404 21548
rect 43812 21496 43864 21548
rect 45192 21496 45244 21548
rect 47400 21496 47452 21548
rect 47584 21496 47636 21548
rect 49240 21496 49292 21548
rect 37188 21428 37240 21480
rect 37924 21428 37976 21480
rect 38292 21471 38344 21480
rect 38292 21437 38301 21471
rect 38301 21437 38335 21471
rect 38335 21437 38344 21471
rect 38292 21428 38344 21437
rect 39580 21428 39632 21480
rect 39764 21471 39816 21480
rect 39764 21437 39773 21471
rect 39773 21437 39807 21471
rect 39807 21437 39816 21471
rect 39764 21428 39816 21437
rect 41052 21428 41104 21480
rect 41512 21471 41564 21480
rect 41512 21437 41521 21471
rect 41521 21437 41555 21471
rect 41555 21437 41564 21471
rect 41512 21428 41564 21437
rect 44272 21428 44324 21480
rect 34244 21360 34296 21412
rect 36544 21360 36596 21412
rect 36636 21360 36688 21412
rect 33508 21292 33560 21344
rect 34980 21292 35032 21344
rect 35164 21335 35216 21344
rect 35164 21301 35173 21335
rect 35173 21301 35207 21335
rect 35207 21301 35216 21335
rect 35164 21292 35216 21301
rect 35716 21335 35768 21344
rect 35716 21301 35725 21335
rect 35725 21301 35759 21335
rect 35759 21301 35768 21335
rect 35716 21292 35768 21301
rect 35992 21292 36044 21344
rect 37004 21292 37056 21344
rect 37280 21292 37332 21344
rect 37648 21335 37700 21344
rect 37648 21301 37657 21335
rect 37657 21301 37691 21335
rect 37691 21301 37700 21335
rect 37648 21292 37700 21301
rect 39488 21360 39540 21412
rect 40868 21335 40920 21344
rect 40868 21301 40877 21335
rect 40877 21301 40911 21335
rect 40911 21301 40920 21335
rect 40868 21292 40920 21301
rect 42800 21292 42852 21344
rect 43536 21292 43588 21344
rect 47768 21471 47820 21480
rect 47768 21437 47777 21471
rect 47777 21437 47811 21471
rect 47811 21437 47820 21471
rect 47768 21428 47820 21437
rect 46296 21360 46348 21412
rect 47216 21360 47268 21412
rect 47400 21292 47452 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 2872 20952 2924 21004
rect 4160 20995 4212 21004
rect 4160 20961 4169 20995
rect 4169 20961 4203 20995
rect 4203 20961 4212 20995
rect 4160 20952 4212 20961
rect 5264 20884 5316 20936
rect 12440 21088 12492 21140
rect 14280 21131 14332 21140
rect 14280 21097 14289 21131
rect 14289 21097 14323 21131
rect 14323 21097 14332 21131
rect 14280 21088 14332 21097
rect 7840 21020 7892 21072
rect 10416 21020 10468 21072
rect 11980 21020 12032 21072
rect 12164 21020 12216 21072
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 6368 20952 6420 21004
rect 9956 20952 10008 21004
rect 13360 20952 13412 21004
rect 7196 20748 7248 20800
rect 7472 20791 7524 20800
rect 7472 20757 7481 20791
rect 7481 20757 7515 20791
rect 7515 20757 7524 20791
rect 7472 20748 7524 20757
rect 8392 20927 8444 20936
rect 8392 20893 8401 20927
rect 8401 20893 8435 20927
rect 8435 20893 8444 20927
rect 8392 20884 8444 20893
rect 8576 20884 8628 20936
rect 11152 20884 11204 20936
rect 11336 20927 11388 20936
rect 11336 20893 11345 20927
rect 11345 20893 11379 20927
rect 11379 20893 11388 20927
rect 11336 20884 11388 20893
rect 11796 20884 11848 20936
rect 12164 20884 12216 20936
rect 8484 20816 8536 20868
rect 10600 20748 10652 20800
rect 11060 20748 11112 20800
rect 11244 20748 11296 20800
rect 12348 20859 12400 20868
rect 12348 20825 12357 20859
rect 12357 20825 12391 20859
rect 12391 20825 12400 20859
rect 12348 20816 12400 20825
rect 12808 20816 12860 20868
rect 24308 21088 24360 21140
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 24952 21088 25004 21140
rect 14556 20952 14608 21004
rect 18512 20952 18564 21004
rect 19708 20952 19760 21004
rect 19800 20952 19852 21004
rect 23296 21020 23348 21072
rect 23480 21020 23532 21072
rect 26056 21020 26108 21072
rect 17040 20884 17092 20936
rect 19340 20884 19392 20936
rect 13728 20748 13780 20800
rect 16120 20816 16172 20868
rect 16212 20748 16264 20800
rect 16304 20748 16356 20800
rect 18420 20748 18472 20800
rect 19432 20748 19484 20800
rect 22560 20952 22612 21004
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 27252 21020 27304 21072
rect 22928 20927 22980 20936
rect 22928 20893 22937 20927
rect 22937 20893 22971 20927
rect 22971 20893 22980 20927
rect 22928 20884 22980 20893
rect 19616 20791 19668 20800
rect 19616 20757 19625 20791
rect 19625 20757 19659 20791
rect 19659 20757 19668 20791
rect 19616 20748 19668 20757
rect 22192 20816 22244 20868
rect 24308 20884 24360 20936
rect 26240 20995 26292 21004
rect 26240 20961 26249 20995
rect 26249 20961 26283 20995
rect 26283 20961 26292 20995
rect 26240 20952 26292 20961
rect 26424 20952 26476 21004
rect 27160 20952 27212 21004
rect 24768 20884 24820 20936
rect 23572 20859 23624 20868
rect 23572 20825 23581 20859
rect 23581 20825 23615 20859
rect 23615 20825 23624 20859
rect 23572 20816 23624 20825
rect 24124 20816 24176 20868
rect 24676 20816 24728 20868
rect 25780 20816 25832 20868
rect 25412 20748 25464 20800
rect 26516 20884 26568 20936
rect 29736 21131 29788 21140
rect 29736 21097 29745 21131
rect 29745 21097 29779 21131
rect 29779 21097 29788 21131
rect 29736 21088 29788 21097
rect 30656 21088 30708 21140
rect 31024 21088 31076 21140
rect 30104 21020 30156 21072
rect 27896 20995 27948 21004
rect 27896 20961 27905 20995
rect 27905 20961 27939 20995
rect 27939 20961 27948 20995
rect 27896 20952 27948 20961
rect 35716 21088 35768 21140
rect 36728 21088 36780 21140
rect 37648 21131 37700 21140
rect 37648 21097 37657 21131
rect 37657 21097 37691 21131
rect 37691 21097 37700 21131
rect 37648 21088 37700 21097
rect 37740 21088 37792 21140
rect 34060 21020 34112 21072
rect 35072 21020 35124 21072
rect 37372 21020 37424 21072
rect 38108 21020 38160 21072
rect 39580 21088 39632 21140
rect 28724 20927 28776 20936
rect 28724 20893 28733 20927
rect 28733 20893 28767 20927
rect 28767 20893 28776 20927
rect 28724 20884 28776 20893
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 32312 20952 32364 21004
rect 33968 20952 34020 21004
rect 34244 20995 34296 21004
rect 34244 20961 34253 20995
rect 34253 20961 34287 20995
rect 34287 20961 34296 20995
rect 34244 20952 34296 20961
rect 35900 20952 35952 21004
rect 36912 20952 36964 21004
rect 32404 20884 32456 20936
rect 32496 20927 32548 20936
rect 32496 20893 32505 20927
rect 32505 20893 32539 20927
rect 32539 20893 32548 20927
rect 32496 20884 32548 20893
rect 34612 20884 34664 20936
rect 35256 20884 35308 20936
rect 26792 20816 26844 20868
rect 27344 20859 27396 20868
rect 27344 20825 27353 20859
rect 27353 20825 27387 20859
rect 27387 20825 27396 20859
rect 27344 20816 27396 20825
rect 28816 20816 28868 20868
rect 30472 20816 30524 20868
rect 30932 20816 30984 20868
rect 31760 20816 31812 20868
rect 31852 20816 31904 20868
rect 32864 20816 32916 20868
rect 37924 20952 37976 21004
rect 39488 20952 39540 21004
rect 39764 20952 39816 21004
rect 30012 20748 30064 20800
rect 30104 20748 30156 20800
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 32220 20748 32272 20800
rect 33692 20748 33744 20800
rect 37556 20816 37608 20868
rect 39120 20859 39172 20868
rect 39120 20825 39129 20859
rect 39129 20825 39163 20859
rect 39163 20825 39172 20859
rect 39120 20816 39172 20825
rect 39764 20816 39816 20868
rect 36268 20748 36320 20800
rect 36912 20791 36964 20800
rect 36912 20757 36921 20791
rect 36921 20757 36955 20791
rect 36955 20757 36964 20791
rect 36912 20748 36964 20757
rect 37280 20791 37332 20800
rect 37280 20757 37289 20791
rect 37289 20757 37323 20791
rect 37323 20757 37332 20791
rect 37280 20748 37332 20757
rect 37740 20748 37792 20800
rect 38752 20748 38804 20800
rect 41696 21088 41748 21140
rect 43536 21088 43588 21140
rect 43812 21088 43864 21140
rect 44456 21131 44508 21140
rect 44456 21097 44465 21131
rect 44465 21097 44499 21131
rect 44499 21097 44508 21131
rect 44456 21088 44508 21097
rect 45192 21131 45244 21140
rect 45192 21097 45201 21131
rect 45201 21097 45235 21131
rect 45235 21097 45244 21131
rect 45192 21088 45244 21097
rect 45836 21131 45888 21140
rect 45836 21097 45845 21131
rect 45845 21097 45879 21131
rect 45879 21097 45888 21131
rect 45836 21088 45888 21097
rect 40868 21020 40920 21072
rect 42432 20995 42484 21004
rect 42432 20961 42441 20995
rect 42441 20961 42475 20995
rect 42475 20961 42484 20995
rect 42432 20952 42484 20961
rect 43352 21020 43404 21072
rect 44364 21020 44416 21072
rect 45376 21020 45428 21072
rect 45376 20927 45428 20936
rect 45376 20893 45385 20927
rect 45385 20893 45419 20927
rect 45419 20893 45428 20927
rect 45376 20884 45428 20893
rect 46848 21020 46900 21072
rect 48320 20952 48372 21004
rect 47860 20884 47912 20936
rect 49332 20927 49384 20936
rect 49332 20893 49341 20927
rect 49341 20893 49375 20927
rect 49375 20893 49384 20927
rect 49332 20884 49384 20893
rect 40132 20816 40184 20868
rect 44180 20816 44232 20868
rect 41328 20748 41380 20800
rect 43352 20748 43404 20800
rect 47308 20791 47360 20800
rect 47308 20757 47317 20791
rect 47317 20757 47351 20791
rect 47351 20757 47360 20791
rect 47308 20748 47360 20757
rect 47400 20748 47452 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 6552 20544 6604 20596
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 11060 20544 11112 20596
rect 1308 20476 1360 20528
rect 8300 20476 8352 20528
rect 13544 20476 13596 20528
rect 13636 20476 13688 20528
rect 15568 20587 15620 20596
rect 15568 20553 15577 20587
rect 15577 20553 15611 20587
rect 15611 20553 15620 20587
rect 15568 20544 15620 20553
rect 15844 20544 15896 20596
rect 16028 20587 16080 20596
rect 16028 20553 16037 20587
rect 16037 20553 16071 20587
rect 16071 20553 16080 20587
rect 16028 20544 16080 20553
rect 17132 20544 17184 20596
rect 18880 20544 18932 20596
rect 19708 20587 19760 20596
rect 19708 20553 19717 20587
rect 19717 20553 19751 20587
rect 19751 20553 19760 20587
rect 19708 20544 19760 20553
rect 19892 20544 19944 20596
rect 2780 20272 2832 20324
rect 6460 20408 6512 20460
rect 9772 20408 9824 20460
rect 10416 20408 10468 20460
rect 11520 20408 11572 20460
rect 11704 20408 11756 20460
rect 12440 20408 12492 20460
rect 12900 20408 12952 20460
rect 13360 20408 13412 20460
rect 13728 20408 13780 20460
rect 13820 20408 13872 20460
rect 16212 20476 16264 20528
rect 22284 20544 22336 20596
rect 22928 20544 22980 20596
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 6368 20340 6420 20392
rect 6644 20340 6696 20392
rect 8392 20340 8444 20392
rect 11060 20340 11112 20392
rect 11152 20340 11204 20392
rect 4528 20204 4580 20256
rect 10140 20272 10192 20324
rect 11060 20204 11112 20256
rect 11612 20204 11664 20256
rect 11888 20204 11940 20256
rect 13452 20247 13504 20256
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 14280 20383 14332 20392
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 19432 20408 19484 20460
rect 22100 20408 22152 20460
rect 23664 20476 23716 20528
rect 17408 20340 17460 20392
rect 20444 20340 20496 20392
rect 21548 20340 21600 20392
rect 16856 20272 16908 20324
rect 16488 20204 16540 20256
rect 17132 20204 17184 20256
rect 17316 20204 17368 20256
rect 20076 20272 20128 20324
rect 19616 20204 19668 20256
rect 19984 20204 20036 20256
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 23756 20408 23808 20460
rect 25688 20544 25740 20596
rect 24032 20476 24084 20528
rect 24216 20476 24268 20528
rect 24584 20476 24636 20528
rect 25872 20476 25924 20528
rect 25964 20408 26016 20460
rect 22744 20272 22796 20324
rect 25596 20383 25648 20392
rect 25596 20349 25605 20383
rect 25605 20349 25639 20383
rect 25639 20349 25648 20383
rect 25596 20340 25648 20349
rect 30840 20544 30892 20596
rect 31484 20544 31536 20596
rect 32496 20544 32548 20596
rect 28264 20476 28316 20528
rect 29644 20476 29696 20528
rect 28540 20340 28592 20392
rect 29092 20340 29144 20392
rect 29460 20340 29512 20392
rect 30104 20340 30156 20392
rect 26056 20272 26108 20324
rect 26148 20272 26200 20324
rect 29368 20272 29420 20324
rect 25504 20204 25556 20256
rect 26424 20204 26476 20256
rect 27344 20204 27396 20256
rect 30288 20272 30340 20324
rect 31576 20476 31628 20528
rect 31668 20476 31720 20528
rect 30656 20340 30708 20392
rect 32220 20476 32272 20528
rect 31852 20340 31904 20392
rect 31944 20383 31996 20392
rect 31944 20349 31953 20383
rect 31953 20349 31987 20383
rect 31987 20349 31996 20383
rect 31944 20340 31996 20349
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 32588 20340 32640 20392
rect 33416 20340 33468 20392
rect 33692 20340 33744 20392
rect 36176 20544 36228 20596
rect 34520 20340 34572 20392
rect 35900 20476 35952 20528
rect 34888 20451 34940 20460
rect 34888 20417 34897 20451
rect 34897 20417 34931 20451
rect 34931 20417 34940 20451
rect 36912 20544 36964 20596
rect 37096 20544 37148 20596
rect 37188 20476 37240 20528
rect 37740 20476 37792 20528
rect 37924 20476 37976 20528
rect 43628 20544 43680 20596
rect 43904 20544 43956 20596
rect 46204 20544 46256 20596
rect 46480 20587 46532 20596
rect 46480 20553 46489 20587
rect 46489 20553 46523 20587
rect 46523 20553 46532 20587
rect 46480 20544 46532 20553
rect 46848 20544 46900 20596
rect 47676 20587 47728 20596
rect 47676 20553 47685 20587
rect 47685 20553 47719 20587
rect 47719 20553 47728 20587
rect 47676 20544 47728 20553
rect 34888 20408 34940 20417
rect 37464 20408 37516 20460
rect 39488 20451 39540 20460
rect 39488 20417 39497 20451
rect 39497 20417 39531 20451
rect 39531 20417 39540 20451
rect 39488 20408 39540 20417
rect 39764 20408 39816 20460
rect 34796 20383 34848 20392
rect 34796 20349 34805 20383
rect 34805 20349 34839 20383
rect 34839 20349 34848 20383
rect 34796 20340 34848 20349
rect 35072 20340 35124 20392
rect 37280 20340 37332 20392
rect 37648 20340 37700 20392
rect 40132 20383 40184 20392
rect 40132 20349 40141 20383
rect 40141 20349 40175 20383
rect 40175 20349 40184 20383
rect 40132 20340 40184 20349
rect 46480 20408 46532 20460
rect 47216 20451 47268 20460
rect 47216 20417 47225 20451
rect 47225 20417 47259 20451
rect 47259 20417 47268 20451
rect 47216 20408 47268 20417
rect 49332 20451 49384 20460
rect 49332 20417 49341 20451
rect 49341 20417 49375 20451
rect 49375 20417 49384 20451
rect 49332 20408 49384 20417
rect 46204 20340 46256 20392
rect 30564 20204 30616 20256
rect 30840 20204 30892 20256
rect 35256 20204 35308 20256
rect 36084 20247 36136 20256
rect 36084 20213 36093 20247
rect 36093 20213 36127 20247
rect 36127 20213 36136 20247
rect 36084 20204 36136 20213
rect 37648 20204 37700 20256
rect 37740 20247 37792 20256
rect 37740 20213 37749 20247
rect 37749 20213 37783 20247
rect 37783 20213 37792 20247
rect 37740 20204 37792 20213
rect 42800 20272 42852 20324
rect 49332 20272 49384 20324
rect 40684 20247 40736 20256
rect 40684 20213 40693 20247
rect 40693 20213 40727 20247
rect 40727 20213 40736 20247
rect 40684 20204 40736 20213
rect 41144 20204 41196 20256
rect 47032 20247 47084 20256
rect 47032 20213 47041 20247
rect 47041 20213 47075 20247
rect 47075 20213 47084 20247
rect 47032 20204 47084 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 4252 19907 4304 19916
rect 4252 19873 4261 19907
rect 4261 19873 4295 19907
rect 4295 19873 4304 19907
rect 4252 19864 4304 19873
rect 6368 19932 6420 19984
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 15016 20000 15068 20052
rect 16488 20000 16540 20052
rect 18328 20000 18380 20052
rect 18420 20000 18472 20052
rect 19892 20000 19944 20052
rect 20076 20000 20128 20052
rect 17316 19932 17368 19984
rect 5724 19864 5776 19916
rect 5448 19796 5500 19848
rect 10968 19864 11020 19916
rect 12348 19864 12400 19916
rect 13452 19864 13504 19916
rect 16304 19907 16356 19916
rect 16304 19873 16313 19907
rect 16313 19873 16347 19907
rect 16347 19873 16356 19907
rect 16304 19864 16356 19873
rect 18880 19932 18932 19984
rect 1492 19728 1544 19780
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 10784 19839 10836 19848
rect 10784 19805 10793 19839
rect 10793 19805 10827 19839
rect 10827 19805 10836 19839
rect 10784 19796 10836 19805
rect 13360 19796 13412 19848
rect 11428 19771 11480 19780
rect 11428 19737 11437 19771
rect 11437 19737 11471 19771
rect 11471 19737 11480 19771
rect 11428 19728 11480 19737
rect 11704 19728 11756 19780
rect 15200 19728 15252 19780
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 10600 19703 10652 19712
rect 10600 19669 10609 19703
rect 10609 19669 10643 19703
rect 10643 19669 10652 19703
rect 10600 19660 10652 19669
rect 10784 19660 10836 19712
rect 15476 19660 15528 19712
rect 15660 19703 15712 19712
rect 15660 19669 15669 19703
rect 15669 19669 15703 19703
rect 15703 19669 15712 19703
rect 15660 19660 15712 19669
rect 18604 19796 18656 19848
rect 19340 19864 19392 19916
rect 21456 19864 21508 19916
rect 22284 19907 22336 19916
rect 22284 19873 22293 19907
rect 22293 19873 22327 19907
rect 22327 19873 22336 19907
rect 22284 19864 22336 19873
rect 16488 19728 16540 19780
rect 17684 19728 17736 19780
rect 20720 19796 20772 19848
rect 20904 19796 20956 19848
rect 24952 20000 25004 20052
rect 25044 20000 25096 20052
rect 25228 20043 25280 20052
rect 25228 20009 25237 20043
rect 25237 20009 25271 20043
rect 25271 20009 25280 20043
rect 25228 20000 25280 20009
rect 25504 20000 25556 20052
rect 25964 20000 26016 20052
rect 26056 20000 26108 20052
rect 28540 20000 28592 20052
rect 23940 19864 23992 19916
rect 25504 19796 25556 19848
rect 27804 19932 27856 19984
rect 28632 19932 28684 19984
rect 26056 19907 26108 19916
rect 26056 19873 26065 19907
rect 26065 19873 26099 19907
rect 26099 19873 26108 19907
rect 26056 19864 26108 19873
rect 27344 19907 27396 19916
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 17316 19703 17368 19712
rect 17316 19669 17325 19703
rect 17325 19669 17359 19703
rect 17359 19669 17368 19703
rect 17316 19660 17368 19669
rect 20628 19728 20680 19780
rect 22284 19728 22336 19780
rect 19524 19660 19576 19712
rect 20444 19660 20496 19712
rect 21364 19660 21416 19712
rect 21732 19660 21784 19712
rect 25320 19728 25372 19780
rect 22652 19703 22704 19712
rect 22652 19669 22661 19703
rect 22661 19669 22695 19703
rect 22695 19669 22704 19703
rect 22652 19660 22704 19669
rect 22744 19660 22796 19712
rect 23756 19660 23808 19712
rect 24216 19660 24268 19712
rect 27344 19873 27353 19907
rect 27353 19873 27387 19907
rect 27387 19873 27396 19907
rect 27344 19864 27396 19873
rect 27528 19864 27580 19916
rect 27160 19796 27212 19848
rect 30932 20000 30984 20052
rect 31576 20000 31628 20052
rect 32772 20000 32824 20052
rect 29460 19932 29512 19984
rect 38200 20000 38252 20052
rect 38292 20000 38344 20052
rect 41052 20043 41104 20052
rect 41052 20009 41061 20043
rect 41061 20009 41095 20043
rect 41095 20009 41104 20043
rect 41052 20000 41104 20009
rect 46388 20000 46440 20052
rect 47124 20000 47176 20052
rect 29092 19864 29144 19916
rect 34704 19932 34756 19984
rect 30104 19839 30156 19848
rect 30104 19805 30113 19839
rect 30113 19805 30147 19839
rect 30147 19805 30156 19839
rect 30104 19796 30156 19805
rect 30932 19796 30984 19848
rect 31024 19796 31076 19848
rect 30380 19728 30432 19780
rect 30472 19728 30524 19780
rect 32312 19728 32364 19780
rect 26792 19703 26844 19712
rect 26792 19669 26801 19703
rect 26801 19669 26835 19703
rect 26835 19669 26844 19703
rect 26792 19660 26844 19669
rect 27160 19703 27212 19712
rect 27160 19669 27169 19703
rect 27169 19669 27203 19703
rect 27203 19669 27212 19703
rect 27160 19660 27212 19669
rect 27620 19660 27672 19712
rect 29644 19660 29696 19712
rect 29736 19703 29788 19712
rect 29736 19669 29745 19703
rect 29745 19669 29779 19703
rect 29779 19669 29788 19703
rect 29736 19660 29788 19669
rect 30012 19660 30064 19712
rect 30288 19660 30340 19712
rect 31300 19703 31352 19712
rect 31300 19669 31309 19703
rect 31309 19669 31343 19703
rect 31343 19669 31352 19703
rect 31300 19660 31352 19669
rect 32128 19703 32180 19712
rect 32128 19669 32137 19703
rect 32137 19669 32171 19703
rect 32171 19669 32180 19703
rect 32128 19660 32180 19669
rect 32772 19864 32824 19916
rect 33600 19907 33652 19916
rect 33600 19873 33609 19907
rect 33609 19873 33643 19907
rect 33643 19873 33652 19907
rect 33600 19864 33652 19873
rect 43352 19932 43404 19984
rect 44180 19932 44232 19984
rect 33784 19839 33836 19848
rect 33784 19805 33793 19839
rect 33793 19805 33827 19839
rect 33827 19805 33836 19839
rect 33784 19796 33836 19805
rect 35072 19907 35124 19916
rect 35072 19873 35081 19907
rect 35081 19873 35115 19907
rect 35115 19873 35124 19907
rect 35072 19864 35124 19873
rect 35348 19864 35400 19916
rect 36176 19864 36228 19916
rect 37372 19864 37424 19916
rect 35716 19796 35768 19848
rect 37832 19796 37884 19848
rect 39396 19864 39448 19916
rect 40316 19907 40368 19916
rect 40316 19873 40325 19907
rect 40325 19873 40359 19907
rect 40359 19873 40368 19907
rect 40316 19864 40368 19873
rect 49240 19864 49292 19916
rect 38200 19839 38252 19848
rect 38200 19805 38209 19839
rect 38209 19805 38243 19839
rect 38243 19805 38252 19839
rect 38200 19796 38252 19805
rect 39856 19796 39908 19848
rect 41052 19796 41104 19848
rect 46020 19839 46072 19848
rect 46020 19805 46029 19839
rect 46029 19805 46063 19839
rect 46063 19805 46072 19839
rect 46020 19796 46072 19805
rect 46848 19839 46900 19848
rect 46848 19805 46857 19839
rect 46857 19805 46891 19839
rect 46891 19805 46900 19839
rect 46848 19796 46900 19805
rect 34244 19728 34296 19780
rect 36360 19728 36412 19780
rect 40040 19728 40092 19780
rect 33324 19660 33376 19712
rect 33600 19660 33652 19712
rect 34336 19660 34388 19712
rect 35808 19660 35860 19712
rect 36084 19703 36136 19712
rect 36084 19669 36093 19703
rect 36093 19669 36127 19703
rect 36127 19669 36136 19703
rect 36084 19660 36136 19669
rect 36544 19703 36596 19712
rect 36544 19669 36553 19703
rect 36553 19669 36587 19703
rect 36587 19669 36596 19703
rect 36544 19660 36596 19669
rect 37556 19703 37608 19712
rect 37556 19669 37565 19703
rect 37565 19669 37599 19703
rect 37599 19669 37608 19703
rect 37556 19660 37608 19669
rect 38384 19660 38436 19712
rect 40868 19660 40920 19712
rect 46664 19660 46716 19712
rect 47584 19796 47636 19848
rect 49424 19796 49476 19848
rect 47676 19728 47728 19780
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 7564 19456 7616 19508
rect 12440 19456 12492 19508
rect 13452 19456 13504 19508
rect 3424 19388 3476 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 9220 19388 9272 19440
rect 12256 19388 12308 19440
rect 13176 19388 13228 19440
rect 15384 19499 15436 19508
rect 15384 19465 15393 19499
rect 15393 19465 15427 19499
rect 15427 19465 15436 19499
rect 15384 19456 15436 19465
rect 15476 19456 15528 19508
rect 16120 19456 16172 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 17316 19456 17368 19508
rect 19892 19456 19944 19508
rect 3884 19252 3936 19304
rect 5816 19320 5868 19372
rect 11612 19320 11664 19372
rect 6828 19252 6880 19304
rect 10416 19252 10468 19304
rect 12900 19320 12952 19372
rect 16028 19388 16080 19440
rect 16948 19388 17000 19440
rect 18328 19388 18380 19440
rect 19524 19388 19576 19440
rect 25412 19456 25464 19508
rect 25504 19456 25556 19508
rect 28264 19456 28316 19508
rect 28724 19456 28776 19508
rect 31392 19456 31444 19508
rect 32864 19456 32916 19508
rect 34244 19499 34296 19508
rect 34244 19465 34253 19499
rect 34253 19465 34287 19499
rect 34287 19465 34296 19499
rect 34244 19456 34296 19465
rect 34888 19456 34940 19508
rect 36544 19456 36596 19508
rect 36912 19456 36964 19508
rect 38476 19456 38528 19508
rect 40040 19456 40092 19508
rect 22100 19431 22152 19440
rect 22100 19397 22109 19431
rect 22109 19397 22143 19431
rect 22143 19397 22152 19431
rect 22100 19388 22152 19397
rect 22652 19388 22704 19440
rect 24492 19388 24544 19440
rect 26148 19431 26200 19440
rect 26148 19397 26157 19431
rect 26157 19397 26191 19431
rect 26191 19397 26200 19431
rect 26148 19388 26200 19397
rect 28632 19388 28684 19440
rect 15936 19320 15988 19372
rect 16672 19320 16724 19372
rect 17132 19320 17184 19372
rect 18420 19320 18472 19372
rect 7472 19184 7524 19236
rect 11980 19227 12032 19236
rect 11980 19193 11989 19227
rect 11989 19193 12023 19227
rect 12023 19193 12032 19227
rect 11980 19184 12032 19193
rect 12624 19252 12676 19304
rect 13728 19252 13780 19304
rect 14556 19252 14608 19304
rect 17040 19252 17092 19304
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 8300 19116 8352 19168
rect 11888 19116 11940 19168
rect 12808 19116 12860 19168
rect 13820 19116 13872 19168
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 15200 19184 15252 19236
rect 16120 19184 16172 19236
rect 15936 19116 15988 19168
rect 16948 19116 17000 19168
rect 23296 19320 23348 19372
rect 25688 19320 25740 19372
rect 26424 19320 26476 19372
rect 28356 19320 28408 19372
rect 31484 19431 31536 19440
rect 31484 19397 31493 19431
rect 31493 19397 31527 19431
rect 31527 19397 31536 19431
rect 31484 19388 31536 19397
rect 31760 19388 31812 19440
rect 33784 19431 33836 19440
rect 33784 19397 33793 19431
rect 33793 19397 33827 19431
rect 33827 19397 33836 19431
rect 33784 19388 33836 19397
rect 34612 19388 34664 19440
rect 34980 19388 35032 19440
rect 47584 19388 47636 19440
rect 30288 19320 30340 19372
rect 19432 19252 19484 19304
rect 19800 19295 19852 19304
rect 19800 19261 19809 19295
rect 19809 19261 19843 19295
rect 19843 19261 19852 19295
rect 19800 19252 19852 19261
rect 19616 19116 19668 19168
rect 20536 19116 20588 19168
rect 20904 19116 20956 19168
rect 24952 19295 25004 19304
rect 24952 19261 24961 19295
rect 24961 19261 24995 19295
rect 24995 19261 25004 19295
rect 24952 19252 25004 19261
rect 25596 19252 25648 19304
rect 26332 19295 26384 19304
rect 26332 19261 26341 19295
rect 26341 19261 26375 19295
rect 26375 19261 26384 19295
rect 26332 19252 26384 19261
rect 27528 19252 27580 19304
rect 27712 19295 27764 19304
rect 27712 19261 27721 19295
rect 27721 19261 27755 19295
rect 27755 19261 27764 19295
rect 27712 19252 27764 19261
rect 22284 19184 22336 19236
rect 23848 19116 23900 19168
rect 25228 19184 25280 19236
rect 26608 19184 26660 19236
rect 26792 19184 26844 19236
rect 28172 19252 28224 19304
rect 28632 19252 28684 19304
rect 28264 19184 28316 19236
rect 29368 19252 29420 19304
rect 30380 19295 30432 19304
rect 30380 19261 30389 19295
rect 30389 19261 30423 19295
rect 30423 19261 30432 19295
rect 33876 19363 33928 19372
rect 33876 19329 33885 19363
rect 33885 19329 33919 19363
rect 33919 19329 33928 19363
rect 33876 19320 33928 19329
rect 34796 19320 34848 19372
rect 30380 19252 30432 19261
rect 32312 19252 32364 19304
rect 32680 19252 32732 19304
rect 33600 19252 33652 19304
rect 34428 19252 34480 19304
rect 35900 19320 35952 19372
rect 38292 19320 38344 19372
rect 40592 19363 40644 19372
rect 40592 19329 40601 19363
rect 40601 19329 40635 19363
rect 40635 19329 40644 19363
rect 40592 19320 40644 19329
rect 47032 19320 47084 19372
rect 48412 19456 48464 19508
rect 49332 19363 49384 19372
rect 49332 19329 49341 19363
rect 49341 19329 49375 19363
rect 49375 19329 49384 19363
rect 49332 19320 49384 19329
rect 29460 19184 29512 19236
rect 29644 19184 29696 19236
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 27712 19116 27764 19168
rect 28448 19116 28500 19168
rect 29092 19116 29144 19168
rect 30288 19184 30340 19236
rect 35992 19295 36044 19304
rect 35992 19261 36001 19295
rect 36001 19261 36035 19295
rect 36035 19261 36044 19295
rect 35992 19252 36044 19261
rect 37832 19252 37884 19304
rect 39396 19295 39448 19304
rect 39396 19261 39405 19295
rect 39405 19261 39439 19295
rect 39439 19261 39448 19295
rect 39396 19252 39448 19261
rect 39672 19295 39724 19304
rect 39672 19261 39681 19295
rect 39681 19261 39715 19295
rect 39715 19261 39724 19295
rect 39672 19252 39724 19261
rect 37740 19184 37792 19236
rect 31760 19116 31812 19168
rect 32496 19116 32548 19168
rect 33416 19116 33468 19168
rect 33692 19116 33744 19168
rect 33784 19116 33836 19168
rect 36452 19116 36504 19168
rect 36636 19159 36688 19168
rect 36636 19125 36645 19159
rect 36645 19125 36679 19159
rect 36679 19125 36688 19159
rect 36636 19116 36688 19125
rect 36912 19159 36964 19168
rect 36912 19125 36921 19159
rect 36921 19125 36955 19159
rect 36955 19125 36964 19159
rect 36912 19116 36964 19125
rect 37832 19116 37884 19168
rect 39856 19184 39908 19236
rect 40500 19116 40552 19168
rect 42064 19116 42116 19168
rect 46664 19159 46716 19168
rect 46664 19125 46673 19159
rect 46673 19125 46707 19159
rect 46707 19125 46716 19159
rect 46664 19116 46716 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 6828 18912 6880 18964
rect 11152 18912 11204 18964
rect 11520 18912 11572 18964
rect 13636 18955 13688 18964
rect 13636 18921 13645 18955
rect 13645 18921 13679 18955
rect 13679 18921 13688 18955
rect 13636 18912 13688 18921
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 3792 18776 3844 18828
rect 11244 18844 11296 18896
rect 11888 18887 11940 18896
rect 11888 18853 11897 18887
rect 11897 18853 11931 18887
rect 11931 18853 11940 18887
rect 11888 18844 11940 18853
rect 13360 18844 13412 18896
rect 1400 18640 1452 18692
rect 7748 18708 7800 18760
rect 12440 18776 12492 18828
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 14556 18776 14608 18828
rect 15016 18776 15068 18828
rect 4344 18640 4396 18692
rect 10232 18640 10284 18692
rect 7380 18572 7432 18624
rect 10692 18683 10744 18692
rect 10692 18649 10701 18683
rect 10701 18649 10735 18683
rect 10735 18649 10744 18683
rect 10692 18640 10744 18649
rect 12256 18708 12308 18760
rect 12440 18640 12492 18692
rect 15660 18708 15712 18760
rect 15936 18912 15988 18964
rect 16120 18912 16172 18964
rect 16488 18912 16540 18964
rect 19892 18955 19944 18964
rect 19892 18921 19901 18955
rect 19901 18921 19935 18955
rect 19935 18921 19944 18955
rect 19892 18912 19944 18921
rect 16764 18844 16816 18896
rect 16580 18776 16632 18828
rect 19708 18776 19760 18828
rect 20720 18844 20772 18896
rect 20444 18819 20496 18828
rect 20444 18785 20453 18819
rect 20453 18785 20487 18819
rect 20487 18785 20496 18819
rect 20444 18776 20496 18785
rect 21180 18776 21232 18828
rect 22284 18955 22336 18964
rect 22284 18921 22293 18955
rect 22293 18921 22327 18955
rect 22327 18921 22336 18955
rect 22284 18912 22336 18921
rect 22744 18912 22796 18964
rect 27620 18912 27672 18964
rect 27712 18912 27764 18964
rect 30012 18912 30064 18964
rect 30932 18955 30984 18964
rect 30932 18921 30941 18955
rect 30941 18921 30975 18955
rect 30975 18921 30984 18955
rect 30932 18912 30984 18921
rect 32956 18912 33008 18964
rect 34980 18912 35032 18964
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 25688 18776 25740 18828
rect 27068 18844 27120 18896
rect 26700 18776 26752 18828
rect 28448 18776 28500 18828
rect 28908 18776 28960 18828
rect 11980 18572 12032 18624
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 14556 18640 14608 18649
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 20904 18708 20956 18760
rect 22284 18708 22336 18760
rect 24124 18708 24176 18760
rect 27436 18708 27488 18760
rect 28172 18751 28224 18760
rect 28172 18717 28181 18751
rect 28181 18717 28215 18751
rect 28215 18717 28224 18751
rect 29644 18776 29696 18828
rect 29920 18819 29972 18828
rect 29920 18785 29929 18819
rect 29929 18785 29963 18819
rect 29963 18785 29972 18819
rect 29920 18776 29972 18785
rect 32680 18844 32732 18896
rect 33232 18844 33284 18896
rect 33692 18844 33744 18896
rect 39396 18912 39448 18964
rect 41512 18912 41564 18964
rect 42064 18955 42116 18964
rect 42064 18921 42073 18955
rect 42073 18921 42107 18955
rect 42107 18921 42116 18955
rect 42064 18912 42116 18921
rect 47492 18912 47544 18964
rect 41880 18844 41932 18896
rect 34152 18819 34204 18828
rect 28172 18708 28224 18717
rect 19340 18640 19392 18692
rect 19616 18640 19668 18692
rect 15568 18572 15620 18624
rect 15844 18572 15896 18624
rect 17408 18615 17460 18624
rect 17408 18581 17417 18615
rect 17417 18581 17451 18615
rect 17451 18581 17460 18615
rect 17408 18572 17460 18581
rect 17500 18572 17552 18624
rect 21364 18572 21416 18624
rect 21640 18572 21692 18624
rect 23480 18640 23532 18692
rect 23848 18640 23900 18692
rect 26148 18640 26200 18692
rect 24768 18572 24820 18624
rect 25044 18615 25096 18624
rect 25044 18581 25053 18615
rect 25053 18581 25087 18615
rect 25087 18581 25096 18615
rect 25044 18572 25096 18581
rect 25136 18572 25188 18624
rect 29368 18640 29420 18692
rect 29828 18640 29880 18692
rect 30748 18683 30800 18692
rect 28356 18615 28408 18624
rect 28356 18581 28365 18615
rect 28365 18581 28399 18615
rect 28399 18581 28408 18615
rect 28356 18572 28408 18581
rect 28632 18615 28684 18624
rect 28632 18581 28641 18615
rect 28641 18581 28675 18615
rect 28675 18581 28684 18615
rect 28632 18572 28684 18581
rect 29184 18572 29236 18624
rect 29644 18572 29696 18624
rect 30748 18649 30757 18683
rect 30757 18649 30791 18683
rect 30791 18649 30800 18683
rect 30748 18640 30800 18649
rect 30472 18615 30524 18624
rect 30472 18581 30481 18615
rect 30481 18581 30515 18615
rect 30515 18581 30524 18615
rect 30472 18572 30524 18581
rect 31024 18572 31076 18624
rect 31300 18572 31352 18624
rect 31852 18615 31904 18624
rect 31852 18581 31861 18615
rect 31861 18581 31895 18615
rect 31895 18581 31904 18615
rect 31852 18572 31904 18581
rect 32680 18708 32732 18760
rect 34152 18785 34161 18819
rect 34161 18785 34195 18819
rect 34195 18785 34204 18819
rect 34152 18776 34204 18785
rect 34520 18776 34572 18828
rect 37280 18776 37332 18828
rect 33508 18708 33560 18760
rect 33876 18708 33928 18760
rect 34612 18708 34664 18760
rect 35532 18708 35584 18760
rect 35348 18640 35400 18692
rect 32772 18572 32824 18624
rect 32956 18572 33008 18624
rect 33784 18572 33836 18624
rect 33876 18615 33928 18624
rect 33876 18581 33885 18615
rect 33885 18581 33919 18615
rect 33919 18581 33928 18615
rect 33876 18572 33928 18581
rect 36084 18572 36136 18624
rect 36820 18572 36872 18624
rect 38568 18819 38620 18828
rect 38568 18785 38577 18819
rect 38577 18785 38611 18819
rect 38611 18785 38620 18819
rect 38568 18776 38620 18785
rect 39672 18776 39724 18828
rect 48412 18776 48464 18828
rect 37556 18572 37608 18624
rect 39672 18640 39724 18692
rect 38016 18615 38068 18624
rect 38016 18581 38025 18615
rect 38025 18581 38059 18615
rect 38059 18581 38068 18615
rect 38016 18572 38068 18581
rect 38476 18615 38528 18624
rect 38476 18581 38485 18615
rect 38485 18581 38519 18615
rect 38519 18581 38528 18615
rect 38476 18572 38528 18581
rect 40132 18572 40184 18624
rect 40500 18640 40552 18692
rect 49424 18708 49476 18760
rect 47308 18615 47360 18624
rect 47308 18581 47317 18615
rect 47317 18581 47351 18615
rect 47351 18581 47360 18615
rect 47308 18572 47360 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 9864 18368 9916 18420
rect 10416 18368 10468 18420
rect 12440 18368 12492 18420
rect 25780 18368 25832 18420
rect 27252 18368 27304 18420
rect 27712 18368 27764 18420
rect 30196 18368 30248 18420
rect 31208 18368 31260 18420
rect 32588 18411 32640 18420
rect 32588 18377 32597 18411
rect 32597 18377 32631 18411
rect 32631 18377 32640 18411
rect 32588 18368 32640 18377
rect 32772 18368 32824 18420
rect 4528 18300 4580 18352
rect 7656 18343 7708 18352
rect 7656 18309 7665 18343
rect 7665 18309 7699 18343
rect 7699 18309 7708 18343
rect 7656 18300 7708 18309
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 4068 18232 4120 18284
rect 11428 18300 11480 18352
rect 13084 18300 13136 18352
rect 13544 18300 13596 18352
rect 16764 18300 16816 18352
rect 16948 18343 17000 18352
rect 16948 18309 16957 18343
rect 16957 18309 16991 18343
rect 16991 18309 17000 18343
rect 16948 18300 17000 18309
rect 4252 18164 4304 18216
rect 11888 18232 11940 18284
rect 10600 18164 10652 18216
rect 11704 18164 11756 18216
rect 11980 18164 12032 18216
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 15016 18232 15068 18284
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 17040 18232 17092 18284
rect 14556 18207 14608 18216
rect 14556 18173 14565 18207
rect 14565 18173 14599 18207
rect 14599 18173 14608 18207
rect 14556 18164 14608 18173
rect 14924 18207 14976 18216
rect 14924 18173 14933 18207
rect 14933 18173 14967 18207
rect 14967 18173 14976 18207
rect 14924 18164 14976 18173
rect 9680 18028 9732 18080
rect 9772 18028 9824 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 13728 18096 13780 18148
rect 15936 18096 15988 18148
rect 17500 18300 17552 18352
rect 16672 18096 16724 18148
rect 18512 18232 18564 18284
rect 19156 18300 19208 18352
rect 20628 18300 20680 18352
rect 22652 18300 22704 18352
rect 21272 18232 21324 18284
rect 19616 18207 19668 18216
rect 19616 18173 19625 18207
rect 19625 18173 19659 18207
rect 19659 18173 19668 18207
rect 19616 18164 19668 18173
rect 22744 18232 22796 18284
rect 24124 18343 24176 18352
rect 24124 18309 24133 18343
rect 24133 18309 24167 18343
rect 24167 18309 24176 18343
rect 24124 18300 24176 18309
rect 24492 18300 24544 18352
rect 23388 18232 23440 18284
rect 24676 18232 24728 18284
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 32128 18300 32180 18352
rect 33232 18300 33284 18352
rect 33968 18300 34020 18352
rect 35348 18411 35400 18420
rect 35348 18377 35357 18411
rect 35357 18377 35391 18411
rect 35391 18377 35400 18411
rect 35348 18368 35400 18377
rect 37188 18368 37240 18420
rect 40868 18411 40920 18420
rect 40868 18377 40877 18411
rect 40877 18377 40911 18411
rect 40911 18377 40920 18411
rect 40868 18368 40920 18377
rect 48412 18368 48464 18420
rect 36084 18300 36136 18352
rect 26700 18164 26752 18216
rect 13544 18028 13596 18080
rect 15292 18028 15344 18080
rect 18604 18028 18656 18080
rect 23664 18096 23716 18148
rect 21180 18028 21232 18080
rect 21456 18028 21508 18080
rect 22468 18028 22520 18080
rect 25044 18028 25096 18080
rect 26056 18096 26108 18148
rect 30104 18232 30156 18284
rect 28908 18207 28960 18216
rect 28908 18173 28917 18207
rect 28917 18173 28951 18207
rect 28951 18173 28960 18207
rect 28908 18164 28960 18173
rect 32036 18232 32088 18284
rect 33140 18232 33192 18284
rect 35256 18232 35308 18284
rect 36268 18275 36320 18284
rect 36268 18241 36277 18275
rect 36277 18241 36311 18275
rect 36311 18241 36320 18275
rect 36268 18232 36320 18241
rect 36912 18232 36964 18284
rect 37280 18300 37332 18352
rect 38016 18300 38068 18352
rect 47308 18300 47360 18352
rect 38384 18232 38436 18284
rect 39764 18275 39816 18284
rect 39764 18241 39773 18275
rect 39773 18241 39807 18275
rect 39807 18241 39816 18275
rect 39764 18232 39816 18241
rect 49332 18275 49384 18284
rect 49332 18241 49341 18275
rect 49341 18241 49375 18275
rect 49375 18241 49384 18275
rect 49332 18232 49384 18241
rect 29000 18096 29052 18148
rect 29276 18096 29328 18148
rect 26332 18028 26384 18080
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 28264 18028 28316 18080
rect 28908 18028 28960 18080
rect 29644 18028 29696 18080
rect 30288 18207 30340 18216
rect 30288 18173 30297 18207
rect 30297 18173 30331 18207
rect 30331 18173 30340 18207
rect 30288 18164 30340 18173
rect 32496 18207 32548 18216
rect 32496 18173 32505 18207
rect 32505 18173 32539 18207
rect 32539 18173 32548 18207
rect 32496 18164 32548 18173
rect 33600 18207 33652 18216
rect 33600 18173 33609 18207
rect 33609 18173 33643 18207
rect 33643 18173 33652 18207
rect 33600 18164 33652 18173
rect 33876 18207 33928 18216
rect 33876 18173 33885 18207
rect 33885 18173 33919 18207
rect 33919 18173 33928 18207
rect 33876 18164 33928 18173
rect 37740 18164 37792 18216
rect 37832 18164 37884 18216
rect 30012 18096 30064 18148
rect 33416 18096 33468 18148
rect 37004 18139 37056 18148
rect 37004 18105 37013 18139
rect 37013 18105 37047 18139
rect 37047 18105 37056 18139
rect 37004 18096 37056 18105
rect 37556 18096 37608 18148
rect 38016 18139 38068 18148
rect 38016 18105 38025 18139
rect 38025 18105 38059 18139
rect 38059 18105 38068 18139
rect 38016 18096 38068 18105
rect 30748 18028 30800 18080
rect 32956 18028 33008 18080
rect 35900 18028 35952 18080
rect 36728 18028 36780 18080
rect 40040 18071 40092 18080
rect 40040 18037 40049 18071
rect 40049 18037 40083 18071
rect 40083 18037 40092 18071
rect 40040 18028 40092 18037
rect 40500 18028 40552 18080
rect 48044 18071 48096 18080
rect 48044 18037 48053 18071
rect 48053 18037 48087 18071
rect 48087 18037 48096 18071
rect 48044 18028 48096 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 10232 17824 10284 17876
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 3332 17756 3384 17808
rect 12440 17824 12492 17876
rect 12532 17824 12584 17876
rect 14556 17824 14608 17876
rect 15108 17824 15160 17876
rect 16580 17824 16632 17876
rect 17224 17824 17276 17876
rect 19432 17867 19484 17876
rect 19432 17833 19441 17867
rect 19441 17833 19475 17867
rect 19475 17833 19484 17867
rect 19432 17824 19484 17833
rect 19616 17824 19668 17876
rect 21088 17824 21140 17876
rect 21180 17824 21232 17876
rect 12532 17688 12584 17740
rect 13452 17688 13504 17740
rect 19524 17756 19576 17808
rect 10416 17620 10468 17672
rect 16028 17731 16080 17740
rect 16028 17697 16037 17731
rect 16037 17697 16071 17731
rect 16071 17697 16080 17731
rect 16028 17688 16080 17697
rect 16396 17688 16448 17740
rect 17316 17688 17368 17740
rect 23296 17867 23348 17876
rect 23296 17833 23305 17867
rect 23305 17833 23339 17867
rect 23339 17833 23348 17867
rect 23296 17824 23348 17833
rect 23572 17824 23624 17876
rect 1032 17552 1084 17604
rect 10324 17527 10376 17536
rect 10324 17493 10333 17527
rect 10333 17493 10367 17527
rect 10367 17493 10376 17527
rect 10324 17484 10376 17493
rect 11796 17552 11848 17604
rect 12072 17595 12124 17604
rect 12072 17561 12081 17595
rect 12081 17561 12115 17595
rect 12115 17561 12124 17595
rect 12072 17552 12124 17561
rect 16672 17620 16724 17672
rect 17776 17620 17828 17672
rect 18420 17620 18472 17672
rect 14004 17552 14056 17604
rect 15016 17552 15068 17604
rect 16028 17552 16080 17604
rect 17500 17552 17552 17604
rect 18604 17552 18656 17604
rect 20352 17620 20404 17672
rect 21640 17688 21692 17740
rect 21732 17731 21784 17740
rect 21732 17697 21741 17731
rect 21741 17697 21775 17731
rect 21775 17697 21784 17731
rect 21732 17688 21784 17697
rect 22100 17688 22152 17740
rect 23756 17731 23808 17740
rect 23756 17697 23765 17731
rect 23765 17697 23799 17731
rect 23799 17697 23808 17731
rect 23756 17688 23808 17697
rect 24952 17688 25004 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 23480 17620 23532 17672
rect 29276 17824 29328 17876
rect 29552 17867 29604 17876
rect 29552 17833 29561 17867
rect 29561 17833 29595 17867
rect 29595 17833 29604 17867
rect 29552 17824 29604 17833
rect 33416 17824 33468 17876
rect 35532 17824 35584 17876
rect 36176 17824 36228 17876
rect 37648 17824 37700 17876
rect 38476 17824 38528 17876
rect 28908 17756 28960 17808
rect 29184 17756 29236 17808
rect 26148 17688 26200 17740
rect 32680 17756 32732 17808
rect 31484 17731 31536 17740
rect 31484 17697 31493 17731
rect 31493 17697 31527 17731
rect 31527 17697 31536 17731
rect 31484 17688 31536 17697
rect 35072 17756 35124 17808
rect 35256 17756 35308 17808
rect 33324 17688 33376 17740
rect 26240 17663 26292 17672
rect 26240 17629 26249 17663
rect 26249 17629 26283 17663
rect 26283 17629 26292 17663
rect 26240 17620 26292 17629
rect 27436 17620 27488 17672
rect 28908 17620 28960 17672
rect 31392 17620 31444 17672
rect 31760 17620 31812 17672
rect 37648 17688 37700 17740
rect 36176 17620 36228 17672
rect 37556 17663 37608 17672
rect 37556 17629 37565 17663
rect 37565 17629 37599 17663
rect 37599 17629 37608 17663
rect 37556 17620 37608 17629
rect 46940 17756 46992 17808
rect 40684 17688 40736 17740
rect 20720 17552 20772 17604
rect 21640 17552 21692 17604
rect 11980 17484 12032 17536
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 16488 17527 16540 17536
rect 16488 17493 16497 17527
rect 16497 17493 16531 17527
rect 16531 17493 16540 17527
rect 16488 17484 16540 17493
rect 18788 17484 18840 17536
rect 22560 17484 22612 17536
rect 25136 17552 25188 17604
rect 25228 17552 25280 17604
rect 28448 17552 28500 17604
rect 29184 17552 29236 17604
rect 30104 17552 30156 17604
rect 30380 17552 30432 17604
rect 31668 17595 31720 17604
rect 31668 17561 31677 17595
rect 31677 17561 31711 17595
rect 31711 17561 31720 17595
rect 31668 17552 31720 17561
rect 24676 17484 24728 17536
rect 25044 17484 25096 17536
rect 26608 17484 26660 17536
rect 27068 17527 27120 17536
rect 27068 17493 27077 17527
rect 27077 17493 27111 17527
rect 27111 17493 27120 17527
rect 27068 17484 27120 17493
rect 28264 17484 28316 17536
rect 29092 17527 29144 17536
rect 29092 17493 29101 17527
rect 29101 17493 29135 17527
rect 29135 17493 29144 17527
rect 29092 17484 29144 17493
rect 32404 17552 32456 17604
rect 32128 17484 32180 17536
rect 33416 17484 33468 17536
rect 33692 17484 33744 17536
rect 34428 17484 34480 17536
rect 35072 17527 35124 17536
rect 35072 17493 35081 17527
rect 35081 17493 35115 17527
rect 35115 17493 35124 17527
rect 35072 17484 35124 17493
rect 35440 17527 35492 17536
rect 35440 17493 35449 17527
rect 35449 17493 35483 17527
rect 35483 17493 35492 17527
rect 35440 17484 35492 17493
rect 35532 17484 35584 17536
rect 36636 17484 36688 17536
rect 38384 17527 38436 17536
rect 38384 17493 38393 17527
rect 38393 17493 38427 17527
rect 38427 17493 38436 17527
rect 38384 17484 38436 17493
rect 40592 17552 40644 17604
rect 38936 17484 38988 17536
rect 39120 17484 39172 17536
rect 40040 17484 40092 17536
rect 40776 17620 40828 17672
rect 49332 17663 49384 17672
rect 49332 17629 49341 17663
rect 49341 17629 49375 17663
rect 49375 17629 49384 17663
rect 49332 17620 49384 17629
rect 47032 17552 47084 17604
rect 43444 17484 43496 17536
rect 47676 17527 47728 17536
rect 47676 17493 47685 17527
rect 47685 17493 47719 17527
rect 47719 17493 47728 17527
rect 47676 17484 47728 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 7380 17280 7432 17332
rect 12440 17280 12492 17332
rect 17040 17280 17092 17332
rect 19156 17323 19208 17332
rect 19156 17289 19165 17323
rect 19165 17289 19199 17323
rect 19199 17289 19208 17323
rect 19156 17280 19208 17289
rect 10324 17212 10376 17264
rect 4344 17144 4396 17196
rect 5816 17144 5868 17196
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 9956 17144 10008 17196
rect 11980 17212 12032 17264
rect 13636 17212 13688 17264
rect 14280 17255 14332 17264
rect 14280 17221 14289 17255
rect 14289 17221 14323 17255
rect 14323 17221 14332 17255
rect 14280 17212 14332 17221
rect 16396 17212 16448 17264
rect 18880 17212 18932 17264
rect 18972 17212 19024 17264
rect 22560 17280 22612 17332
rect 23480 17280 23532 17332
rect 24860 17323 24912 17332
rect 24860 17289 24869 17323
rect 24869 17289 24903 17323
rect 24903 17289 24912 17323
rect 24860 17280 24912 17289
rect 27804 17280 27856 17332
rect 20536 17212 20588 17264
rect 21272 17212 21324 17264
rect 21548 17212 21600 17264
rect 21732 17212 21784 17264
rect 22100 17212 22152 17264
rect 22744 17212 22796 17264
rect 24124 17212 24176 17264
rect 14188 17144 14240 17196
rect 940 17076 992 17128
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 5448 17008 5500 17060
rect 10600 17076 10652 17128
rect 12348 17076 12400 17128
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 15384 17144 15436 17196
rect 11796 17008 11848 17060
rect 13912 17008 13964 17060
rect 15568 17051 15620 17060
rect 15568 17017 15577 17051
rect 15577 17017 15611 17051
rect 15611 17017 15620 17051
rect 15568 17008 15620 17017
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 18604 17144 18656 17196
rect 19064 17144 19116 17196
rect 25964 17255 26016 17264
rect 25964 17221 25973 17255
rect 25973 17221 26007 17255
rect 26007 17221 26016 17255
rect 25964 17212 26016 17221
rect 26884 17212 26936 17264
rect 19892 17076 19944 17128
rect 16488 17008 16540 17060
rect 12256 16940 12308 16992
rect 13360 16940 13412 16992
rect 13728 16983 13780 16992
rect 13728 16949 13737 16983
rect 13737 16949 13771 16983
rect 13771 16949 13780 16983
rect 13728 16940 13780 16949
rect 15844 16940 15896 16992
rect 15936 16940 15988 16992
rect 21640 17051 21692 17060
rect 21640 17017 21649 17051
rect 21649 17017 21683 17051
rect 21683 17017 21692 17051
rect 21640 17008 21692 17017
rect 22284 17008 22336 17060
rect 25596 17144 25648 17196
rect 27620 17144 27672 17196
rect 24492 17076 24544 17128
rect 25504 17119 25556 17128
rect 25504 17085 25513 17119
rect 25513 17085 25547 17119
rect 25547 17085 25556 17119
rect 25504 17076 25556 17085
rect 26976 17076 27028 17128
rect 27988 17144 28040 17196
rect 29552 17212 29604 17264
rect 30656 17280 30708 17332
rect 31392 17280 31444 17332
rect 32036 17212 32088 17264
rect 27896 17119 27948 17128
rect 27896 17085 27905 17119
rect 27905 17085 27939 17119
rect 27939 17085 27948 17119
rect 27896 17076 27948 17085
rect 27252 17008 27304 17060
rect 22376 16940 22428 16992
rect 29736 17076 29788 17128
rect 30564 17144 30616 17196
rect 30104 17119 30156 17128
rect 30104 17085 30113 17119
rect 30113 17085 30147 17119
rect 30147 17085 30156 17119
rect 30104 17076 30156 17085
rect 30380 17076 30432 17128
rect 30288 17008 30340 17060
rect 30748 17076 30800 17128
rect 32220 17144 32272 17196
rect 33600 17280 33652 17332
rect 35072 17280 35124 17332
rect 38476 17323 38528 17332
rect 38476 17289 38485 17323
rect 38485 17289 38519 17323
rect 38519 17289 38528 17323
rect 38476 17280 38528 17289
rect 38660 17280 38712 17332
rect 40040 17280 40092 17332
rect 41052 17280 41104 17332
rect 47032 17323 47084 17332
rect 47032 17289 47041 17323
rect 47041 17289 47075 17323
rect 47075 17289 47084 17323
rect 47032 17280 47084 17289
rect 34428 17212 34480 17264
rect 35440 17212 35492 17264
rect 39120 17212 39172 17264
rect 40132 17212 40184 17264
rect 47676 17212 47728 17264
rect 48228 17212 48280 17264
rect 35164 17144 35216 17196
rect 36360 17187 36412 17196
rect 36360 17153 36369 17187
rect 36369 17153 36403 17187
rect 36403 17153 36412 17187
rect 36360 17144 36412 17153
rect 38936 17144 38988 17196
rect 32588 17119 32640 17128
rect 32588 17085 32597 17119
rect 32597 17085 32631 17119
rect 32631 17085 32640 17119
rect 32588 17076 32640 17085
rect 32680 17076 32732 17128
rect 34796 17119 34848 17128
rect 34796 17085 34805 17119
rect 34805 17085 34839 17119
rect 34839 17085 34848 17119
rect 34796 17076 34848 17085
rect 36544 17076 36596 17128
rect 37832 17076 37884 17128
rect 31576 17008 31628 17060
rect 33876 17008 33928 17060
rect 40684 17119 40736 17128
rect 40684 17085 40693 17119
rect 40693 17085 40727 17119
rect 40727 17085 40736 17119
rect 40684 17076 40736 17085
rect 30196 16940 30248 16992
rect 31760 16983 31812 16992
rect 31760 16949 31769 16983
rect 31769 16949 31803 16983
rect 31803 16949 31812 16983
rect 31760 16940 31812 16949
rect 35348 16940 35400 16992
rect 36636 16940 36688 16992
rect 37280 16940 37332 16992
rect 37464 16983 37516 16992
rect 37464 16949 37473 16983
rect 37473 16949 37507 16983
rect 37507 16949 37516 16983
rect 37464 16940 37516 16949
rect 38844 16940 38896 16992
rect 40776 16940 40828 16992
rect 41696 16940 41748 16992
rect 47952 17119 48004 17128
rect 47952 17085 47961 17119
rect 47961 17085 47995 17119
rect 47995 17085 48004 17119
rect 47952 17076 48004 17085
rect 48320 16940 48372 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 9864 16668 9916 16720
rect 11980 16736 12032 16788
rect 12256 16736 12308 16788
rect 13728 16736 13780 16788
rect 13912 16736 13964 16788
rect 14924 16736 14976 16788
rect 16212 16736 16264 16788
rect 18972 16736 19024 16788
rect 19064 16736 19116 16788
rect 23388 16736 23440 16788
rect 26332 16736 26384 16788
rect 27620 16736 27672 16788
rect 28540 16736 28592 16788
rect 28724 16736 28776 16788
rect 29368 16779 29420 16788
rect 29368 16745 29377 16779
rect 29377 16745 29411 16779
rect 29411 16745 29420 16779
rect 29368 16736 29420 16745
rect 30104 16736 30156 16788
rect 10600 16668 10652 16720
rect 4436 16600 4488 16652
rect 3332 16532 3384 16584
rect 1032 16464 1084 16516
rect 9036 16600 9088 16652
rect 9496 16600 9548 16652
rect 10508 16600 10560 16652
rect 11152 16643 11204 16652
rect 11152 16609 11161 16643
rect 11161 16609 11195 16643
rect 11195 16609 11204 16643
rect 11152 16600 11204 16609
rect 11796 16600 11848 16652
rect 12624 16600 12676 16652
rect 7564 16532 7616 16584
rect 11980 16532 12032 16584
rect 12164 16532 12216 16584
rect 12256 16532 12308 16584
rect 14740 16668 14792 16720
rect 13912 16600 13964 16652
rect 14188 16643 14240 16652
rect 14188 16609 14197 16643
rect 14197 16609 14231 16643
rect 14231 16609 14240 16643
rect 14188 16600 14240 16609
rect 15844 16600 15896 16652
rect 16948 16668 17000 16720
rect 17500 16668 17552 16720
rect 20996 16711 21048 16720
rect 20996 16677 21005 16711
rect 21005 16677 21039 16711
rect 21039 16677 21048 16711
rect 20996 16668 21048 16677
rect 21272 16668 21324 16720
rect 13820 16532 13872 16584
rect 15752 16532 15804 16584
rect 18236 16600 18288 16652
rect 18604 16643 18656 16652
rect 18604 16609 18613 16643
rect 18613 16609 18647 16643
rect 18647 16609 18656 16643
rect 18604 16600 18656 16609
rect 18880 16643 18932 16652
rect 18880 16609 18889 16643
rect 18889 16609 18923 16643
rect 18923 16609 18932 16643
rect 18880 16600 18932 16609
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 26056 16668 26108 16720
rect 27988 16668 28040 16720
rect 25872 16600 25924 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27436 16600 27488 16652
rect 29460 16600 29512 16652
rect 30012 16643 30064 16652
rect 30012 16609 30021 16643
rect 30021 16609 30055 16643
rect 30055 16609 30064 16643
rect 30012 16600 30064 16609
rect 17500 16532 17552 16584
rect 9680 16464 9732 16516
rect 10508 16507 10560 16516
rect 10508 16473 10517 16507
rect 10517 16473 10551 16507
rect 10551 16473 10560 16507
rect 10508 16464 10560 16473
rect 12808 16464 12860 16516
rect 14648 16464 14700 16516
rect 20720 16532 20772 16584
rect 24584 16575 24636 16584
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 11336 16439 11388 16448
rect 11336 16405 11345 16439
rect 11345 16405 11379 16439
rect 11379 16405 11388 16439
rect 11336 16396 11388 16405
rect 12164 16396 12216 16448
rect 12716 16396 12768 16448
rect 13452 16396 13504 16448
rect 14924 16396 14976 16448
rect 15476 16396 15528 16448
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 16212 16396 16264 16448
rect 17132 16439 17184 16448
rect 17132 16405 17141 16439
rect 17141 16405 17175 16439
rect 17175 16405 17184 16439
rect 17132 16396 17184 16405
rect 28908 16532 28960 16584
rect 29000 16532 29052 16584
rect 18328 16396 18380 16448
rect 18972 16396 19024 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 20720 16396 20772 16448
rect 28448 16507 28500 16516
rect 28448 16473 28457 16507
rect 28457 16473 28491 16507
rect 28491 16473 28500 16507
rect 33876 16736 33928 16788
rect 34428 16736 34480 16788
rect 36176 16736 36228 16788
rect 36360 16736 36412 16788
rect 36636 16736 36688 16788
rect 30564 16668 30616 16720
rect 31116 16643 31168 16652
rect 31116 16609 31125 16643
rect 31125 16609 31159 16643
rect 31159 16609 31168 16643
rect 31116 16600 31168 16609
rect 28448 16464 28500 16473
rect 22836 16396 22888 16448
rect 23296 16439 23348 16448
rect 23296 16405 23305 16439
rect 23305 16405 23339 16439
rect 23339 16405 23348 16439
rect 23296 16396 23348 16405
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 27528 16396 27580 16448
rect 28172 16396 28224 16448
rect 29368 16396 29420 16448
rect 31024 16532 31076 16584
rect 32220 16643 32272 16652
rect 32220 16609 32229 16643
rect 32229 16609 32263 16643
rect 32263 16609 32272 16643
rect 32220 16600 32272 16609
rect 32496 16643 32548 16652
rect 32496 16609 32505 16643
rect 32505 16609 32539 16643
rect 32539 16609 32548 16643
rect 32496 16600 32548 16609
rect 37556 16668 37608 16720
rect 37096 16600 37148 16652
rect 40224 16736 40276 16788
rect 41052 16779 41104 16788
rect 41052 16745 41061 16779
rect 41061 16745 41095 16779
rect 41095 16745 41104 16779
rect 41052 16736 41104 16745
rect 41236 16779 41288 16788
rect 41236 16745 41245 16779
rect 41245 16745 41279 16779
rect 41279 16745 41288 16779
rect 41236 16736 41288 16745
rect 48780 16668 48832 16720
rect 38844 16600 38896 16652
rect 40316 16600 40368 16652
rect 41052 16600 41104 16652
rect 31944 16532 31996 16584
rect 34428 16532 34480 16584
rect 35440 16532 35492 16584
rect 36636 16532 36688 16584
rect 39488 16575 39540 16584
rect 39488 16541 39497 16575
rect 39497 16541 39531 16575
rect 39531 16541 39540 16575
rect 39488 16532 39540 16541
rect 40684 16532 40736 16584
rect 32128 16464 32180 16516
rect 35900 16464 35952 16516
rect 38660 16464 38712 16516
rect 40224 16464 40276 16516
rect 41236 16464 41288 16516
rect 31300 16439 31352 16448
rect 31300 16405 31309 16439
rect 31309 16405 31343 16439
rect 31343 16405 31352 16439
rect 31300 16396 31352 16405
rect 31852 16396 31904 16448
rect 33968 16439 34020 16448
rect 33968 16405 33977 16439
rect 33977 16405 34011 16439
rect 34011 16405 34020 16439
rect 33968 16396 34020 16405
rect 34336 16439 34388 16448
rect 34336 16405 34345 16439
rect 34345 16405 34379 16439
rect 34379 16405 34388 16439
rect 34336 16396 34388 16405
rect 35532 16396 35584 16448
rect 36728 16396 36780 16448
rect 38568 16396 38620 16448
rect 40960 16396 41012 16448
rect 49332 16575 49384 16584
rect 49332 16541 49341 16575
rect 49341 16541 49375 16575
rect 49375 16541 49384 16575
rect 49332 16532 49384 16541
rect 41604 16396 41656 16448
rect 47860 16396 47912 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 9772 16192 9824 16244
rect 11060 16192 11112 16244
rect 11336 16192 11388 16244
rect 10876 16124 10928 16176
rect 15936 16192 15988 16244
rect 17408 16235 17460 16244
rect 17408 16201 17417 16235
rect 17417 16201 17451 16235
rect 17451 16201 17460 16235
rect 17408 16192 17460 16201
rect 18328 16192 18380 16244
rect 18604 16192 18656 16244
rect 23296 16192 23348 16244
rect 4252 16056 4304 16108
rect 11060 16099 11112 16108
rect 1032 15988 1084 16040
rect 9036 15988 9088 16040
rect 11060 16065 11069 16099
rect 11069 16065 11103 16099
rect 11103 16065 11112 16099
rect 11060 16056 11112 16065
rect 13912 16056 13964 16108
rect 9772 15920 9824 15972
rect 9864 15852 9916 15904
rect 10600 15852 10652 15904
rect 10784 15920 10836 15972
rect 12440 15988 12492 16040
rect 13452 15988 13504 16040
rect 13544 15988 13596 16040
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 17132 16124 17184 16176
rect 14740 16056 14792 16108
rect 11520 15852 11572 15904
rect 14280 15920 14332 15972
rect 14648 15988 14700 16040
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 15752 16031 15804 16040
rect 15752 15997 15761 16031
rect 15761 15997 15795 16031
rect 15795 15997 15804 16031
rect 15752 15988 15804 15997
rect 14464 15920 14516 15972
rect 16856 16056 16908 16108
rect 17408 16056 17460 16108
rect 17224 15988 17276 16040
rect 20720 16124 20772 16176
rect 21640 16124 21692 16176
rect 18880 16056 18932 16108
rect 24584 16124 24636 16176
rect 17592 15920 17644 15972
rect 19984 15988 20036 16040
rect 16488 15852 16540 15904
rect 16948 15852 17000 15904
rect 17316 15852 17368 15904
rect 19064 15920 19116 15972
rect 18420 15852 18472 15904
rect 18788 15852 18840 15904
rect 19156 15852 19208 15904
rect 23572 16056 23624 16108
rect 27804 16124 27856 16176
rect 26608 16056 26660 16108
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 28264 16056 28316 16108
rect 28908 16124 28960 16176
rect 29092 16124 29144 16176
rect 30380 16192 30432 16244
rect 31760 16192 31812 16244
rect 34796 16192 34848 16244
rect 30656 16124 30708 16176
rect 30840 16167 30892 16176
rect 30840 16133 30849 16167
rect 30849 16133 30883 16167
rect 30883 16133 30892 16167
rect 30840 16124 30892 16133
rect 20812 15988 20864 16040
rect 21916 15988 21968 16040
rect 20720 15920 20772 15972
rect 22192 15920 22244 15972
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 21640 15852 21692 15904
rect 23480 15920 23532 15972
rect 24492 15988 24544 16040
rect 26792 15988 26844 16040
rect 24676 15920 24728 15972
rect 27436 15988 27488 16040
rect 26976 15920 27028 15972
rect 28632 16031 28684 16040
rect 28632 15997 28641 16031
rect 28641 15997 28675 16031
rect 28675 15997 28684 16031
rect 28632 15988 28684 15997
rect 29828 15988 29880 16040
rect 31944 15988 31996 16040
rect 32220 15988 32272 16040
rect 36176 16124 36228 16176
rect 33324 16056 33376 16108
rect 37004 16192 37056 16244
rect 40960 16235 41012 16244
rect 40960 16201 40969 16235
rect 40969 16201 41003 16235
rect 41003 16201 41012 16235
rect 40960 16192 41012 16201
rect 38568 16124 38620 16176
rect 38752 16124 38804 16176
rect 37372 16056 37424 16108
rect 48320 16056 48372 16108
rect 48688 16099 48740 16108
rect 48688 16065 48697 16099
rect 48697 16065 48731 16099
rect 48731 16065 48740 16099
rect 48688 16056 48740 16065
rect 32772 15988 32824 16040
rect 26884 15852 26936 15904
rect 27344 15852 27396 15904
rect 33416 15920 33468 15972
rect 37464 16031 37516 16040
rect 37464 15997 37473 16031
rect 37473 15997 37507 16031
rect 37507 15997 37516 16031
rect 37464 15988 37516 15997
rect 38568 15988 38620 16040
rect 41788 15988 41840 16040
rect 30748 15852 30800 15904
rect 31392 15852 31444 15904
rect 31760 15852 31812 15904
rect 33692 15852 33744 15904
rect 34152 15852 34204 15904
rect 35164 15895 35216 15904
rect 35164 15861 35173 15895
rect 35173 15861 35207 15895
rect 35207 15861 35216 15895
rect 35164 15852 35216 15861
rect 37648 15920 37700 15972
rect 37188 15852 37240 15904
rect 40316 15852 40368 15904
rect 41604 15895 41656 15904
rect 41604 15861 41613 15895
rect 41613 15861 41647 15895
rect 41647 15861 41656 15895
rect 41604 15852 41656 15861
rect 49332 15895 49384 15904
rect 49332 15861 49341 15895
rect 49341 15861 49375 15895
rect 49375 15861 49384 15895
rect 49332 15852 49384 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 10692 15648 10744 15700
rect 12440 15648 12492 15700
rect 12992 15648 13044 15700
rect 14372 15648 14424 15700
rect 14924 15648 14976 15700
rect 16764 15691 16816 15700
rect 16764 15657 16773 15691
rect 16773 15657 16807 15691
rect 16807 15657 16816 15691
rect 16764 15648 16816 15657
rect 17868 15691 17920 15700
rect 17868 15657 17877 15691
rect 17877 15657 17911 15691
rect 17911 15657 17920 15691
rect 17868 15648 17920 15657
rect 18696 15648 18748 15700
rect 18788 15648 18840 15700
rect 19064 15648 19116 15700
rect 19340 15691 19392 15700
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20904 15648 20956 15700
rect 22560 15648 22612 15700
rect 25136 15648 25188 15700
rect 26148 15648 26200 15700
rect 26240 15648 26292 15700
rect 27068 15648 27120 15700
rect 28816 15648 28868 15700
rect 29092 15648 29144 15700
rect 29552 15648 29604 15700
rect 11060 15512 11112 15564
rect 13728 15580 13780 15632
rect 13912 15580 13964 15632
rect 15016 15580 15068 15632
rect 16488 15580 16540 15632
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 14464 15512 14516 15564
rect 14832 15555 14884 15564
rect 14832 15521 14841 15555
rect 14841 15521 14875 15555
rect 14875 15521 14884 15555
rect 14832 15512 14884 15521
rect 15752 15512 15804 15564
rect 10232 15444 10284 15496
rect 15108 15444 15160 15496
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 16028 15444 16080 15496
rect 17408 15512 17460 15564
rect 21364 15512 21416 15564
rect 21456 15512 21508 15564
rect 18420 15444 18472 15496
rect 18604 15487 18656 15496
rect 18604 15453 18613 15487
rect 18613 15453 18647 15487
rect 18647 15453 18656 15487
rect 18604 15444 18656 15453
rect 18972 15444 19024 15496
rect 21548 15444 21600 15496
rect 24860 15580 24912 15632
rect 22100 15512 22152 15564
rect 24308 15512 24360 15564
rect 26700 15580 26752 15632
rect 32588 15580 32640 15632
rect 25320 15512 25372 15564
rect 26608 15512 26660 15564
rect 31116 15512 31168 15564
rect 34428 15691 34480 15700
rect 34428 15657 34437 15691
rect 34437 15657 34471 15691
rect 34471 15657 34480 15691
rect 34428 15648 34480 15657
rect 37648 15648 37700 15700
rect 37740 15691 37792 15700
rect 37740 15657 37749 15691
rect 37749 15657 37783 15691
rect 37783 15657 37792 15691
rect 37740 15648 37792 15657
rect 41604 15648 41656 15700
rect 48320 15648 48372 15700
rect 49148 15691 49200 15700
rect 49148 15657 49157 15691
rect 49157 15657 49191 15691
rect 49191 15657 49200 15691
rect 49148 15648 49200 15657
rect 41788 15623 41840 15632
rect 41788 15589 41797 15623
rect 41797 15589 41831 15623
rect 41831 15589 41840 15623
rect 41788 15580 41840 15589
rect 27160 15444 27212 15496
rect 28172 15444 28224 15496
rect 30104 15444 30156 15496
rect 34796 15512 34848 15564
rect 35900 15512 35952 15564
rect 36176 15512 36228 15564
rect 34336 15444 34388 15496
rect 36452 15512 36504 15564
rect 37372 15512 37424 15564
rect 39488 15555 39540 15564
rect 39488 15521 39497 15555
rect 39497 15521 39531 15555
rect 39531 15521 39540 15555
rect 39488 15512 39540 15521
rect 40316 15555 40368 15564
rect 40316 15521 40325 15555
rect 40325 15521 40359 15555
rect 40359 15521 40368 15555
rect 40316 15512 40368 15521
rect 48596 15487 48648 15496
rect 48596 15453 48605 15487
rect 48605 15453 48639 15487
rect 48639 15453 48648 15487
rect 48596 15444 48648 15453
rect 49332 15487 49384 15496
rect 49332 15453 49341 15487
rect 49341 15453 49375 15487
rect 49375 15453 49384 15487
rect 49332 15444 49384 15453
rect 940 15376 992 15428
rect 4160 15376 4212 15428
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 11244 15308 11296 15360
rect 12624 15376 12676 15428
rect 13360 15419 13412 15428
rect 13360 15385 13369 15419
rect 13369 15385 13403 15419
rect 13403 15385 13412 15419
rect 13360 15376 13412 15385
rect 12992 15308 13044 15360
rect 13544 15308 13596 15360
rect 13820 15308 13872 15360
rect 14556 15308 14608 15360
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 15752 15308 15804 15360
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 17868 15308 17920 15360
rect 19708 15308 19760 15360
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 21272 15308 21324 15360
rect 21456 15308 21508 15360
rect 24124 15351 24176 15360
rect 24124 15317 24133 15351
rect 24133 15317 24167 15351
rect 24167 15317 24176 15351
rect 24124 15308 24176 15317
rect 25044 15419 25096 15428
rect 25044 15385 25053 15419
rect 25053 15385 25087 15419
rect 25087 15385 25096 15419
rect 25044 15376 25096 15385
rect 25688 15376 25740 15428
rect 26240 15419 26292 15428
rect 26240 15385 26249 15419
rect 26249 15385 26283 15419
rect 26283 15385 26292 15419
rect 26240 15376 26292 15385
rect 26332 15419 26384 15428
rect 26332 15385 26341 15419
rect 26341 15385 26375 15419
rect 26375 15385 26384 15419
rect 26332 15376 26384 15385
rect 28816 15376 28868 15428
rect 30472 15376 30524 15428
rect 30748 15419 30800 15428
rect 30748 15385 30757 15419
rect 30757 15385 30791 15419
rect 30791 15385 30800 15419
rect 30748 15376 30800 15385
rect 31760 15376 31812 15428
rect 25136 15351 25188 15360
rect 25136 15317 25145 15351
rect 25145 15317 25179 15351
rect 25179 15317 25188 15351
rect 25136 15308 25188 15317
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 26792 15308 26844 15360
rect 27160 15308 27212 15360
rect 27436 15351 27488 15360
rect 27436 15317 27445 15351
rect 27445 15317 27479 15351
rect 27479 15317 27488 15351
rect 27436 15308 27488 15317
rect 30012 15351 30064 15360
rect 30012 15317 30021 15351
rect 30021 15317 30055 15351
rect 30055 15317 30064 15351
rect 30012 15308 30064 15317
rect 30288 15308 30340 15360
rect 31668 15308 31720 15360
rect 32036 15308 32088 15360
rect 33048 15351 33100 15360
rect 33048 15317 33057 15351
rect 33057 15317 33091 15351
rect 33091 15317 33100 15351
rect 33048 15308 33100 15317
rect 34888 15376 34940 15428
rect 38752 15376 38804 15428
rect 33876 15351 33928 15360
rect 33876 15317 33885 15351
rect 33885 15317 33919 15351
rect 33919 15317 33928 15351
rect 33876 15308 33928 15317
rect 35900 15308 35952 15360
rect 37832 15308 37884 15360
rect 38568 15308 38620 15360
rect 41052 15376 41104 15428
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 11244 15104 11296 15156
rect 11796 15104 11848 15156
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 12992 15147 13044 15156
rect 12992 15113 13001 15147
rect 13001 15113 13035 15147
rect 13035 15113 13044 15147
rect 12992 15104 13044 15113
rect 13912 15104 13964 15156
rect 10876 15079 10928 15088
rect 10876 15045 10885 15079
rect 10885 15045 10919 15079
rect 10919 15045 10928 15079
rect 10876 15036 10928 15045
rect 11060 15079 11112 15088
rect 11060 15045 11069 15079
rect 11069 15045 11103 15079
rect 11103 15045 11112 15079
rect 11060 15036 11112 15045
rect 940 14968 992 15020
rect 4160 14968 4212 15020
rect 10692 14968 10744 15020
rect 12348 15011 12400 15020
rect 12348 14977 12357 15011
rect 12357 14977 12391 15011
rect 12391 14977 12400 15011
rect 12348 14968 12400 14977
rect 14372 15036 14424 15088
rect 15016 15104 15068 15156
rect 18788 15147 18840 15156
rect 18788 15113 18797 15147
rect 18797 15113 18831 15147
rect 18831 15113 18840 15147
rect 18788 15104 18840 15113
rect 19248 15104 19300 15156
rect 22836 15104 22888 15156
rect 23756 15104 23808 15156
rect 25136 15104 25188 15156
rect 25688 15104 25740 15156
rect 9772 14900 9824 14952
rect 11980 14832 12032 14884
rect 12072 14832 12124 14884
rect 10692 14764 10744 14816
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 15660 15036 15712 15088
rect 18604 15036 18656 15088
rect 20720 15036 20772 15088
rect 21824 15079 21876 15088
rect 21824 15045 21833 15079
rect 21833 15045 21867 15079
rect 21867 15045 21876 15079
rect 21824 15036 21876 15045
rect 25872 15036 25924 15088
rect 27068 15079 27120 15088
rect 27068 15045 27077 15079
rect 27077 15045 27111 15079
rect 27111 15045 27120 15079
rect 27068 15036 27120 15045
rect 29000 15036 29052 15088
rect 29828 15104 29880 15156
rect 30472 15104 30524 15156
rect 31300 15104 31352 15156
rect 19064 14968 19116 15020
rect 20904 14968 20956 15020
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 24124 14968 24176 15020
rect 24584 15011 24636 15020
rect 24584 14977 24593 15011
rect 24593 14977 24627 15011
rect 24627 14977 24636 15011
rect 24584 14968 24636 14977
rect 27344 14968 27396 15020
rect 27804 14968 27856 15020
rect 29552 14968 29604 15020
rect 33876 15147 33928 15156
rect 33876 15113 33885 15147
rect 33885 15113 33919 15147
rect 33919 15113 33928 15147
rect 33876 15104 33928 15113
rect 37464 15104 37516 15156
rect 34060 15036 34112 15088
rect 35808 15036 35860 15088
rect 36360 15036 36412 15088
rect 39948 15104 40000 15156
rect 13636 14900 13688 14952
rect 14280 14900 14332 14952
rect 14740 14900 14792 14952
rect 15200 14900 15252 14952
rect 16212 14764 16264 14816
rect 17224 14832 17276 14884
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 18052 14875 18104 14884
rect 18052 14841 18061 14875
rect 18061 14841 18095 14875
rect 18095 14841 18104 14875
rect 18052 14832 18104 14841
rect 20996 14900 21048 14952
rect 21088 14900 21140 14952
rect 18972 14832 19024 14884
rect 21548 14900 21600 14952
rect 24032 14900 24084 14952
rect 24216 14900 24268 14952
rect 17776 14764 17828 14816
rect 19248 14764 19300 14816
rect 20536 14764 20588 14816
rect 22744 14832 22796 14884
rect 21732 14764 21784 14816
rect 22192 14764 22244 14816
rect 24124 14764 24176 14816
rect 25872 14807 25924 14816
rect 25872 14773 25881 14807
rect 25881 14773 25915 14807
rect 25915 14773 25924 14807
rect 25872 14764 25924 14773
rect 26148 14832 26200 14884
rect 29736 14900 29788 14952
rect 29920 14900 29972 14952
rect 30288 14900 30340 14952
rect 31852 14900 31904 14952
rect 32496 14900 32548 14952
rect 33048 14900 33100 14952
rect 33416 14900 33468 14952
rect 29276 14832 29328 14884
rect 33784 14943 33836 14952
rect 33784 14909 33793 14943
rect 33793 14909 33827 14943
rect 33827 14909 33836 14943
rect 33784 14900 33836 14909
rect 33968 14832 34020 14884
rect 28080 14764 28132 14816
rect 28816 14764 28868 14816
rect 29552 14764 29604 14816
rect 30196 14807 30248 14816
rect 30196 14773 30205 14807
rect 30205 14773 30239 14807
rect 30239 14773 30248 14807
rect 30196 14764 30248 14773
rect 30472 14764 30524 14816
rect 34612 14832 34664 14884
rect 35348 14832 35400 14884
rect 34244 14807 34296 14816
rect 34244 14773 34253 14807
rect 34253 14773 34287 14807
rect 34287 14773 34296 14807
rect 34244 14764 34296 14773
rect 35440 14807 35492 14816
rect 35440 14773 35449 14807
rect 35449 14773 35483 14807
rect 35483 14773 35492 14807
rect 35440 14764 35492 14773
rect 37740 15079 37792 15088
rect 37740 15045 37749 15079
rect 37749 15045 37783 15079
rect 37783 15045 37792 15079
rect 37740 15036 37792 15045
rect 38752 15036 38804 15088
rect 40592 15036 40644 15088
rect 37372 14968 37424 15020
rect 38476 14900 38528 14952
rect 40224 14943 40276 14952
rect 40224 14909 40233 14943
rect 40233 14909 40267 14943
rect 40267 14909 40276 14943
rect 40224 14900 40276 14909
rect 49332 15011 49384 15020
rect 49332 14977 49341 15011
rect 49341 14977 49375 15011
rect 49375 14977 49384 15011
rect 49332 14968 49384 14977
rect 46940 14900 46992 14952
rect 36544 14832 36596 14884
rect 35992 14764 36044 14816
rect 48044 14875 48096 14884
rect 48044 14841 48053 14875
rect 48053 14841 48087 14875
rect 48087 14841 48096 14875
rect 48044 14832 48096 14841
rect 38752 14764 38804 14816
rect 45652 14764 45704 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 11428 14560 11480 14612
rect 12808 14560 12860 14612
rect 14556 14560 14608 14612
rect 17500 14560 17552 14612
rect 10232 14535 10284 14544
rect 10232 14501 10241 14535
rect 10241 14501 10275 14535
rect 10275 14501 10284 14535
rect 10232 14492 10284 14501
rect 18420 14560 18472 14612
rect 21548 14560 21600 14612
rect 22468 14560 22520 14612
rect 25504 14560 25556 14612
rect 26424 14560 26476 14612
rect 30564 14560 30616 14612
rect 31392 14560 31444 14612
rect 33600 14560 33652 14612
rect 34244 14560 34296 14612
rect 940 14424 992 14476
rect 13268 14424 13320 14476
rect 13452 14424 13504 14476
rect 19248 14492 19300 14544
rect 20168 14492 20220 14544
rect 15200 14424 15252 14476
rect 17040 14424 17092 14476
rect 20076 14467 20128 14476
rect 20076 14433 20085 14467
rect 20085 14433 20119 14467
rect 20119 14433 20128 14467
rect 20076 14424 20128 14433
rect 20628 14424 20680 14476
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 14280 14356 14332 14408
rect 17408 14356 17460 14408
rect 18052 14356 18104 14408
rect 18420 14356 18472 14408
rect 18788 14356 18840 14408
rect 19616 14356 19668 14408
rect 9956 14288 10008 14340
rect 10416 14331 10468 14340
rect 10416 14297 10425 14331
rect 10425 14297 10459 14331
rect 10459 14297 10468 14331
rect 10416 14288 10468 14297
rect 12808 14288 12860 14340
rect 10508 14220 10560 14272
rect 12716 14220 12768 14272
rect 13912 14220 13964 14272
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 16856 14263 16908 14272
rect 16856 14229 16865 14263
rect 16865 14229 16899 14263
rect 16899 14229 16908 14263
rect 16856 14220 16908 14229
rect 17868 14263 17920 14272
rect 17868 14229 17877 14263
rect 17877 14229 17911 14263
rect 17911 14229 17920 14263
rect 17868 14220 17920 14229
rect 19800 14288 19852 14340
rect 20536 14331 20588 14340
rect 20536 14297 20545 14331
rect 20545 14297 20579 14331
rect 20579 14297 20588 14331
rect 20536 14288 20588 14297
rect 22560 14492 22612 14544
rect 25044 14492 25096 14544
rect 21088 14467 21140 14476
rect 21088 14433 21097 14467
rect 21097 14433 21131 14467
rect 21131 14433 21140 14467
rect 21088 14424 21140 14433
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 21732 14424 21784 14476
rect 25780 14424 25832 14476
rect 26056 14424 26108 14476
rect 27804 14424 27856 14476
rect 28540 14492 28592 14544
rect 33784 14492 33836 14544
rect 36636 14603 36688 14612
rect 36636 14569 36645 14603
rect 36645 14569 36679 14603
rect 36679 14569 36688 14603
rect 36636 14560 36688 14569
rect 38384 14560 38436 14612
rect 38476 14560 38528 14612
rect 38844 14560 38896 14612
rect 22836 14356 22888 14408
rect 27344 14399 27396 14408
rect 27344 14365 27353 14399
rect 27353 14365 27387 14399
rect 27387 14365 27396 14399
rect 27344 14356 27396 14365
rect 29276 14424 29328 14476
rect 29644 14424 29696 14476
rect 30656 14424 30708 14476
rect 30840 14424 30892 14476
rect 31208 14424 31260 14476
rect 31484 14424 31536 14476
rect 32312 14424 32364 14476
rect 34796 14424 34848 14476
rect 37096 14424 37148 14476
rect 37372 14424 37424 14476
rect 21640 14288 21692 14340
rect 18512 14220 18564 14272
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 19708 14220 19760 14272
rect 23204 14263 23256 14272
rect 23204 14229 23213 14263
rect 23213 14229 23247 14263
rect 23247 14229 23256 14263
rect 23204 14220 23256 14229
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 25136 14263 25188 14272
rect 25136 14229 25145 14263
rect 25145 14229 25179 14263
rect 25179 14229 25188 14263
rect 25136 14220 25188 14229
rect 25688 14288 25740 14340
rect 28080 14399 28132 14408
rect 28080 14365 28089 14399
rect 28089 14365 28123 14399
rect 28123 14365 28132 14399
rect 28080 14356 28132 14365
rect 28632 14356 28684 14408
rect 30012 14356 30064 14408
rect 27712 14288 27764 14340
rect 29000 14263 29052 14272
rect 29000 14229 29009 14263
rect 29009 14229 29043 14263
rect 29043 14229 29052 14263
rect 29000 14220 29052 14229
rect 29368 14220 29420 14272
rect 30104 14263 30156 14272
rect 30104 14229 30113 14263
rect 30113 14229 30147 14263
rect 30147 14229 30156 14263
rect 30104 14220 30156 14229
rect 30564 14220 30616 14272
rect 32864 14356 32916 14408
rect 33692 14399 33744 14408
rect 33692 14365 33701 14399
rect 33701 14365 33735 14399
rect 33735 14365 33744 14399
rect 33692 14356 33744 14365
rect 39304 14399 39356 14408
rect 39304 14365 39313 14399
rect 39313 14365 39347 14399
rect 39347 14365 39356 14399
rect 39304 14356 39356 14365
rect 47952 14399 48004 14408
rect 47952 14365 47961 14399
rect 47961 14365 47995 14399
rect 47995 14365 48004 14399
rect 47952 14356 48004 14365
rect 49332 14399 49384 14408
rect 49332 14365 49341 14399
rect 49341 14365 49375 14399
rect 49375 14365 49384 14399
rect 49332 14356 49384 14365
rect 33324 14288 33376 14340
rect 34796 14288 34848 14340
rect 35164 14331 35216 14340
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 36452 14288 36504 14340
rect 38844 14288 38896 14340
rect 32588 14220 32640 14272
rect 32772 14220 32824 14272
rect 33416 14220 33468 14272
rect 34244 14220 34296 14272
rect 35440 14220 35492 14272
rect 36820 14220 36872 14272
rect 37188 14220 37240 14272
rect 37556 14220 37608 14272
rect 38476 14220 38528 14272
rect 39488 14263 39540 14272
rect 39488 14229 39497 14263
rect 39497 14229 39531 14263
rect 39531 14229 39540 14263
rect 39488 14220 39540 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 9864 14016 9916 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 11244 14016 11296 14068
rect 11888 14016 11940 14068
rect 14280 14016 14332 14068
rect 15660 14016 15712 14068
rect 16764 14059 16816 14068
rect 16764 14025 16773 14059
rect 16773 14025 16807 14059
rect 16807 14025 16816 14059
rect 16764 14016 16816 14025
rect 16856 14016 16908 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 19432 14016 19484 14068
rect 20168 14016 20220 14068
rect 21364 14016 21416 14068
rect 22100 14016 22152 14068
rect 1032 13948 1084 14000
rect 10508 13948 10560 14000
rect 13268 13991 13320 14000
rect 13268 13957 13277 13991
rect 13277 13957 13311 13991
rect 13311 13957 13320 13991
rect 13268 13948 13320 13957
rect 15016 13991 15068 14000
rect 15016 13957 15025 13991
rect 15025 13957 15059 13991
rect 15059 13957 15068 13991
rect 15016 13948 15068 13957
rect 19524 13948 19576 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 14648 13880 14700 13932
rect 16212 13880 16264 13932
rect 16764 13880 16816 13932
rect 18604 13880 18656 13932
rect 19616 13880 19668 13932
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 9772 13744 9824 13796
rect 12532 13812 12584 13864
rect 10784 13744 10836 13796
rect 12072 13676 12124 13728
rect 14464 13744 14516 13796
rect 17040 13812 17092 13864
rect 17500 13812 17552 13864
rect 16304 13744 16356 13796
rect 17868 13812 17920 13864
rect 13636 13676 13688 13728
rect 16028 13676 16080 13728
rect 16120 13676 16172 13728
rect 17408 13676 17460 13728
rect 17960 13744 18012 13796
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 18972 13812 19024 13864
rect 22192 13948 22244 14000
rect 21640 13880 21692 13932
rect 23204 14016 23256 14068
rect 25320 14016 25372 14068
rect 25504 14016 25556 14068
rect 25688 13948 25740 14000
rect 26516 14016 26568 14068
rect 27620 14059 27672 14068
rect 27620 14025 27629 14059
rect 27629 14025 27663 14059
rect 27663 14025 27672 14059
rect 27620 14016 27672 14025
rect 27804 14016 27856 14068
rect 30012 14016 30064 14068
rect 31116 14016 31168 14068
rect 41328 14016 41380 14068
rect 47216 14016 47268 14068
rect 28816 13948 28868 14000
rect 34704 13948 34756 14000
rect 34888 13991 34940 14000
rect 34888 13957 34897 13991
rect 34897 13957 34931 13991
rect 34931 13957 34940 13991
rect 34888 13948 34940 13957
rect 35164 13948 35216 14000
rect 37004 13948 37056 14000
rect 37280 13948 37332 14000
rect 38844 13948 38896 14000
rect 39488 13948 39540 14000
rect 47860 13948 47912 14000
rect 24492 13880 24544 13932
rect 28908 13923 28960 13932
rect 28908 13889 28917 13923
rect 28917 13889 28951 13923
rect 28951 13889 28960 13923
rect 28908 13880 28960 13889
rect 31116 13923 31168 13932
rect 31116 13889 31125 13923
rect 31125 13889 31159 13923
rect 31159 13889 31168 13923
rect 31116 13880 31168 13889
rect 31484 13880 31536 13932
rect 31760 13880 31812 13932
rect 35256 13880 35308 13932
rect 35624 13880 35676 13932
rect 36176 13880 36228 13932
rect 37188 13880 37240 13932
rect 40224 13880 40276 13932
rect 45652 13923 45704 13932
rect 45652 13889 45661 13923
rect 45661 13889 45695 13923
rect 45695 13889 45704 13923
rect 45652 13880 45704 13889
rect 21916 13812 21968 13864
rect 19708 13676 19760 13728
rect 19984 13719 20036 13728
rect 19984 13685 20014 13719
rect 20014 13685 20036 13719
rect 22008 13744 22060 13796
rect 23940 13812 23992 13864
rect 27344 13812 27396 13864
rect 24308 13744 24360 13796
rect 28448 13744 28500 13796
rect 29092 13744 29144 13796
rect 32496 13812 32548 13864
rect 32588 13812 32640 13864
rect 33416 13812 33468 13864
rect 34060 13855 34112 13864
rect 34060 13821 34069 13855
rect 34069 13821 34103 13855
rect 34103 13821 34112 13855
rect 34060 13812 34112 13821
rect 34704 13744 34756 13796
rect 36636 13812 36688 13864
rect 36452 13744 36504 13796
rect 46756 13812 46808 13864
rect 46940 13812 46992 13864
rect 49332 13923 49384 13932
rect 49332 13889 49341 13923
rect 49341 13889 49375 13923
rect 49375 13889 49384 13923
rect 49332 13880 49384 13889
rect 47676 13855 47728 13864
rect 47676 13821 47685 13855
rect 47685 13821 47719 13855
rect 47719 13821 47728 13855
rect 47676 13812 47728 13821
rect 47768 13812 47820 13864
rect 38200 13744 38252 13796
rect 19984 13676 20036 13685
rect 22744 13676 22796 13728
rect 27436 13676 27488 13728
rect 30840 13676 30892 13728
rect 36176 13676 36228 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 13452 13472 13504 13524
rect 14004 13472 14056 13524
rect 14924 13472 14976 13524
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 10784 13379 10836 13388
rect 10784 13345 10793 13379
rect 10793 13345 10827 13379
rect 10827 13345 10836 13379
rect 10784 13336 10836 13345
rect 12532 13379 12584 13388
rect 12532 13345 12541 13379
rect 12541 13345 12575 13379
rect 12575 13345 12584 13379
rect 12532 13336 12584 13345
rect 12808 13336 12860 13388
rect 14832 13336 14884 13388
rect 17960 13472 18012 13524
rect 18328 13472 18380 13524
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 20076 13472 20128 13524
rect 20260 13472 20312 13524
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 20352 13404 20404 13456
rect 15476 13379 15528 13388
rect 15476 13345 15485 13379
rect 15485 13345 15519 13379
rect 15519 13345 15528 13379
rect 15476 13336 15528 13345
rect 15752 13336 15804 13388
rect 18972 13336 19024 13388
rect 19984 13336 20036 13388
rect 20996 13336 21048 13388
rect 21548 13379 21600 13388
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 22744 13472 22796 13524
rect 23664 13472 23716 13524
rect 25596 13515 25648 13524
rect 25596 13481 25605 13515
rect 25605 13481 25639 13515
rect 25639 13481 25648 13515
rect 25596 13472 25648 13481
rect 28356 13472 28408 13524
rect 28908 13472 28960 13524
rect 33784 13472 33836 13524
rect 36268 13472 36320 13524
rect 24308 13404 24360 13456
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 14924 13268 14976 13320
rect 9036 13200 9088 13252
rect 11060 13243 11112 13252
rect 11060 13209 11069 13243
rect 11069 13209 11103 13243
rect 11103 13209 11112 13243
rect 11060 13200 11112 13209
rect 11704 13132 11756 13184
rect 15016 13200 15068 13252
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 16304 13268 16356 13320
rect 18052 13268 18104 13320
rect 13728 13132 13780 13184
rect 14004 13132 14056 13184
rect 14096 13132 14148 13184
rect 15844 13132 15896 13184
rect 16764 13200 16816 13252
rect 17132 13200 17184 13252
rect 20996 13200 21048 13252
rect 21640 13200 21692 13252
rect 23388 13200 23440 13252
rect 23848 13268 23900 13320
rect 25228 13404 25280 13456
rect 26056 13336 26108 13388
rect 29920 13404 29972 13456
rect 29828 13379 29880 13388
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 30380 13336 30432 13388
rect 25136 13268 25188 13320
rect 27804 13268 27856 13320
rect 24216 13200 24268 13252
rect 19800 13132 19852 13184
rect 19984 13175 20036 13184
rect 19984 13141 19993 13175
rect 19993 13141 20027 13175
rect 20027 13141 20036 13175
rect 19984 13132 20036 13141
rect 21272 13175 21324 13184
rect 21272 13141 21281 13175
rect 21281 13141 21315 13175
rect 21315 13141 21324 13175
rect 21272 13132 21324 13141
rect 23664 13132 23716 13184
rect 23848 13132 23900 13184
rect 25872 13200 25924 13252
rect 26700 13200 26752 13252
rect 28448 13200 28500 13252
rect 29000 13268 29052 13320
rect 30196 13268 30248 13320
rect 31576 13336 31628 13388
rect 34428 13404 34480 13456
rect 33692 13336 33744 13388
rect 37832 13472 37884 13524
rect 38200 13515 38252 13524
rect 38200 13481 38209 13515
rect 38209 13481 38243 13515
rect 38243 13481 38252 13515
rect 38200 13472 38252 13481
rect 38844 13472 38896 13524
rect 39488 13472 39540 13524
rect 47768 13472 47820 13524
rect 36728 13336 36780 13388
rect 39580 13336 39632 13388
rect 29736 13200 29788 13252
rect 31484 13268 31536 13320
rect 34060 13268 34112 13320
rect 34888 13268 34940 13320
rect 24492 13175 24544 13184
rect 24492 13141 24501 13175
rect 24501 13141 24535 13175
rect 24535 13141 24544 13175
rect 24492 13132 24544 13141
rect 25964 13132 26016 13184
rect 26056 13175 26108 13184
rect 26056 13141 26065 13175
rect 26065 13141 26099 13175
rect 26099 13141 26108 13175
rect 26056 13132 26108 13141
rect 27712 13175 27764 13184
rect 27712 13141 27721 13175
rect 27721 13141 27755 13175
rect 27755 13141 27764 13175
rect 27712 13132 27764 13141
rect 28540 13132 28592 13184
rect 28724 13175 28776 13184
rect 28724 13141 28733 13175
rect 28733 13141 28767 13175
rect 28767 13141 28776 13175
rect 28724 13132 28776 13141
rect 33968 13200 34020 13252
rect 35900 13200 35952 13252
rect 31668 13132 31720 13184
rect 33416 13132 33468 13184
rect 34152 13132 34204 13184
rect 35164 13175 35216 13184
rect 35164 13141 35173 13175
rect 35173 13141 35207 13175
rect 35207 13141 35216 13175
rect 35164 13132 35216 13141
rect 35716 13132 35768 13184
rect 41328 13311 41380 13320
rect 41328 13277 41337 13311
rect 41337 13277 41371 13311
rect 41371 13277 41380 13311
rect 41328 13268 41380 13277
rect 46756 13268 46808 13320
rect 49148 13311 49200 13320
rect 49148 13277 49157 13311
rect 49157 13277 49191 13311
rect 49191 13277 49200 13311
rect 49148 13268 49200 13277
rect 36636 13200 36688 13252
rect 38844 13200 38896 13252
rect 37464 13132 37516 13184
rect 37648 13132 37700 13184
rect 39304 13132 39356 13184
rect 45928 13132 45980 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 9496 12928 9548 12980
rect 11336 12971 11388 12980
rect 11336 12937 11345 12971
rect 11345 12937 11379 12971
rect 11379 12937 11388 12971
rect 11336 12928 11388 12937
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 12532 12928 12584 12980
rect 12900 12928 12952 12980
rect 13268 12928 13320 12980
rect 13636 12928 13688 12980
rect 1308 12860 1360 12912
rect 11704 12860 11756 12912
rect 14004 12860 14056 12912
rect 14556 12903 14608 12912
rect 14556 12869 14565 12903
rect 14565 12869 14599 12903
rect 14599 12869 14608 12903
rect 14556 12860 14608 12869
rect 15200 12928 15252 12980
rect 16396 12860 16448 12912
rect 16672 12903 16724 12912
rect 16672 12869 16681 12903
rect 16681 12869 16715 12903
rect 16715 12869 16724 12903
rect 16672 12860 16724 12869
rect 17040 12860 17092 12912
rect 18972 12860 19024 12912
rect 20904 12928 20956 12980
rect 23480 12928 23532 12980
rect 23664 12928 23716 12980
rect 1308 12656 1360 12708
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 15752 12792 15804 12844
rect 16764 12792 16816 12844
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17316 12792 17368 12844
rect 18880 12792 18932 12844
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 19800 12792 19852 12844
rect 20996 12792 21048 12844
rect 21916 12792 21968 12844
rect 13820 12724 13872 12776
rect 15936 12724 15988 12776
rect 16580 12724 16632 12776
rect 19524 12724 19576 12776
rect 19708 12767 19760 12776
rect 19708 12733 19717 12767
rect 19717 12733 19751 12767
rect 19751 12733 19760 12767
rect 19708 12724 19760 12733
rect 20260 12724 20312 12776
rect 20444 12724 20496 12776
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 22744 12767 22796 12776
rect 22744 12733 22753 12767
rect 22753 12733 22787 12767
rect 22787 12733 22796 12767
rect 22744 12724 22796 12733
rect 22928 12767 22980 12776
rect 22928 12733 22937 12767
rect 22937 12733 22971 12767
rect 22971 12733 22980 12767
rect 22928 12724 22980 12733
rect 15292 12699 15344 12708
rect 15292 12665 15301 12699
rect 15301 12665 15335 12699
rect 15335 12665 15344 12699
rect 15292 12656 15344 12665
rect 16396 12656 16448 12708
rect 2320 12631 2372 12640
rect 2320 12597 2329 12631
rect 2329 12597 2363 12631
rect 2363 12597 2372 12631
rect 2320 12588 2372 12597
rect 2872 12588 2924 12640
rect 12624 12588 12676 12640
rect 13820 12588 13872 12640
rect 14096 12588 14148 12640
rect 14188 12588 14240 12640
rect 15016 12588 15068 12640
rect 16580 12588 16632 12640
rect 17040 12588 17092 12640
rect 20996 12656 21048 12708
rect 21456 12656 21508 12708
rect 23848 12860 23900 12912
rect 23572 12724 23624 12776
rect 23664 12724 23716 12776
rect 24400 12928 24452 12980
rect 24584 12928 24636 12980
rect 24860 12860 24912 12912
rect 25320 12903 25372 12912
rect 25320 12869 25329 12903
rect 25329 12869 25363 12903
rect 25363 12869 25372 12903
rect 25320 12860 25372 12869
rect 25964 12928 26016 12980
rect 27068 12928 27120 12980
rect 28540 12928 28592 12980
rect 24952 12724 25004 12776
rect 25228 12724 25280 12776
rect 26240 12860 26292 12912
rect 27160 12903 27212 12912
rect 27160 12869 27169 12903
rect 27169 12869 27203 12903
rect 27203 12869 27212 12903
rect 27160 12860 27212 12869
rect 28448 12860 28500 12912
rect 29368 12860 29420 12912
rect 29736 12860 29788 12912
rect 31760 12928 31812 12980
rect 34060 12928 34112 12980
rect 32036 12860 32088 12912
rect 32128 12860 32180 12912
rect 32772 12860 32824 12912
rect 33416 12903 33468 12912
rect 33416 12869 33425 12903
rect 33425 12869 33459 12903
rect 33459 12869 33468 12903
rect 33416 12860 33468 12869
rect 34428 12860 34480 12912
rect 34980 12928 35032 12980
rect 36728 12928 36780 12980
rect 37188 12928 37240 12980
rect 40316 12928 40368 12980
rect 34888 12860 34940 12912
rect 36912 12860 36964 12912
rect 30012 12835 30064 12844
rect 30012 12801 30021 12835
rect 30021 12801 30055 12835
rect 30055 12801 30064 12835
rect 30012 12792 30064 12801
rect 31392 12792 31444 12844
rect 31760 12792 31812 12844
rect 33324 12792 33376 12844
rect 34612 12792 34664 12844
rect 29644 12724 29696 12776
rect 32036 12724 32088 12776
rect 24124 12656 24176 12708
rect 33692 12724 33744 12776
rect 35164 12724 35216 12776
rect 35348 12724 35400 12776
rect 22928 12588 22980 12640
rect 24860 12588 24912 12640
rect 25688 12588 25740 12640
rect 25964 12631 26016 12640
rect 25964 12597 25973 12631
rect 25973 12597 26007 12631
rect 26007 12597 26016 12631
rect 25964 12588 26016 12597
rect 28816 12588 28868 12640
rect 34520 12656 34572 12708
rect 35808 12724 35860 12776
rect 37648 12860 37700 12912
rect 37464 12835 37516 12844
rect 37464 12801 37473 12835
rect 37473 12801 37507 12835
rect 37507 12801 37516 12835
rect 37464 12792 37516 12801
rect 38844 12792 38896 12844
rect 40040 12835 40092 12844
rect 40040 12801 40049 12835
rect 40049 12801 40083 12835
rect 40083 12801 40092 12835
rect 40040 12792 40092 12801
rect 45928 12835 45980 12844
rect 45928 12801 45937 12835
rect 45937 12801 45971 12835
rect 45971 12801 45980 12835
rect 45928 12792 45980 12801
rect 47216 12792 47268 12844
rect 49148 12835 49200 12844
rect 49148 12801 49157 12835
rect 49157 12801 49191 12835
rect 49191 12801 49200 12835
rect 49148 12792 49200 12801
rect 36452 12767 36504 12776
rect 36452 12733 36461 12767
rect 36461 12733 36495 12767
rect 36495 12733 36504 12767
rect 36452 12724 36504 12733
rect 37188 12724 37240 12776
rect 38292 12724 38344 12776
rect 39304 12724 39356 12776
rect 32312 12588 32364 12640
rect 32588 12588 32640 12640
rect 32864 12588 32916 12640
rect 35808 12588 35860 12640
rect 36912 12588 36964 12640
rect 46940 12656 46992 12708
rect 39120 12588 39172 12640
rect 47952 12588 48004 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 4344 12384 4396 12436
rect 11796 12384 11848 12436
rect 13544 12384 13596 12436
rect 13728 12384 13780 12436
rect 14188 12384 14240 12436
rect 11060 12316 11112 12368
rect 5816 12248 5868 12300
rect 10784 12248 10836 12300
rect 13360 12316 13412 12368
rect 16120 12384 16172 12436
rect 17868 12384 17920 12436
rect 19340 12384 19392 12436
rect 21732 12384 21784 12436
rect 26056 12384 26108 12436
rect 26332 12427 26384 12436
rect 26332 12393 26341 12427
rect 26341 12393 26375 12427
rect 26375 12393 26384 12427
rect 26332 12384 26384 12393
rect 26976 12384 27028 12436
rect 31760 12384 31812 12436
rect 16212 12316 16264 12368
rect 16396 12316 16448 12368
rect 13728 12248 13780 12300
rect 15292 12248 15344 12300
rect 15752 12248 15804 12300
rect 2228 12180 2280 12232
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 11612 12180 11664 12232
rect 9772 12155 9824 12164
rect 9772 12121 9781 12155
rect 9781 12121 9815 12155
rect 9815 12121 9824 12155
rect 9772 12112 9824 12121
rect 11060 12112 11112 12164
rect 13544 12112 13596 12164
rect 14464 12112 14516 12164
rect 16948 12248 17000 12300
rect 17408 12316 17460 12368
rect 17500 12248 17552 12300
rect 19432 12248 19484 12300
rect 17040 12180 17092 12232
rect 19064 12180 19116 12232
rect 21272 12316 21324 12368
rect 23756 12316 23808 12368
rect 25964 12316 26016 12368
rect 26700 12359 26752 12368
rect 26700 12325 26709 12359
rect 26709 12325 26743 12359
rect 26743 12325 26752 12359
rect 26700 12316 26752 12325
rect 31024 12316 31076 12368
rect 39304 12427 39356 12436
rect 39304 12393 39313 12427
rect 39313 12393 39347 12427
rect 39347 12393 39356 12427
rect 39304 12384 39356 12393
rect 39488 12427 39540 12436
rect 39488 12393 39497 12427
rect 39497 12393 39531 12427
rect 39531 12393 39540 12427
rect 39488 12384 39540 12393
rect 19892 12248 19944 12300
rect 20996 12291 21048 12300
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 18788 12112 18840 12164
rect 18880 12155 18932 12164
rect 18880 12121 18889 12155
rect 18889 12121 18923 12155
rect 18923 12121 18932 12155
rect 18880 12112 18932 12121
rect 19524 12112 19576 12164
rect 20536 12180 20588 12232
rect 21180 12180 21232 12232
rect 21732 12180 21784 12232
rect 22376 12291 22428 12300
rect 22376 12257 22385 12291
rect 22385 12257 22419 12291
rect 22419 12257 22428 12291
rect 22376 12248 22428 12257
rect 23480 12248 23532 12300
rect 23664 12248 23716 12300
rect 24492 12248 24544 12300
rect 24952 12248 25004 12300
rect 12992 12044 13044 12096
rect 14372 12044 14424 12096
rect 15660 12044 15712 12096
rect 16764 12087 16816 12096
rect 16764 12053 16773 12087
rect 16773 12053 16807 12087
rect 16807 12053 16816 12087
rect 16764 12044 16816 12053
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 20076 12112 20128 12164
rect 21456 12112 21508 12164
rect 17224 12044 17276 12053
rect 20904 12044 20956 12096
rect 21180 12087 21232 12096
rect 21180 12053 21189 12087
rect 21189 12053 21223 12087
rect 21223 12053 21232 12087
rect 24124 12180 24176 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 27160 12291 27212 12300
rect 27160 12257 27169 12291
rect 27169 12257 27203 12291
rect 27203 12257 27212 12291
rect 27160 12248 27212 12257
rect 27344 12248 27396 12300
rect 30012 12248 30064 12300
rect 31484 12248 31536 12300
rect 27620 12180 27672 12232
rect 28816 12180 28868 12232
rect 31116 12180 31168 12232
rect 21180 12044 21232 12053
rect 23388 12044 23440 12096
rect 26884 12112 26936 12164
rect 27068 12112 27120 12164
rect 27528 12112 27580 12164
rect 29920 12112 29972 12164
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 31392 12044 31444 12096
rect 33876 12291 33928 12300
rect 33876 12257 33885 12291
rect 33885 12257 33919 12291
rect 33919 12257 33928 12291
rect 33876 12248 33928 12257
rect 38384 12291 38436 12300
rect 38384 12257 38393 12291
rect 38393 12257 38427 12291
rect 38427 12257 38436 12291
rect 38384 12248 38436 12257
rect 38752 12248 38804 12300
rect 39948 12316 40000 12368
rect 47400 12316 47452 12368
rect 32128 12223 32180 12232
rect 32128 12189 32137 12223
rect 32137 12189 32171 12223
rect 32171 12189 32180 12223
rect 32128 12180 32180 12189
rect 34152 12180 34204 12232
rect 34888 12223 34940 12232
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 37096 12180 37148 12232
rect 49148 12291 49200 12300
rect 49148 12257 49157 12291
rect 49157 12257 49191 12291
rect 49191 12257 49200 12291
rect 49148 12248 49200 12257
rect 32312 12112 32364 12164
rect 32864 12112 32916 12164
rect 34612 12112 34664 12164
rect 35164 12155 35216 12164
rect 35164 12121 35173 12155
rect 35173 12121 35207 12155
rect 35207 12121 35216 12155
rect 35164 12112 35216 12121
rect 34336 12044 34388 12096
rect 36544 12044 36596 12096
rect 36728 12044 36780 12096
rect 37280 12044 37332 12096
rect 40408 12112 40460 12164
rect 38660 12087 38712 12096
rect 38660 12053 38669 12087
rect 38669 12053 38703 12087
rect 38703 12053 38712 12087
rect 38660 12044 38712 12053
rect 40960 12087 41012 12096
rect 40960 12053 40969 12087
rect 40969 12053 41003 12087
rect 41003 12053 41012 12087
rect 40960 12044 41012 12053
rect 47952 12223 48004 12232
rect 47952 12189 47961 12223
rect 47961 12189 47995 12223
rect 47995 12189 48004 12223
rect 47952 12180 48004 12189
rect 46112 12087 46164 12096
rect 46112 12053 46121 12087
rect 46121 12053 46155 12087
rect 46155 12053 46164 12087
rect 46112 12044 46164 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 2228 11883 2280 11892
rect 2228 11849 2237 11883
rect 2237 11849 2271 11883
rect 2271 11849 2280 11883
rect 2228 11840 2280 11849
rect 4252 11840 4304 11892
rect 11704 11840 11756 11892
rect 12072 11840 12124 11892
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 13636 11840 13688 11892
rect 14280 11883 14332 11892
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 14648 11840 14700 11892
rect 17960 11840 18012 11892
rect 19984 11840 20036 11892
rect 20720 11883 20772 11892
rect 20720 11849 20729 11883
rect 20729 11849 20763 11883
rect 20763 11849 20772 11883
rect 20720 11840 20772 11849
rect 22008 11840 22060 11892
rect 11244 11772 11296 11824
rect 1308 11704 1360 11756
rect 2320 11704 2372 11756
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 14372 11772 14424 11824
rect 12992 11704 13044 11756
rect 15384 11772 15436 11824
rect 11796 11636 11848 11688
rect 14740 11704 14792 11756
rect 14280 11636 14332 11688
rect 14556 11636 14608 11688
rect 11888 11500 11940 11552
rect 15476 11568 15528 11620
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 14832 11500 14884 11552
rect 15384 11500 15436 11552
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 16948 11772 17000 11824
rect 20444 11772 20496 11824
rect 20536 11772 20588 11824
rect 22376 11840 22428 11892
rect 24492 11840 24544 11892
rect 27344 11840 27396 11892
rect 28632 11840 28684 11892
rect 22192 11772 22244 11824
rect 18696 11704 18748 11756
rect 19800 11747 19852 11756
rect 19800 11713 19809 11747
rect 19809 11713 19843 11747
rect 19843 11713 19852 11747
rect 19800 11704 19852 11713
rect 18788 11636 18840 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 20812 11704 20864 11756
rect 22468 11704 22520 11756
rect 24124 11772 24176 11824
rect 25596 11772 25648 11824
rect 26976 11772 27028 11824
rect 28448 11772 28500 11824
rect 31116 11840 31168 11892
rect 31852 11840 31904 11892
rect 32404 11840 32456 11892
rect 32680 11883 32732 11892
rect 32680 11849 32689 11883
rect 32689 11849 32723 11883
rect 32723 11849 32732 11883
rect 32680 11840 32732 11849
rect 25688 11704 25740 11756
rect 25780 11704 25832 11756
rect 20352 11636 20404 11688
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 21180 11636 21232 11645
rect 21548 11636 21600 11688
rect 23480 11636 23532 11688
rect 26332 11636 26384 11688
rect 18696 11500 18748 11552
rect 19156 11543 19208 11552
rect 19156 11509 19165 11543
rect 19165 11509 19199 11543
rect 19199 11509 19208 11543
rect 19156 11500 19208 11509
rect 21272 11500 21324 11552
rect 21640 11500 21692 11552
rect 22008 11500 22060 11552
rect 22468 11500 22520 11552
rect 24676 11500 24728 11552
rect 24768 11500 24820 11552
rect 26148 11568 26200 11620
rect 27436 11679 27488 11688
rect 27436 11645 27445 11679
rect 27445 11645 27479 11679
rect 27479 11645 27488 11679
rect 27436 11636 27488 11645
rect 27804 11568 27856 11620
rect 31392 11772 31444 11824
rect 33784 11840 33836 11892
rect 34336 11840 34388 11892
rect 31116 11747 31168 11756
rect 31116 11713 31125 11747
rect 31125 11713 31159 11747
rect 31159 11713 31168 11747
rect 31116 11704 31168 11713
rect 35072 11772 35124 11824
rect 35256 11840 35308 11892
rect 38660 11883 38712 11892
rect 38660 11849 38669 11883
rect 38669 11849 38703 11883
rect 38703 11849 38712 11883
rect 38660 11840 38712 11849
rect 39120 11883 39172 11892
rect 39120 11849 39129 11883
rect 39129 11849 39163 11883
rect 39163 11849 39172 11883
rect 39120 11840 39172 11849
rect 35716 11772 35768 11824
rect 36728 11772 36780 11824
rect 28816 11636 28868 11688
rect 28908 11568 28960 11620
rect 30288 11679 30340 11688
rect 30288 11645 30297 11679
rect 30297 11645 30331 11679
rect 30331 11645 30340 11679
rect 30288 11636 30340 11645
rect 30840 11679 30892 11688
rect 30840 11645 30849 11679
rect 30849 11645 30883 11679
rect 30883 11645 30892 11679
rect 30840 11636 30892 11645
rect 31760 11636 31812 11688
rect 32864 11636 32916 11688
rect 33692 11704 33744 11756
rect 36820 11704 36872 11756
rect 39028 11747 39080 11756
rect 39028 11713 39037 11747
rect 39037 11713 39071 11747
rect 39071 11713 39080 11747
rect 39028 11704 39080 11713
rect 33968 11636 34020 11688
rect 34244 11636 34296 11688
rect 34888 11636 34940 11688
rect 31392 11568 31444 11620
rect 27252 11500 27304 11552
rect 30196 11500 30248 11552
rect 31484 11500 31536 11552
rect 34244 11543 34296 11552
rect 34244 11509 34253 11543
rect 34253 11509 34287 11543
rect 34287 11509 34296 11543
rect 34244 11500 34296 11509
rect 34428 11500 34480 11552
rect 36452 11636 36504 11688
rect 36636 11636 36688 11688
rect 39948 11815 40000 11824
rect 39948 11781 39957 11815
rect 39957 11781 39991 11815
rect 39991 11781 40000 11815
rect 39948 11772 40000 11781
rect 40408 11815 40460 11824
rect 40408 11781 40417 11815
rect 40417 11781 40451 11815
rect 40451 11781 40460 11815
rect 40408 11772 40460 11781
rect 40960 11772 41012 11824
rect 49148 11815 49200 11824
rect 49148 11781 49157 11815
rect 49157 11781 49191 11815
rect 49191 11781 49200 11815
rect 49148 11772 49200 11781
rect 46112 11704 46164 11756
rect 38384 11568 38436 11620
rect 35624 11500 35676 11552
rect 40224 11500 40276 11552
rect 46664 11568 46716 11620
rect 47032 11500 47084 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 11428 11296 11480 11348
rect 12440 11296 12492 11348
rect 1308 11228 1360 11280
rect 2688 11228 2740 11280
rect 11244 11228 11296 11280
rect 1216 11092 1268 11144
rect 11060 11160 11112 11212
rect 11796 11160 11848 11212
rect 13544 11296 13596 11348
rect 13912 11296 13964 11348
rect 14464 11296 14516 11348
rect 15568 11296 15620 11348
rect 16672 11296 16724 11348
rect 18880 11296 18932 11348
rect 22468 11296 22520 11348
rect 23296 11339 23348 11348
rect 23296 11305 23305 11339
rect 23305 11305 23339 11339
rect 23339 11305 23348 11339
rect 23296 11296 23348 11305
rect 18420 11228 18472 11280
rect 14740 11160 14792 11212
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15108 11160 15160 11212
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 15844 11203 15896 11212
rect 15844 11169 15853 11203
rect 15853 11169 15887 11203
rect 15887 11169 15896 11203
rect 15844 11160 15896 11169
rect 17408 11203 17460 11212
rect 17408 11169 17417 11203
rect 17417 11169 17451 11203
rect 17451 11169 17460 11203
rect 17408 11160 17460 11169
rect 17684 11160 17736 11212
rect 19156 11228 19208 11280
rect 20352 11228 20404 11280
rect 20444 11271 20496 11280
rect 20444 11237 20453 11271
rect 20453 11237 20487 11271
rect 20487 11237 20496 11271
rect 20444 11228 20496 11237
rect 19432 11160 19484 11212
rect 20076 11160 20128 11212
rect 23756 11203 23808 11212
rect 2780 11092 2832 11144
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 16856 11092 16908 11144
rect 19064 11092 19116 11144
rect 23756 11169 23765 11203
rect 23765 11169 23799 11203
rect 23799 11169 23808 11203
rect 23756 11160 23808 11169
rect 25228 11296 25280 11348
rect 26608 11296 26660 11348
rect 28540 11296 28592 11348
rect 28816 11296 28868 11348
rect 30472 11339 30524 11348
rect 30472 11305 30481 11339
rect 30481 11305 30515 11339
rect 30515 11305 30524 11339
rect 30472 11296 30524 11305
rect 31392 11296 31444 11348
rect 33324 11296 33376 11348
rect 34428 11296 34480 11348
rect 24492 11160 24544 11212
rect 11796 11024 11848 11076
rect 13452 11024 13504 11076
rect 14740 11067 14792 11076
rect 14740 11033 14749 11067
rect 14749 11033 14783 11067
rect 14783 11033 14792 11067
rect 14740 11024 14792 11033
rect 16672 11024 16724 11076
rect 18512 11024 18564 11076
rect 11704 10956 11756 11008
rect 12532 10956 12584 11008
rect 15292 10956 15344 11008
rect 17132 10956 17184 11008
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 17316 10956 17368 11008
rect 18788 11024 18840 11076
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 29368 11092 29420 11144
rect 31024 11228 31076 11280
rect 32864 11271 32916 11280
rect 32864 11237 32873 11271
rect 32873 11237 32907 11271
rect 32907 11237 32916 11271
rect 32864 11228 32916 11237
rect 34244 11228 34296 11280
rect 30196 11160 30248 11212
rect 32128 11160 32180 11212
rect 35716 11160 35768 11212
rect 30288 11092 30340 11144
rect 33324 11135 33376 11144
rect 33324 11101 33333 11135
rect 33333 11101 33367 11135
rect 33367 11101 33376 11135
rect 33324 11092 33376 11101
rect 37464 11160 37516 11212
rect 38660 11296 38712 11348
rect 39488 11296 39540 11348
rect 39580 11339 39632 11348
rect 39580 11305 39589 11339
rect 39589 11305 39623 11339
rect 39623 11305 39632 11339
rect 39580 11296 39632 11305
rect 44364 11296 44416 11348
rect 39580 11092 39632 11144
rect 40224 11092 40276 11144
rect 49148 11203 49200 11212
rect 49148 11169 49157 11203
rect 49157 11169 49191 11203
rect 49191 11169 49200 11203
rect 49148 11160 49200 11169
rect 46940 11092 46992 11144
rect 20168 11024 20220 11076
rect 20444 11024 20496 11076
rect 23572 11024 23624 11076
rect 23940 11024 23992 11076
rect 26700 11024 26752 11076
rect 27160 11067 27212 11076
rect 27160 11033 27169 11067
rect 27169 11033 27203 11067
rect 27203 11033 27212 11067
rect 27160 11024 27212 11033
rect 28540 11024 28592 11076
rect 28908 11024 28960 11076
rect 29460 11024 29512 11076
rect 19800 10956 19852 11008
rect 25596 10956 25648 11008
rect 29000 10956 29052 11008
rect 30380 11024 30432 11076
rect 31300 11024 31352 11076
rect 31484 11024 31536 11076
rect 30840 10956 30892 11008
rect 31576 10956 31628 11008
rect 34796 11024 34848 11076
rect 35532 11024 35584 11076
rect 35900 11024 35952 11076
rect 38384 11024 38436 11076
rect 47216 11024 47268 11076
rect 46112 10956 46164 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 2780 10752 2832 10804
rect 11796 10752 11848 10804
rect 12808 10752 12860 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 14004 10684 14056 10736
rect 1308 10616 1360 10668
rect 1216 10548 1268 10600
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 12072 10616 12124 10668
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 15844 10752 15896 10804
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 18144 10752 18196 10804
rect 16764 10684 16816 10736
rect 17592 10727 17644 10736
rect 17592 10693 17601 10727
rect 17601 10693 17635 10727
rect 17635 10693 17644 10727
rect 17592 10684 17644 10693
rect 3424 10548 3476 10600
rect 15016 10616 15068 10668
rect 14648 10548 14700 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 16488 10616 16540 10668
rect 19708 10752 19760 10804
rect 22652 10752 22704 10804
rect 24216 10795 24268 10804
rect 24216 10761 24225 10795
rect 24225 10761 24259 10795
rect 24259 10761 24268 10795
rect 24216 10752 24268 10761
rect 26332 10795 26384 10804
rect 26332 10761 26341 10795
rect 26341 10761 26375 10795
rect 26375 10761 26384 10795
rect 26332 10752 26384 10761
rect 27068 10752 27120 10804
rect 28724 10752 28776 10804
rect 22284 10684 22336 10736
rect 23848 10684 23900 10736
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 19800 10616 19852 10668
rect 20260 10616 20312 10668
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 12532 10412 12584 10464
rect 15660 10480 15712 10532
rect 15936 10480 15988 10532
rect 17960 10548 18012 10600
rect 19156 10548 19208 10600
rect 21088 10548 21140 10600
rect 20628 10480 20680 10532
rect 12808 10412 12860 10464
rect 14740 10412 14792 10464
rect 16672 10412 16724 10464
rect 17500 10412 17552 10464
rect 17592 10412 17644 10464
rect 21272 10412 21324 10464
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 23940 10548 23992 10600
rect 26700 10616 26752 10668
rect 27344 10684 27396 10736
rect 29920 10752 29972 10804
rect 31116 10752 31168 10804
rect 29552 10684 29604 10736
rect 30288 10684 30340 10736
rect 31484 10684 31536 10736
rect 33324 10727 33376 10736
rect 33324 10693 33333 10727
rect 33333 10693 33367 10727
rect 33367 10693 33376 10727
rect 33324 10684 33376 10693
rect 36636 10684 36688 10736
rect 36820 10795 36872 10804
rect 36820 10761 36829 10795
rect 36829 10761 36863 10795
rect 36863 10761 36872 10795
rect 36820 10752 36872 10761
rect 37280 10684 37332 10736
rect 49240 10684 49292 10736
rect 26608 10548 26660 10600
rect 27344 10591 27396 10600
rect 27344 10557 27353 10591
rect 27353 10557 27387 10591
rect 27387 10557 27396 10591
rect 27344 10548 27396 10557
rect 29736 10616 29788 10668
rect 23572 10480 23624 10532
rect 24768 10480 24820 10532
rect 29460 10548 29512 10600
rect 29552 10591 29604 10600
rect 29552 10557 29561 10591
rect 29561 10557 29595 10591
rect 29595 10557 29604 10591
rect 29552 10548 29604 10557
rect 29828 10548 29880 10600
rect 30472 10591 30524 10600
rect 30472 10557 30481 10591
rect 30481 10557 30515 10591
rect 30515 10557 30524 10591
rect 30472 10548 30524 10557
rect 30656 10616 30708 10668
rect 35624 10659 35676 10668
rect 35624 10625 35633 10659
rect 35633 10625 35667 10659
rect 35667 10625 35676 10659
rect 35624 10616 35676 10625
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 32220 10548 32272 10600
rect 32312 10548 32364 10600
rect 34704 10548 34756 10600
rect 36360 10591 36412 10600
rect 36360 10557 36369 10591
rect 36369 10557 36403 10591
rect 36403 10557 36412 10591
rect 36360 10548 36412 10557
rect 47216 10616 47268 10668
rect 22100 10412 22152 10464
rect 26056 10455 26108 10464
rect 26056 10421 26065 10455
rect 26065 10421 26099 10455
rect 26099 10421 26108 10455
rect 26056 10412 26108 10421
rect 26700 10412 26752 10464
rect 27436 10412 27488 10464
rect 30748 10412 30800 10464
rect 31760 10412 31812 10464
rect 31852 10455 31904 10464
rect 31852 10421 31861 10455
rect 31861 10421 31895 10455
rect 31895 10421 31904 10455
rect 31852 10412 31904 10421
rect 32220 10412 32272 10464
rect 35624 10480 35676 10532
rect 36544 10480 36596 10532
rect 38936 10480 38988 10532
rect 46940 10480 46992 10532
rect 36912 10412 36964 10464
rect 38568 10412 38620 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 1308 10208 1360 10260
rect 5448 10208 5500 10260
rect 16028 10208 16080 10260
rect 16672 10251 16724 10260
rect 16672 10217 16681 10251
rect 16681 10217 16715 10251
rect 16715 10217 16724 10251
rect 16672 10208 16724 10217
rect 17224 10208 17276 10260
rect 18328 10208 18380 10260
rect 19156 10208 19208 10260
rect 20260 10251 20312 10260
rect 20260 10217 20269 10251
rect 20269 10217 20303 10251
rect 20303 10217 20312 10251
rect 20260 10208 20312 10217
rect 1308 10072 1360 10124
rect 14740 10140 14792 10192
rect 17316 10140 17368 10192
rect 17500 10140 17552 10192
rect 19800 10140 19852 10192
rect 16580 10072 16632 10124
rect 17868 10072 17920 10124
rect 18328 10072 18380 10124
rect 18604 10115 18656 10124
rect 18604 10081 18613 10115
rect 18613 10081 18647 10115
rect 18647 10081 18656 10115
rect 18604 10072 18656 10081
rect 19432 10072 19484 10124
rect 19616 10072 19668 10124
rect 3332 10004 3384 10056
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 13084 10047 13136 10056
rect 12440 10004 12492 10013
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 13544 10004 13596 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 18512 10004 18564 10056
rect 23756 10251 23808 10260
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 24308 10208 24360 10260
rect 26332 10208 26384 10260
rect 29092 10208 29144 10260
rect 29828 10208 29880 10260
rect 30380 10251 30432 10260
rect 30380 10217 30389 10251
rect 30389 10217 30423 10251
rect 30423 10217 30432 10251
rect 30380 10208 30432 10217
rect 32036 10208 32088 10260
rect 21088 10072 21140 10124
rect 26608 10140 26660 10192
rect 29000 10183 29052 10192
rect 29000 10149 29009 10183
rect 29009 10149 29043 10183
rect 29043 10149 29052 10183
rect 29000 10140 29052 10149
rect 29368 10183 29420 10192
rect 29368 10149 29377 10183
rect 29377 10149 29411 10183
rect 29411 10149 29420 10183
rect 29368 10140 29420 10149
rect 30012 10140 30064 10192
rect 26884 10072 26936 10124
rect 29552 10072 29604 10124
rect 30656 10072 30708 10124
rect 34428 10140 34480 10192
rect 32128 10115 32180 10124
rect 32128 10081 32137 10115
rect 32137 10081 32171 10115
rect 32171 10081 32180 10115
rect 32128 10072 32180 10081
rect 32220 10072 32272 10124
rect 32772 10072 32824 10124
rect 34704 10072 34756 10124
rect 35164 10115 35216 10124
rect 35164 10081 35173 10115
rect 35173 10081 35207 10115
rect 35207 10081 35216 10115
rect 35164 10072 35216 10081
rect 14464 9936 14516 9988
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 14740 9868 14792 9920
rect 15016 9868 15068 9920
rect 15844 9936 15896 9988
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 24032 10004 24084 10056
rect 30748 10004 30800 10056
rect 32496 10004 32548 10056
rect 33508 10004 33560 10056
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17224 9868 17276 9920
rect 19800 9936 19852 9988
rect 20444 9936 20496 9988
rect 21456 9868 21508 9920
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 36636 10251 36688 10260
rect 36636 10217 36645 10251
rect 36645 10217 36679 10251
rect 36679 10217 36688 10251
rect 36636 10208 36688 10217
rect 47124 10072 47176 10124
rect 49148 10115 49200 10124
rect 49148 10081 49157 10115
rect 49157 10081 49191 10115
rect 49191 10081 49200 10115
rect 49148 10072 49200 10081
rect 38936 10004 38988 10056
rect 22468 9979 22520 9988
rect 22468 9945 22477 9979
rect 22477 9945 22511 9979
rect 22511 9945 22520 9979
rect 22468 9936 22520 9945
rect 23848 9979 23900 9988
rect 23848 9945 23857 9979
rect 23857 9945 23891 9979
rect 23891 9945 23900 9979
rect 23848 9936 23900 9945
rect 23940 9868 23992 9920
rect 25044 9868 25096 9920
rect 26056 9936 26108 9988
rect 26700 9911 26752 9920
rect 26700 9877 26709 9911
rect 26709 9877 26743 9911
rect 26743 9877 26752 9911
rect 26700 9868 26752 9877
rect 27252 9979 27304 9988
rect 27252 9945 27261 9979
rect 27261 9945 27295 9979
rect 27295 9945 27304 9979
rect 27252 9936 27304 9945
rect 28540 9936 28592 9988
rect 28724 9936 28776 9988
rect 31944 9936 31996 9988
rect 32680 9936 32732 9988
rect 34244 9936 34296 9988
rect 35440 9936 35492 9988
rect 35716 9936 35768 9988
rect 45836 10004 45888 10056
rect 46112 10047 46164 10056
rect 46112 10013 46121 10047
rect 46121 10013 46155 10047
rect 46155 10013 46164 10047
rect 46112 10004 46164 10013
rect 46664 10004 46716 10056
rect 44364 9979 44416 9988
rect 44364 9945 44373 9979
rect 44373 9945 44407 9979
rect 44407 9945 44416 9979
rect 44364 9936 44416 9945
rect 46756 9936 46808 9988
rect 47308 9979 47360 9988
rect 47308 9945 47317 9979
rect 47317 9945 47351 9979
rect 47351 9945 47360 9979
rect 47308 9936 47360 9945
rect 32036 9868 32088 9920
rect 32404 9868 32456 9920
rect 36820 9868 36872 9920
rect 36912 9911 36964 9920
rect 36912 9877 36921 9911
rect 36921 9877 36955 9911
rect 36955 9877 36964 9911
rect 36912 9868 36964 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 16672 9664 16724 9716
rect 3792 9596 3844 9648
rect 12624 9596 12676 9648
rect 13728 9596 13780 9648
rect 14648 9596 14700 9648
rect 15200 9596 15252 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 2688 9528 2740 9580
rect 2228 9460 2280 9512
rect 12348 9528 12400 9580
rect 16028 9596 16080 9648
rect 16120 9596 16172 9648
rect 19708 9596 19760 9648
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 26056 9664 26108 9716
rect 26700 9664 26752 9716
rect 21548 9639 21600 9648
rect 21548 9605 21557 9639
rect 21557 9605 21591 9639
rect 21591 9605 21600 9639
rect 21548 9596 21600 9605
rect 22560 9596 22612 9648
rect 24676 9596 24728 9648
rect 15844 9528 15896 9580
rect 16488 9571 16540 9580
rect 16488 9537 16497 9571
rect 16497 9537 16531 9571
rect 16531 9537 16540 9571
rect 16488 9528 16540 9537
rect 17500 9528 17552 9580
rect 23388 9528 23440 9580
rect 23848 9528 23900 9580
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 11060 9460 11112 9512
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 17592 9460 17644 9512
rect 18604 9503 18656 9512
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 18880 9503 18932 9512
rect 18880 9469 18889 9503
rect 18889 9469 18923 9503
rect 18923 9469 18932 9503
rect 18880 9460 18932 9469
rect 19616 9503 19668 9512
rect 19616 9469 19625 9503
rect 19625 9469 19659 9503
rect 19659 9469 19668 9503
rect 19616 9460 19668 9469
rect 23756 9460 23808 9512
rect 24308 9460 24360 9512
rect 27252 9596 27304 9648
rect 28724 9664 28776 9716
rect 30196 9664 30248 9716
rect 31576 9664 31628 9716
rect 30104 9596 30156 9648
rect 30748 9596 30800 9648
rect 31484 9596 31536 9648
rect 31852 9664 31904 9716
rect 32036 9664 32088 9716
rect 32312 9664 32364 9716
rect 32496 9596 32548 9648
rect 34888 9664 34940 9716
rect 35164 9664 35216 9716
rect 35716 9664 35768 9716
rect 25964 9503 26016 9512
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 25780 9392 25832 9444
rect 31668 9528 31720 9580
rect 36084 9596 36136 9648
rect 36912 9664 36964 9716
rect 49332 9596 49384 9648
rect 47400 9528 47452 9580
rect 27160 9460 27212 9512
rect 29276 9503 29328 9512
rect 29276 9469 29285 9503
rect 29285 9469 29319 9503
rect 29319 9469 29328 9503
rect 29276 9460 29328 9469
rect 29552 9460 29604 9512
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 14924 9324 14976 9376
rect 16028 9367 16080 9376
rect 16028 9333 16037 9367
rect 16037 9333 16071 9367
rect 16071 9333 16080 9367
rect 16028 9324 16080 9333
rect 18788 9324 18840 9376
rect 19800 9324 19852 9376
rect 22008 9324 22060 9376
rect 22284 9367 22336 9376
rect 22284 9333 22293 9367
rect 22293 9333 22327 9367
rect 22327 9333 22336 9367
rect 22284 9324 22336 9333
rect 23756 9324 23808 9376
rect 28816 9324 28868 9376
rect 29276 9324 29328 9376
rect 29644 9392 29696 9444
rect 30104 9460 30156 9512
rect 31760 9503 31812 9512
rect 31760 9469 31769 9503
rect 31769 9469 31803 9503
rect 31803 9469 31812 9503
rect 31760 9460 31812 9469
rect 31944 9460 31996 9512
rect 32772 9460 32824 9512
rect 35900 9503 35952 9512
rect 35900 9469 35909 9503
rect 35909 9469 35943 9503
rect 35943 9469 35952 9503
rect 35900 9460 35952 9469
rect 32220 9392 32272 9444
rect 30472 9324 30524 9376
rect 31760 9324 31812 9376
rect 32588 9324 32640 9376
rect 33232 9324 33284 9376
rect 35532 9324 35584 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 2780 9120 2832 9172
rect 13820 9120 13872 9172
rect 15752 9120 15804 9172
rect 17132 9120 17184 9172
rect 17408 9120 17460 9172
rect 19616 9120 19668 9172
rect 22100 9120 22152 9172
rect 22468 9120 22520 9172
rect 25044 9120 25096 9172
rect 32404 9120 32456 9172
rect 32588 9120 32640 9172
rect 36360 9120 36412 9172
rect 43720 9120 43772 9172
rect 15844 9052 15896 9104
rect 16856 9052 16908 9104
rect 29644 9052 29696 9104
rect 1308 8916 1360 8968
rect 4068 8984 4120 9036
rect 12532 8984 12584 9036
rect 15108 8984 15160 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 16488 8984 16540 9036
rect 18880 8984 18932 9036
rect 19432 8984 19484 9036
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 24032 9027 24084 9036
rect 24032 8993 24041 9027
rect 24041 8993 24075 9027
rect 24075 8993 24084 9027
rect 24032 8984 24084 8993
rect 30196 8984 30248 9036
rect 31484 8984 31536 9036
rect 33324 9052 33376 9104
rect 35992 9052 36044 9104
rect 32496 9027 32548 9036
rect 32496 8993 32505 9027
rect 32505 8993 32539 9027
rect 32539 8993 32548 9027
rect 32496 8984 32548 8993
rect 32772 8984 32824 9036
rect 33048 8984 33100 9036
rect 34244 8984 34296 9036
rect 34980 9027 35032 9036
rect 34980 8993 34989 9027
rect 34989 8993 35023 9027
rect 35023 8993 35032 9027
rect 34980 8984 35032 8993
rect 35072 8984 35124 9036
rect 35532 8984 35584 9036
rect 1216 8848 1268 8900
rect 12164 8916 12216 8968
rect 15660 8916 15712 8968
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 19800 8916 19852 8968
rect 21456 8916 21508 8968
rect 25964 8916 26016 8968
rect 30932 8916 30984 8968
rect 33876 8916 33928 8968
rect 34520 8916 34572 8968
rect 2596 8780 2648 8832
rect 15292 8848 15344 8900
rect 16580 8848 16632 8900
rect 17868 8891 17920 8900
rect 17868 8857 17877 8891
rect 17877 8857 17911 8891
rect 17911 8857 17920 8891
rect 17868 8848 17920 8857
rect 22008 8848 22060 8900
rect 14648 8780 14700 8832
rect 31760 8848 31812 8900
rect 22192 8780 22244 8832
rect 23388 8780 23440 8832
rect 24860 8823 24912 8832
rect 24860 8789 24869 8823
rect 24869 8789 24903 8823
rect 24903 8789 24912 8823
rect 24860 8780 24912 8789
rect 25780 8823 25832 8832
rect 25780 8789 25789 8823
rect 25789 8789 25823 8823
rect 25823 8789 25832 8823
rect 25780 8780 25832 8789
rect 27804 8823 27856 8832
rect 27804 8789 27813 8823
rect 27813 8789 27847 8823
rect 27847 8789 27856 8823
rect 27804 8780 27856 8789
rect 30196 8780 30248 8832
rect 30748 8780 30800 8832
rect 32128 8780 32180 8832
rect 36452 8848 36504 8900
rect 49240 8984 49292 9036
rect 39396 8916 39448 8968
rect 46480 8916 46532 8968
rect 47032 8916 47084 8968
rect 47584 8848 47636 8900
rect 34244 8780 34296 8832
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 35624 8823 35676 8832
rect 35624 8789 35633 8823
rect 35633 8789 35667 8823
rect 35667 8789 35676 8823
rect 35624 8780 35676 8789
rect 37832 8823 37884 8832
rect 37832 8789 37841 8823
rect 37841 8789 37875 8823
rect 37875 8789 37884 8823
rect 37832 8780 37884 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 2596 8440 2648 8492
rect 2780 8440 2832 8492
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 12716 8576 12768 8628
rect 15200 8576 15252 8628
rect 17500 8576 17552 8628
rect 17868 8576 17920 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 19064 8619 19116 8628
rect 19064 8585 19073 8619
rect 19073 8585 19107 8619
rect 19107 8585 19116 8619
rect 19064 8576 19116 8585
rect 19892 8576 19944 8628
rect 14188 8508 14240 8560
rect 16580 8508 16632 8560
rect 16764 8508 16816 8560
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 19800 8508 19852 8560
rect 15200 8440 15252 8492
rect 16488 8440 16540 8492
rect 15108 8372 15160 8424
rect 16396 8415 16448 8424
rect 16396 8381 16405 8415
rect 16405 8381 16439 8415
rect 16439 8381 16448 8415
rect 16396 8372 16448 8381
rect 17224 8372 17276 8424
rect 21180 8372 21232 8424
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 16672 8304 16724 8356
rect 22008 8440 22060 8492
rect 30472 8576 30524 8628
rect 32128 8576 32180 8628
rect 32496 8576 32548 8628
rect 29092 8551 29144 8560
rect 29092 8517 29101 8551
rect 29101 8517 29135 8551
rect 29135 8517 29144 8551
rect 29092 8508 29144 8517
rect 30748 8508 30800 8560
rect 24032 8440 24084 8492
rect 22100 8372 22152 8424
rect 28816 8415 28868 8424
rect 28816 8381 28825 8415
rect 28825 8381 28859 8415
rect 28859 8381 28868 8415
rect 28816 8372 28868 8381
rect 32588 8508 32640 8560
rect 33324 8576 33376 8628
rect 34980 8576 35032 8628
rect 40040 8576 40092 8628
rect 33876 8508 33928 8560
rect 34336 8508 34388 8560
rect 31116 8440 31168 8492
rect 32312 8483 32364 8492
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 22468 8304 22520 8356
rect 24860 8304 24912 8356
rect 31852 8372 31904 8424
rect 32220 8372 32272 8424
rect 32956 8372 33008 8424
rect 33048 8372 33100 8424
rect 35624 8508 35676 8560
rect 36084 8440 36136 8492
rect 36820 8440 36872 8492
rect 37832 8508 37884 8560
rect 47768 8508 47820 8560
rect 49148 8551 49200 8560
rect 49148 8517 49157 8551
rect 49157 8517 49191 8551
rect 49191 8517 49200 8551
rect 49148 8508 49200 8517
rect 40316 8483 40368 8492
rect 40316 8449 40325 8483
rect 40325 8449 40359 8483
rect 40359 8449 40368 8483
rect 40316 8440 40368 8449
rect 45836 8483 45888 8492
rect 45836 8449 45845 8483
rect 45845 8449 45879 8483
rect 45879 8449 45888 8483
rect 45836 8440 45888 8449
rect 46756 8440 46808 8492
rect 39396 8372 39448 8424
rect 31944 8304 31996 8356
rect 32036 8236 32088 8288
rect 38752 8304 38804 8356
rect 44916 8304 44968 8356
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 47676 8304 47728 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 2780 8032 2832 8084
rect 18512 8032 18564 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 21916 8032 21968 8084
rect 30564 8032 30616 8084
rect 35256 8032 35308 8084
rect 18880 7964 18932 8016
rect 27528 7964 27580 8016
rect 3516 7896 3568 7948
rect 16396 7896 16448 7948
rect 16764 7939 16816 7948
rect 16764 7905 16773 7939
rect 16773 7905 16807 7939
rect 16807 7905 16816 7939
rect 16764 7896 16816 7905
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 18604 7896 18656 7948
rect 19892 7896 19944 7948
rect 23572 7896 23624 7948
rect 29920 7939 29972 7948
rect 29920 7905 29929 7939
rect 29929 7905 29963 7939
rect 29963 7905 29972 7939
rect 29920 7896 29972 7905
rect 32220 7896 32272 7948
rect 34612 7896 34664 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 2228 7828 2280 7880
rect 14924 7828 14976 7880
rect 18328 7828 18380 7880
rect 19800 7828 19852 7880
rect 14372 7760 14424 7812
rect 18420 7692 18472 7744
rect 19616 7760 19668 7812
rect 20996 7760 21048 7812
rect 21456 7828 21508 7880
rect 22192 7828 22244 7880
rect 30564 7828 30616 7880
rect 32680 7871 32732 7880
rect 32680 7837 32689 7871
rect 32689 7837 32723 7871
rect 32723 7837 32732 7871
rect 32680 7828 32732 7837
rect 49332 7896 49384 7948
rect 21272 7760 21324 7812
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 30748 7803 30800 7812
rect 30748 7769 30757 7803
rect 30757 7769 30791 7803
rect 30791 7769 30800 7803
rect 30748 7760 30800 7769
rect 31668 7760 31720 7812
rect 31760 7760 31812 7812
rect 39028 7828 39080 7880
rect 46940 7828 46992 7880
rect 25780 7692 25832 7744
rect 30472 7735 30524 7744
rect 30472 7701 30481 7735
rect 30481 7701 30515 7735
rect 30515 7701 30524 7735
rect 30472 7692 30524 7701
rect 31392 7735 31444 7744
rect 31392 7701 31401 7735
rect 31401 7701 31435 7735
rect 31435 7701 31444 7735
rect 31392 7692 31444 7701
rect 32588 7735 32640 7744
rect 32588 7701 32597 7735
rect 32597 7701 32631 7735
rect 32631 7701 32640 7735
rect 32588 7692 32640 7701
rect 38752 7803 38804 7812
rect 38752 7769 38761 7803
rect 38761 7769 38795 7803
rect 38795 7769 38804 7803
rect 38752 7760 38804 7769
rect 40592 7760 40644 7812
rect 38660 7692 38712 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 3608 7488 3660 7540
rect 21272 7488 21324 7540
rect 22284 7488 22336 7540
rect 31116 7531 31168 7540
rect 31116 7497 31125 7531
rect 31125 7497 31159 7531
rect 31159 7497 31168 7531
rect 31116 7488 31168 7497
rect 31392 7488 31444 7540
rect 1308 7352 1360 7404
rect 21180 7420 21232 7472
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 17960 7352 18012 7404
rect 19800 7352 19852 7404
rect 31852 7463 31904 7472
rect 31852 7429 31861 7463
rect 31861 7429 31895 7463
rect 31895 7429 31904 7463
rect 31852 7420 31904 7429
rect 32772 7420 32824 7472
rect 34428 7420 34480 7472
rect 38660 7420 38712 7472
rect 46940 7420 46992 7472
rect 49240 7420 49292 7472
rect 30472 7352 30524 7404
rect 21456 7284 21508 7336
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 20720 7216 20772 7268
rect 28632 7216 28684 7268
rect 44916 7395 44968 7404
rect 44916 7361 44925 7395
rect 44925 7361 44959 7395
rect 44959 7361 44968 7395
rect 44916 7352 44968 7361
rect 47124 7352 47176 7404
rect 2780 7148 2832 7200
rect 32588 7148 32640 7200
rect 37280 7148 37332 7200
rect 37924 7191 37976 7200
rect 37924 7157 37933 7191
rect 37933 7157 37967 7191
rect 37967 7157 37976 7191
rect 37924 7148 37976 7157
rect 47860 7216 47912 7268
rect 45744 7148 45796 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 30472 6944 30524 6996
rect 38476 6944 38528 6996
rect 37924 6876 37976 6928
rect 47032 6876 47084 6928
rect 49148 6851 49200 6860
rect 49148 6817 49157 6851
rect 49157 6817 49191 6851
rect 49191 6817 49200 6851
rect 49148 6808 49200 6817
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 1308 6672 1360 6724
rect 16856 6740 16908 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 40592 6740 40644 6792
rect 47768 6740 47820 6792
rect 2872 6647 2924 6656
rect 2872 6613 2881 6647
rect 2881 6613 2915 6647
rect 2915 6613 2924 6647
rect 2872 6604 2924 6613
rect 10600 6672 10652 6724
rect 48688 6672 48740 6724
rect 19248 6604 19300 6656
rect 21916 6604 21968 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 2780 6375 2832 6384
rect 2780 6341 2789 6375
rect 2789 6341 2823 6375
rect 2823 6341 2832 6375
rect 2780 6332 2832 6341
rect 27804 6332 27856 6384
rect 30840 6332 30892 6384
rect 40040 6332 40092 6384
rect 49332 6332 49384 6384
rect 1308 6264 1360 6316
rect 10968 6264 11020 6316
rect 23940 6264 23992 6316
rect 27068 6264 27120 6316
rect 36820 6264 36872 6316
rect 37004 6264 37056 6316
rect 47216 6264 47268 6316
rect 47584 6264 47636 6316
rect 15844 6196 15896 6248
rect 18328 6196 18380 6248
rect 26976 6196 27028 6248
rect 37740 6196 37792 6248
rect 11704 6128 11756 6180
rect 28356 6128 28408 6180
rect 39212 6128 39264 6180
rect 47124 6128 47176 6180
rect 2136 6060 2188 6112
rect 12440 6060 12492 6112
rect 19432 6060 19484 6112
rect 37648 6103 37700 6112
rect 37648 6069 37657 6103
rect 37657 6069 37691 6103
rect 37691 6069 37700 6103
rect 37648 6060 37700 6069
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 37648 5856 37700 5908
rect 47400 5856 47452 5908
rect 49240 5720 49292 5772
rect 1400 5652 1452 5704
rect 1308 5584 1360 5636
rect 43720 5695 43772 5704
rect 43720 5661 43729 5695
rect 43729 5661 43763 5695
rect 43763 5661 43772 5695
rect 43720 5652 43772 5661
rect 47676 5652 47728 5704
rect 3424 5584 3476 5636
rect 45652 5584 45704 5636
rect 2872 5516 2924 5568
rect 16028 5516 16080 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 3424 5355 3476 5364
rect 3424 5321 3433 5355
rect 3433 5321 3467 5355
rect 3467 5321 3476 5355
rect 3424 5312 3476 5321
rect 11888 5244 11940 5296
rect 37280 5244 37332 5296
rect 38476 5287 38528 5296
rect 38476 5253 38485 5287
rect 38485 5253 38519 5287
rect 38519 5253 38528 5287
rect 38476 5244 38528 5253
rect 49148 5287 49200 5296
rect 49148 5253 49157 5287
rect 49157 5253 49191 5287
rect 49191 5253 49200 5287
rect 49148 5244 49200 5253
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 45744 5176 45796 5228
rect 47860 5176 47912 5228
rect 1308 5108 1360 5160
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 48320 5108 48372 5160
rect 13360 5040 13412 5092
rect 40040 5040 40092 5092
rect 1400 4972 1452 5024
rect 20628 4972 20680 5024
rect 37832 5015 37884 5024
rect 37832 4981 37841 5015
rect 37841 4981 37875 5015
rect 37875 4981 37884 5015
rect 37832 4972 37884 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 3516 4768 3568 4820
rect 5540 4768 5592 4820
rect 23388 4768 23440 4820
rect 25780 4768 25832 4820
rect 36452 4768 36504 4820
rect 36820 4811 36872 4820
rect 36820 4777 36829 4811
rect 36829 4777 36863 4811
rect 36863 4777 36872 4811
rect 36820 4768 36872 4777
rect 37832 4768 37884 4820
rect 47308 4768 47360 4820
rect 19064 4700 19116 4752
rect 1308 4564 1360 4616
rect 19248 4632 19300 4684
rect 21916 4675 21968 4684
rect 21916 4641 21925 4675
rect 21925 4641 21959 4675
rect 21959 4641 21968 4675
rect 21916 4632 21968 4641
rect 26148 4700 26200 4752
rect 46480 4743 46532 4752
rect 46480 4709 46489 4743
rect 46489 4709 46523 4743
rect 46523 4709 46532 4743
rect 46480 4700 46532 4709
rect 47216 4743 47268 4752
rect 47216 4709 47225 4743
rect 47225 4709 47259 4743
rect 47259 4709 47268 4743
rect 47216 4700 47268 4709
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 19984 4564 20036 4616
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 23572 4632 23624 4684
rect 49424 4632 49476 4684
rect 23204 4564 23256 4616
rect 15844 4496 15896 4548
rect 36820 4564 36872 4616
rect 37740 4564 37792 4616
rect 46940 4564 46992 4616
rect 28724 4496 28776 4548
rect 39764 4496 39816 4548
rect 10968 4428 11020 4480
rect 21272 4428 21324 4480
rect 24768 4428 24820 4480
rect 37372 4471 37424 4480
rect 37372 4437 37381 4471
rect 37381 4437 37415 4471
rect 37415 4437 37424 4471
rect 37372 4428 37424 4437
rect 47676 4496 47728 4548
rect 49792 4428 49844 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 2688 4224 2740 4276
rect 37372 4224 37424 4276
rect 45836 4224 45888 4276
rect 1216 4088 1268 4140
rect 18328 4156 18380 4208
rect 1308 4020 1360 4072
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 22100 4156 22152 4208
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 1124 3952 1176 4004
rect 23204 4088 23256 4140
rect 24768 4156 24820 4208
rect 23296 4020 23348 4072
rect 24860 4020 24912 4072
rect 27804 4020 27856 4072
rect 27896 4063 27948 4072
rect 27896 4029 27905 4063
rect 27905 4029 27939 4063
rect 27939 4029 27948 4063
rect 27896 4020 27948 4029
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 13360 3884 13412 3936
rect 22836 3884 22888 3936
rect 36544 4088 36596 4140
rect 47032 4088 47084 4140
rect 49332 4088 49384 4140
rect 35072 4020 35124 4072
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 27528 3884 27580 3936
rect 47676 3927 47728 3936
rect 47676 3893 47685 3927
rect 47685 3893 47719 3927
rect 47719 3893 47728 3927
rect 47676 3884 47728 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 7472 3680 7524 3732
rect 5540 3612 5592 3664
rect 19984 3680 20036 3732
rect 23296 3680 23348 3732
rect 23572 3723 23624 3732
rect 23572 3689 23581 3723
rect 23581 3689 23615 3723
rect 23615 3689 23624 3723
rect 23572 3680 23624 3689
rect 25964 3680 26016 3732
rect 36544 3723 36596 3732
rect 36544 3689 36553 3723
rect 36553 3689 36587 3723
rect 36587 3689 36596 3723
rect 36544 3680 36596 3689
rect 1308 3544 1360 3596
rect 5356 3544 5408 3596
rect 15292 3544 15344 3596
rect 17684 3612 17736 3664
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 2688 3476 2740 3528
rect 10324 3476 10376 3528
rect 10416 3476 10468 3528
rect 15844 3476 15896 3528
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 22836 3476 22888 3528
rect 3332 3408 3384 3460
rect 18972 3408 19024 3460
rect 19340 3408 19392 3460
rect 23756 3476 23808 3528
rect 28356 3544 28408 3596
rect 33968 3544 34020 3596
rect 49148 3587 49200 3596
rect 49148 3553 49157 3587
rect 49157 3553 49191 3587
rect 49191 3553 49200 3587
rect 49148 3544 49200 3553
rect 26516 3476 26568 3528
rect 31760 3476 31812 3528
rect 36452 3519 36504 3528
rect 36452 3485 36461 3519
rect 36461 3485 36495 3519
rect 36495 3485 36504 3519
rect 36452 3476 36504 3485
rect 40040 3476 40092 3528
rect 47124 3476 47176 3528
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 10692 3340 10744 3392
rect 14832 3340 14884 3392
rect 22284 3340 22336 3392
rect 22744 3383 22796 3392
rect 22744 3349 22753 3383
rect 22753 3349 22787 3383
rect 22787 3349 22796 3383
rect 22744 3340 22796 3349
rect 29000 3408 29052 3460
rect 26516 3340 26568 3392
rect 28356 3340 28408 3392
rect 31300 3408 31352 3460
rect 45560 3451 45612 3460
rect 45560 3417 45569 3451
rect 45569 3417 45603 3451
rect 45603 3417 45612 3451
rect 45560 3408 45612 3417
rect 48688 3408 48740 3460
rect 29552 3383 29604 3392
rect 29552 3349 29561 3383
rect 29561 3349 29595 3383
rect 29595 3349 29604 3383
rect 29552 3340 29604 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 4068 3136 4120 3188
rect 10324 3179 10376 3188
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 1308 3000 1360 3052
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 9588 3000 9640 3052
rect 13360 3000 13412 3052
rect 15200 3136 15252 3188
rect 19340 3136 19392 3188
rect 14832 3111 14884 3120
rect 14832 3077 14841 3111
rect 14841 3077 14875 3111
rect 14875 3077 14884 3111
rect 14832 3068 14884 3077
rect 16580 3068 16632 3120
rect 19064 3068 19116 3120
rect 24584 3136 24636 3188
rect 25964 3179 26016 3188
rect 25964 3145 25973 3179
rect 25973 3145 26007 3179
rect 26007 3145 26016 3179
rect 25964 3136 26016 3145
rect 27528 3179 27580 3188
rect 27528 3145 27537 3179
rect 27537 3145 27571 3179
rect 27571 3145 27580 3179
rect 27528 3136 27580 3145
rect 27804 3136 27856 3188
rect 31300 3136 31352 3188
rect 31760 3111 31812 3120
rect 31760 3077 31769 3111
rect 31769 3077 31803 3111
rect 31803 3077 31812 3111
rect 31760 3068 31812 3077
rect 11704 2932 11756 2984
rect 14464 2932 14516 2984
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 3608 2864 3660 2916
rect 3884 2796 3936 2848
rect 9588 2796 9640 2848
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 20996 2932 21048 2984
rect 22100 2864 22152 2916
rect 22192 2907 22244 2916
rect 22192 2873 22201 2907
rect 22201 2873 22235 2907
rect 22235 2873 22244 2907
rect 22192 2864 22244 2873
rect 22744 2864 22796 2916
rect 26148 3000 26200 3052
rect 28356 3000 28408 3052
rect 28816 3000 28868 3052
rect 31392 3043 31444 3052
rect 31392 3009 31401 3043
rect 31401 3009 31435 3043
rect 31435 3009 31444 3043
rect 31392 3000 31444 3009
rect 33692 3000 33744 3052
rect 35256 3043 35308 3052
rect 35256 3009 35265 3043
rect 35265 3009 35299 3043
rect 35299 3009 35308 3043
rect 35256 3000 35308 3009
rect 49240 3068 49292 3120
rect 39764 3000 39816 3052
rect 45652 3000 45704 3052
rect 47400 3000 47452 3052
rect 26332 2932 26384 2984
rect 26516 2932 26568 2984
rect 28724 2932 28776 2984
rect 38292 2975 38344 2984
rect 38292 2941 38301 2975
rect 38301 2941 38335 2975
rect 38335 2941 38344 2975
rect 38292 2932 38344 2941
rect 46756 2932 46808 2984
rect 46848 2975 46900 2984
rect 46848 2941 46857 2975
rect 46857 2941 46891 2975
rect 46891 2941 46900 2975
rect 46848 2932 46900 2941
rect 22284 2796 22336 2848
rect 23296 2839 23348 2848
rect 23296 2805 23305 2839
rect 23305 2805 23339 2839
rect 23339 2805 23348 2839
rect 23296 2796 23348 2805
rect 27160 2796 27212 2848
rect 40684 2864 40736 2916
rect 35072 2839 35124 2848
rect 35072 2805 35081 2839
rect 35081 2805 35115 2839
rect 35115 2805 35124 2839
rect 35072 2796 35124 2805
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 2780 2592 2832 2644
rect 10416 2592 10468 2644
rect 26332 2635 26384 2644
rect 26332 2601 26341 2635
rect 26341 2601 26375 2635
rect 26375 2601 26384 2635
rect 26332 2592 26384 2601
rect 29000 2635 29052 2644
rect 29000 2601 29009 2635
rect 29009 2601 29043 2635
rect 29043 2601 29052 2635
rect 29000 2592 29052 2601
rect 31392 2592 31444 2644
rect 33692 2635 33744 2644
rect 33692 2601 33701 2635
rect 33701 2601 33735 2635
rect 33735 2601 33744 2635
rect 33692 2592 33744 2601
rect 35256 2592 35308 2644
rect 38292 2592 38344 2644
rect 12808 2524 12860 2576
rect 1216 2388 1268 2440
rect 3792 2456 3844 2508
rect 13820 2456 13872 2508
rect 15292 2499 15344 2508
rect 15292 2465 15301 2499
rect 15301 2465 15335 2499
rect 15335 2465 15344 2499
rect 15292 2456 15344 2465
rect 1308 2320 1360 2372
rect 4068 2388 4120 2440
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 14464 2388 14516 2440
rect 24860 2524 24912 2576
rect 34152 2524 34204 2576
rect 19984 2456 20036 2508
rect 20168 2456 20220 2508
rect 22284 2456 22336 2508
rect 24400 2456 24452 2508
rect 26516 2456 26568 2508
rect 29000 2456 29052 2508
rect 29552 2456 29604 2508
rect 3884 2320 3936 2372
rect 12072 2320 12124 2372
rect 15936 2320 15988 2372
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 22100 2388 22152 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 41328 2456 41380 2508
rect 49148 2499 49200 2508
rect 49148 2465 49157 2499
rect 49157 2465 49191 2499
rect 49191 2465 49200 2499
rect 49148 2456 49200 2465
rect 30748 2388 30800 2440
rect 40684 2431 40736 2440
rect 40684 2397 40693 2431
rect 40693 2397 40727 2431
rect 40727 2397 40736 2431
rect 40684 2388 40736 2397
rect 45836 2431 45888 2440
rect 45836 2397 45845 2431
rect 45845 2397 45879 2431
rect 45879 2397 45888 2431
rect 45836 2388 45888 2397
rect 47308 2388 47360 2440
rect 48504 2320 48556 2372
rect 32864 2252 32916 2304
rect 34980 2252 35032 2304
rect 37096 2295 37148 2304
rect 37096 2261 37105 2295
rect 37105 2261 37139 2295
rect 37139 2261 37148 2295
rect 37096 2252 37148 2261
rect 43444 2252 43496 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26330 2926 27000
rect 2870 26302 3372 26330
rect 2870 26200 2926 26302
rect 1596 22778 1624 26200
rect 1768 23044 1820 23050
rect 1768 22986 1820 22992
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1032 21956 1084 21962
rect 1032 21898 1084 21904
rect 1044 20777 1072 21898
rect 1780 21593 1808 22986
rect 2240 22234 2268 26200
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2778 24440 2834 24449
rect 2950 24443 3258 24452
rect 2778 24375 2834 24384
rect 2320 24132 2372 24138
rect 2320 24074 2372 24080
rect 2332 23866 2360 24074
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2792 23526 2820 24375
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2780 22500 2832 22506
rect 2780 22442 2832 22448
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 1766 21584 1822 21593
rect 1766 21519 1822 21528
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1030 20768 1086 20777
rect 1030 20703 1086 20712
rect 1308 20528 1360 20534
rect 1308 20470 1360 20476
rect 1320 20369 1348 20470
rect 1306 20360 1362 20369
rect 1306 20295 1362 20304
rect 1780 19961 1808 21422
rect 2792 21185 2820 22442
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3344 21622 3372 26302
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26200 4858 27000
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26330 8078 27000
rect 7852 26302 8078 26330
rect 3528 24274 3556 26200
rect 4066 25664 4122 25673
rect 4066 25599 4122 25608
rect 3698 25256 3754 25265
rect 4080 25226 4108 25599
rect 3698 25191 3754 25200
rect 4068 25220 4120 25226
rect 3606 24848 3662 24857
rect 3606 24783 3662 24792
rect 3620 24614 3648 24783
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3514 24032 3570 24041
rect 3514 23967 3570 23976
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2778 21176 2834 21185
rect 2950 21179 3258 21188
rect 2778 21111 2834 21120
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 1766 19952 1822 19961
rect 1766 19887 1822 19896
rect 1492 19780 1544 19786
rect 1492 19722 1544 19728
rect 1504 18737 1532 19722
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1490 18728 1546 18737
rect 1400 18692 1452 18698
rect 1490 18663 1546 18672
rect 1400 18634 1452 18640
rect 1412 17921 1440 18634
rect 1780 18329 1808 19314
rect 2792 19145 2820 20266
rect 2884 19553 2912 20946
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2870 19544 2926 19553
rect 2870 19479 2926 19488
rect 3436 19446 3464 22714
rect 3528 22098 3556 23967
rect 3608 23044 3660 23050
rect 3608 22986 3660 22992
rect 3516 22092 3568 22098
rect 3516 22034 3568 22040
rect 3514 21992 3570 22001
rect 3514 21927 3516 21936
rect 3568 21927 3570 21936
rect 3516 21898 3568 21904
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3620 18426 3648 22986
rect 3712 21622 3740 25191
rect 4068 25162 4120 25168
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3790 23216 3846 23225
rect 3790 23151 3846 23160
rect 3804 22438 3832 23151
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3700 21616 3752 21622
rect 3700 21558 3752 21564
rect 3804 18834 3832 22034
rect 3896 19310 3924 24142
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 3974 23624 4030 23633
rect 3974 23559 3976 23568
rect 4028 23559 4030 23568
rect 3976 23530 4028 23536
rect 3974 22808 4030 22817
rect 3974 22743 4030 22752
rect 3988 22166 4016 22743
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 1766 18320 1822 18329
rect 4080 18290 4108 23666
rect 4172 23662 4200 26200
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4724 23322 4752 23666
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4158 22536 4214 22545
rect 4158 22471 4214 22480
rect 4172 21010 4200 22471
rect 4252 22228 4304 22234
rect 4252 22170 4304 22176
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4264 19922 4292 22170
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 1766 18255 1822 18264
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 1032 17604 1084 17610
rect 1032 17546 1084 17552
rect 940 17128 992 17134
rect 1044 17105 1072 17546
rect 1780 17513 1808 18158
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3332 17808 3384 17814
rect 3332 17750 3384 17756
rect 1766 17504 1822 17513
rect 1766 17439 1822 17448
rect 940 17070 992 17076
rect 1030 17096 1086 17105
rect 952 16697 980 17070
rect 1030 17031 1086 17040
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 938 16688 994 16697
rect 938 16623 994 16632
rect 3344 16590 3372 17750
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 1032 16516 1084 16522
rect 1032 16458 1084 16464
rect 1044 16289 1072 16458
rect 1030 16280 1086 16289
rect 1030 16215 1086 16224
rect 4264 16114 4292 18158
rect 4356 17202 4384 18634
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4448 16658 4476 23054
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4632 21554 4660 22918
rect 4816 22710 4844 26200
rect 5460 23662 5488 26200
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5816 23588 5868 23594
rect 5816 23530 5868 23536
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 5356 22024 5408 22030
rect 5356 21966 5408 21972
rect 5368 21690 5396 21966
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4540 18358 4568 20198
rect 5276 19145 5304 20878
rect 5460 19854 5488 22918
rect 5644 21962 5672 23190
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5736 19922 5764 23462
rect 5828 21486 5856 23530
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 6012 22642 6040 23462
rect 6104 23186 6132 26200
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 6460 22500 6512 22506
rect 6460 22442 6512 22448
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 6012 21010 6040 22374
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6380 21010 6408 21490
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6472 20466 6500 22442
rect 6564 22094 6592 24550
rect 6748 24274 6776 26200
rect 6736 24268 6788 24274
rect 6736 24210 6788 24216
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6656 23118 6684 24006
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 7116 22574 7144 24142
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 6564 22066 6684 22094
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6564 20602 6592 21490
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6656 20398 6684 22066
rect 7208 20806 7236 22578
rect 7392 22574 7420 26200
rect 7470 24304 7526 24313
rect 7470 24239 7526 24248
rect 7484 24206 7512 24239
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 22642 7512 24006
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26200 10654 27000
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26330 12586 27000
rect 13174 26330 13230 27000
rect 12530 26302 12848 26330
rect 12530 26200 12586 26302
rect 8680 24274 8708 26200
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7840 23044 7892 23050
rect 7840 22986 7892 22992
rect 7564 22704 7616 22710
rect 7564 22646 7616 22652
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6380 19990 6408 20334
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5828 19174 5856 19314
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 5816 19168 5868 19174
rect 5262 19136 5318 19145
rect 5816 19110 5868 19116
rect 5262 19071 5318 19080
rect 4528 18352 4580 18358
rect 4528 18294 4580 18300
rect 5828 17202 5856 19110
rect 6840 18970 6868 19246
rect 7484 19242 7512 20742
rect 7576 19514 7604 22646
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 17338 7420 18566
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 1032 16040 1084 16046
rect 1032 15982 1084 15988
rect 1044 15881 1072 15982
rect 1030 15872 1086 15881
rect 1030 15807 1086 15816
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 938 15464 994 15473
rect 938 15399 940 15408
rect 992 15399 994 15408
rect 4160 15428 4212 15434
rect 940 15370 992 15376
rect 4160 15370 4212 15376
rect 938 15056 994 15065
rect 4172 15026 4200 15370
rect 938 14991 940 15000
rect 992 14991 994 15000
rect 4160 15020 4212 15026
rect 940 14962 992 14968
rect 4160 14962 4212 14968
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 938 14648 994 14657
rect 2950 14651 3258 14660
rect 938 14583 994 14592
rect 952 14482 980 14583
rect 940 14476 992 14482
rect 940 14418 992 14424
rect 1030 14240 1086 14249
rect 1030 14175 1086 14184
rect 1044 14006 1072 14175
rect 1032 14000 1084 14006
rect 1032 13942 1084 13948
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 1766 13832 1822 13841
rect 1766 13767 1822 13776
rect 1780 13394 1808 13767
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3528 13433 3556 13874
rect 3514 13424 3570 13433
rect 1768 13388 1820 13394
rect 3514 13359 3570 13368
rect 1768 13330 1820 13336
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 12918 1348 12951
rect 1308 12912 1360 12918
rect 1308 12854 1360 12860
rect 1308 12708 1360 12714
rect 1308 12650 1360 12656
rect 1320 12617 1348 12650
rect 2320 12640 2372 12646
rect 1306 12608 1362 12617
rect 2320 12582 2372 12588
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 1306 12543 1362 12552
rect 2228 12232 2280 12238
rect 1214 12200 1270 12209
rect 2228 12174 2280 12180
rect 1214 12135 1270 12144
rect 1228 11150 1256 12135
rect 2240 11898 2268 12174
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1306 11792 1362 11801
rect 2332 11762 2360 12582
rect 2884 12238 2912 12582
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 4264 11898 4292 16050
rect 4344 12436 4396 12442
rect 4448 12434 4476 16594
rect 4396 12406 4476 12434
rect 4344 12378 4396 12384
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 1306 11727 1308 11736
rect 1360 11727 1362 11736
rect 2320 11756 2372 11762
rect 1308 11698 1360 11704
rect 2320 11698 2372 11704
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 1306 11384 1362 11393
rect 1306 11319 1362 11328
rect 1320 11286 1348 11319
rect 2700 11286 2728 11698
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 1308 11280 1360 11286
rect 1308 11222 1360 11228
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 1216 11144 1268 11150
rect 1216 11086 1268 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 1306 10976 1362 10985
rect 1306 10911 1362 10920
rect 1320 10674 1348 10911
rect 2792 10810 2820 11086
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 1216 10600 1268 10606
rect 1216 10542 1268 10548
rect 1228 10169 1256 10542
rect 1320 10266 1348 10610
rect 3424 10600 3476 10606
rect 1582 10568 1638 10577
rect 3424 10542 3476 10548
rect 1582 10503 1638 10512
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1214 10160 1270 10169
rect 1214 10095 1270 10104
rect 1308 10124 1360 10130
rect 1308 10066 1360 10072
rect 1320 9761 1348 10066
rect 1306 9752 1362 9761
rect 1306 9687 1362 9696
rect 1596 9586 1624 10503
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 3344 10062 3372 10406
rect 3436 10062 3464 10542
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3804 9654 3832 10610
rect 5460 10266 5488 17002
rect 5828 12306 5856 17138
rect 7576 16590 7604 19450
rect 7668 18358 7696 21286
rect 7760 18766 7788 22374
rect 7852 21078 7880 22986
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8404 21894 8432 23598
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 8312 20754 8340 21830
rect 8392 20936 8444 20942
rect 8390 20904 8392 20913
rect 8444 20904 8446 20913
rect 8496 20874 8524 21898
rect 8588 20942 8616 23666
rect 9140 23118 9168 24006
rect 9220 23656 9272 23662
rect 9324 23644 9352 26200
rect 9772 25220 9824 25226
rect 9772 25162 9824 25168
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9272 23616 9352 23644
rect 9220 23598 9272 23604
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 22030 9168 22442
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9600 21690 9628 24074
rect 9784 22098 9812 25162
rect 9864 24336 9916 24342
rect 9864 24278 9916 24284
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8390 20839 8446 20848
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8312 20726 8432 20754
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 19174 8340 20470
rect 8404 20398 8432 20726
rect 9692 20602 9720 22034
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16250 8340 19110
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9048 16454 9076 16594
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 9048 16046 9076 16390
rect 9232 16250 9260 19382
rect 9784 18086 9812 20402
rect 9876 18426 9904 24278
rect 9968 22710 9996 26200
rect 10612 23662 10640 26200
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10324 23588 10376 23594
rect 10324 23530 10376 23536
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9968 19718 9996 20946
rect 10336 20602 10364 23530
rect 11164 22642 11192 24006
rect 11256 23186 11284 26200
rect 11900 24342 11928 26200
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23798 11836 24006
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 11978 23216 12034 23225
rect 11244 23180 11296 23186
rect 11978 23151 12034 23160
rect 11244 23122 11296 23128
rect 11888 23112 11940 23118
rect 11334 23080 11390 23089
rect 11888 23054 11940 23060
rect 11334 23015 11390 23024
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10428 20466 10456 21014
rect 11348 20942 11376 23015
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11440 21962 11468 22578
rect 11900 22234 11928 23054
rect 11992 22438 12020 23151
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11992 22098 12020 22374
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11440 21486 11468 21898
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10152 19854 10180 20266
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10612 19718 10640 20742
rect 11072 20602 11100 20742
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11164 20398 11192 20878
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11060 20392 11112 20398
rect 11058 20360 11060 20369
rect 11152 20392 11204 20398
rect 11112 20360 11114 20369
rect 11152 20334 11204 20340
rect 11058 20295 11114 20304
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10784 19848 10836 19854
rect 10782 19816 10784 19825
rect 10836 19816 10838 19825
rect 10782 19751 10838 19760
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9508 16658 9536 17070
rect 9692 16674 9720 18022
rect 9968 17202 9996 19654
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10244 17882 10272 18634
rect 10428 18426 10456 19246
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10612 17882 10640 18158
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10598 17776 10654 17785
rect 10598 17711 10654 17720
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10336 17270 10364 17478
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9876 16726 9904 17138
rect 10428 16794 10456 17614
rect 10612 17134 10640 17711
rect 10600 17128 10652 17134
rect 10520 17088 10600 17116
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 9864 16720 9916 16726
rect 9496 16652 9548 16658
rect 9692 16646 9812 16674
rect 9864 16662 9916 16668
rect 10520 16658 10548 17088
rect 10600 17070 10652 17076
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 9496 16594 9548 16600
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9048 15366 9076 15982
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 9048 13258 9076 15302
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 9508 12986 9536 16594
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9692 15162 9720 16458
rect 9784 16250 9812 16646
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15162 9812 15914
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9784 13802 9812 14894
rect 9876 14074 9904 15846
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10244 14550 10272 15438
rect 10520 15337 10548 16458
rect 10612 15910 10640 16662
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10704 15706 10732 18634
rect 10796 15978 10824 19654
rect 10980 16266 11008 19858
rect 11072 19281 11100 20198
rect 11058 19272 11114 19281
rect 11058 19207 11114 19216
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11164 16658 11192 18906
rect 11256 18902 11284 20742
rect 11532 20618 11560 21626
rect 11624 21457 11652 21966
rect 11610 21448 11666 21457
rect 11610 21383 11666 21392
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11532 20590 11652 20618
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11426 19952 11482 19961
rect 11426 19887 11482 19896
rect 11440 19786 11468 19887
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11532 18970 11560 20402
rect 11624 20262 11652 20590
rect 11716 20466 11744 21286
rect 11808 20942 11836 21354
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 11992 21078 12020 21286
rect 12176 21078 12204 23666
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12268 21554 12296 22374
rect 12360 22080 12388 24210
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12636 22778 12664 23598
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12820 22710 12848 26302
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 23186 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26200 16450 27000
rect 17038 26200 17094 27000
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26330 24178 27000
rect 24122 26302 24348 26330
rect 24122 26200 24178 26302
rect 13832 24274 13860 26200
rect 14476 24290 14504 26200
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 14384 24262 14504 24290
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 12808 22704 12860 22710
rect 13556 22681 13584 22714
rect 12808 22646 12860 22652
rect 13542 22672 13598 22681
rect 13542 22607 13598 22616
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12452 22080 12664 22094
rect 12360 22066 12664 22080
rect 12360 22052 12480 22066
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 11980 21072 12032 21078
rect 11980 21014 12032 21020
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 11808 20777 11836 20878
rect 11794 20768 11850 20777
rect 11794 20703 11850 20712
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11886 20360 11942 20369
rect 11886 20295 11942 20304
rect 11900 20262 11928 20295
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11520 18964 11572 18970
rect 11520 18906 11572 18912
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 10980 16250 11100 16266
rect 11348 16250 11376 16390
rect 10980 16244 11112 16250
rect 10980 16238 11060 16244
rect 11060 16186 11112 16192
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10506 15328 10562 15337
rect 10506 15263 10562 15272
rect 10888 15094 10916 16118
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 16017 11100 16050
rect 11058 16008 11114 16017
rect 11058 15943 11114 15952
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11072 15094 11100 15506
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11256 15162 11284 15302
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10704 14822 10732 14962
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 9968 14249 9996 14282
rect 9954 14240 10010 14249
rect 9954 14175 10010 14184
rect 9968 14074 9996 14175
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10428 13818 10456 14282
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 14006 10548 14214
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10508 13864 10560 13870
rect 10506 13832 10508 13841
rect 10560 13832 10562 13841
rect 9772 13796 9824 13802
rect 10428 13790 10506 13818
rect 10506 13767 10562 13776
rect 9772 13738 9824 13744
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 9784 12170 9812 13738
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1320 8974 1348 9279
rect 2240 9178 2268 9454
rect 2700 9178 2728 9522
rect 3700 9512 3752 9518
rect 3698 9480 3700 9489
rect 3752 9480 3754 9489
rect 3698 9415 3754 9424
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 9178 2820 9318
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 1308 8968 1360 8974
rect 1308 8910 1360 8916
rect 1582 8936 1638 8945
rect 1216 8900 1268 8906
rect 1582 8871 1638 8880
rect 1216 8842 1268 8848
rect 1228 8537 1256 8842
rect 1214 8528 1270 8537
rect 1214 8463 1270 8472
rect 1596 7886 1624 8871
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8498 2636 8774
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2424 8129 2452 8366
rect 2410 8120 2466 8129
rect 2792 8090 2820 8434
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2410 8055 2466 8064
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1320 7410 1348 7647
rect 2240 7546 2268 7822
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 1582 7304 1638 7313
rect 1582 7239 1638 7248
rect 1596 6798 1624 7239
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1320 6497 1348 6666
rect 1306 6488 1362 6497
rect 1306 6423 1362 6432
rect 2792 6390 2820 7142
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3344 6905 3372 7346
rect 3330 6896 3386 6905
rect 3330 6831 3386 6840
rect 2870 6760 2926 6769
rect 2870 6695 2926 6704
rect 2884 6662 2912 6695
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 2136 6112 2188 6118
rect 1306 6080 1362 6089
rect 2136 6054 2188 6060
rect 1306 6015 1362 6024
rect 1400 5704 1452 5710
rect 1306 5672 1362 5681
rect 1400 5646 1452 5652
rect 1306 5607 1308 5616
rect 1360 5607 1362 5616
rect 1308 5578 1360 5584
rect 1412 5273 1440 5646
rect 1398 5264 1454 5273
rect 1398 5199 1454 5208
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4865 1348 5102
rect 1412 5030 1440 5199
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1320 4457 1348 4558
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 1124 4004 1176 4010
rect 1124 3946 1176 3952
rect 1136 800 1164 3946
rect 1228 3641 1256 4082
rect 1308 4072 1360 4078
rect 1306 4040 1308 4049
rect 1360 4040 1362 4049
rect 1306 3975 1362 3984
rect 1214 3632 1270 3641
rect 1214 3567 1270 3576
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 1320 3233 1348 3538
rect 2148 3534 2176 6054
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5234 2912 5510
rect 3436 5370 3464 5578
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3528 4826 3556 7890
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 4282 2728 4558
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3534 2728 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 1306 3224 1362 3233
rect 1306 3159 1362 3168
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 1320 2825 1348 2994
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 2792 2650 2820 2994
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 1216 2440 1268 2446
rect 1216 2382 1268 2388
rect 1306 2408 1362 2417
rect 1228 2009 1256 2382
rect 1306 2343 1308 2352
rect 1360 2343 1362 2352
rect 1308 2314 1360 2320
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 3344 1714 3372 3402
rect 3620 2922 3648 7482
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3804 2514 3832 3334
rect 4080 3194 4108 8978
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 10704 6914 10732 14758
rect 11440 14618 11468 18294
rect 11624 16289 11652 19314
rect 11716 18222 11744 19722
rect 11980 19236 12032 19242
rect 11980 19178 12032 19184
rect 11888 19168 11940 19174
rect 11992 19145 12020 19178
rect 11888 19110 11940 19116
rect 11978 19136 12034 19145
rect 11900 18902 11928 19110
rect 11978 19071 12034 19080
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 17626 11744 18022
rect 11716 17610 11836 17626
rect 11716 17604 11848 17610
rect 11716 17598 11796 17604
rect 11796 17546 11848 17552
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11808 16658 11836 17002
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11610 16280 11666 16289
rect 11610 16215 11666 16224
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15473 11560 15846
rect 11518 15464 11574 15473
rect 11518 15399 11574 15408
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11242 14512 11298 14521
rect 11242 14447 11298 14456
rect 11256 14414 11284 14447
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11256 14074 11284 14350
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10796 13394 10824 13738
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10796 12306 10824 13330
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11072 12374 11100 13194
rect 11334 13152 11390 13161
rect 11334 13087 11390 13096
rect 11348 12986 11376 13087
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11072 11218 11100 12106
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11256 11286 11284 11766
rect 11428 11348 11480 11354
rect 11532 11336 11560 15399
rect 11900 15162 11928 18226
rect 11992 18222 12020 18566
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11992 17542 12020 18158
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11992 16794 12020 17206
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11808 15042 11836 15098
rect 11992 15042 12020 16526
rect 11808 15014 12020 15042
rect 11900 14074 11928 15014
rect 12084 14890 12112 17546
rect 12176 16590 12204 20878
rect 12268 19802 12296 21490
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12360 20874 12388 21354
rect 12452 21146 12480 21422
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 12360 19922 12388 20810
rect 12438 20496 12494 20505
rect 12438 20431 12440 20440
rect 12492 20431 12494 20440
rect 12440 20402 12492 20408
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12268 19774 12388 19802
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12268 18766 12296 19382
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12360 18465 12388 19774
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12452 18834 12480 19450
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12346 18456 12402 18465
rect 12452 18426 12480 18634
rect 12346 18391 12402 18400
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12544 17882 12572 21966
rect 12636 21690 12664 22066
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12636 19310 12664 21490
rect 12728 20369 12756 21898
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12820 21026 12848 21558
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12898 21040 12954 21049
rect 12820 20998 12898 21026
rect 13372 21010 13400 21830
rect 12898 20975 12954 20984
rect 13360 21004 13412 21010
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12714 20360 12770 20369
rect 12714 20295 12770 20304
rect 12624 19304 12676 19310
rect 12820 19258 12848 20810
rect 12912 20466 12940 20975
rect 13360 20946 13412 20952
rect 13648 20534 13676 24142
rect 13740 22030 13768 24142
rect 14384 23798 14412 24262
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13924 21690 13952 23054
rect 14188 22976 14240 22982
rect 14188 22918 14240 22924
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14200 22778 14228 22918
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14384 22438 14412 22918
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14384 22166 14412 22374
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 20806 13768 21286
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13636 20528 13688 20534
rect 13636 20470 13688 20476
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19854 13400 20402
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 19922 13492 20198
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13360 19848 13412 19854
rect 13188 19808 13360 19836
rect 13188 19446 13216 19808
rect 13360 19790 13412 19796
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12624 19246 12676 19252
rect 12728 19230 12848 19258
rect 12912 19258 12940 19314
rect 12912 19230 13400 19258
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12452 17338 12480 17818
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16794 12296 16934
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11716 12918 11744 13126
rect 11992 12986 12020 14826
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11612 12232 11664 12238
rect 11716 12220 11744 12854
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 12442 11836 12718
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11664 12192 11744 12220
rect 11612 12174 11664 12180
rect 11716 11898 11744 12192
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11480 11308 11560 11336
rect 11428 11290 11480 11296
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 9518 11100 11154
rect 11716 11098 11744 11834
rect 11808 11694 11836 12378
rect 12084 11898 12112 13670
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11218 11836 11630
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11716 11082 11836 11098
rect 11716 11076 11848 11082
rect 11716 11070 11796 11076
rect 11796 11018 11848 11024
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10612 6886 10732 6914
rect 10612 6730 10640 6886
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5552 3670 5580 4762
rect 10980 4486 11008 6258
rect 11716 6186 11744 10950
rect 11808 10810 11836 11018
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 11900 5302 11928 11494
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 10470 12112 10610
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3896 2378 3924 2790
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 3252 1686 3372 1714
rect 3252 800 3280 1686
rect 4080 1601 4108 2382
rect 4066 1592 4122 1601
rect 4066 1527 4122 1536
rect 5368 800 5396 3538
rect 7484 800 7512 3674
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 10336 3194 10364 3470
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9600 2854 9628 2994
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9600 800 9628 2790
rect 10428 2650 10456 3470
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10704 2446 10732 3334
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 11716 800 11744 2926
rect 12084 2378 12112 10406
rect 12176 8974 12204 16390
rect 12268 12753 12296 16526
rect 12360 15609 12388 17070
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12452 15706 12480 15982
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12346 15600 12402 15609
rect 12544 15570 12572 17682
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12346 15535 12402 15544
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12636 15434 12664 16594
rect 12728 16454 12756 19230
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18748 12848 19110
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18902 13400 19230
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13084 18828 13136 18834
rect 13004 18788 13084 18816
rect 13004 18748 13032 18788
rect 13084 18770 13136 18776
rect 12820 18720 13032 18748
rect 13096 18358 13124 18770
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13464 18290 13492 19450
rect 13556 18358 13584 20470
rect 13740 20466 13768 20742
rect 13818 20496 13874 20505
rect 13728 20460 13780 20466
rect 13818 20431 13820 20440
rect 13728 20402 13780 20408
rect 13872 20431 13874 20440
rect 13820 20402 13872 20408
rect 13634 20224 13690 20233
rect 13634 20159 13690 20168
rect 13648 18970 13676 20159
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13464 17746 13492 18226
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13556 17542 13584 18022
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12438 15328 12494 15337
rect 12438 15263 12494 15272
rect 12346 15056 12402 15065
rect 12346 14991 12348 15000
rect 12400 14991 12402 15000
rect 12348 14962 12400 14968
rect 12452 13410 12480 15263
rect 12820 14618 12848 16458
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13004 15366 13032 15642
rect 13266 15600 13322 15609
rect 13266 15535 13322 15544
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 15162 13032 15302
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13280 14804 13308 15535
rect 13372 15434 13400 16934
rect 13556 16572 13584 17478
rect 13648 17270 13676 18906
rect 13740 18154 13768 19246
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18970 13860 19110
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13832 18329 13860 18906
rect 13818 18320 13874 18329
rect 13818 18255 13874 18264
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16794 13768 16934
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13832 16590 13860 18255
rect 13924 17066 13952 21490
rect 14016 21418 14044 21626
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 14292 21146 14320 21558
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14292 20398 14320 21082
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14476 20058 14504 24142
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14568 21486 14596 22714
rect 14660 22642 14688 22918
rect 15120 22710 15148 26200
rect 15568 24132 15620 24138
rect 15568 24074 15620 24080
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14568 21010 14596 21422
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14568 18834 14596 19246
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14568 18222 14596 18634
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14568 17882 14596 18158
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14278 17640 14334 17649
rect 14004 17604 14056 17610
rect 14278 17575 14334 17584
rect 14004 17546 14056 17552
rect 13912 17060 13964 17066
rect 13912 17002 13964 17008
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13924 16658 13952 16730
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13820 16584 13872 16590
rect 13556 16544 13676 16572
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 16130 13492 16390
rect 13464 16102 13584 16130
rect 13556 16046 13584 16102
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13280 14776 13400 14804
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12360 13382 12480 13410
rect 12544 13394 12572 13806
rect 12532 13388 12584 13394
rect 12254 12744 12310 12753
rect 12254 12679 12310 12688
rect 12360 12050 12388 13382
rect 12532 13330 12584 13336
rect 12728 13172 12756 14214
rect 12820 13394 12848 14282
rect 13280 14006 13308 14418
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13280 13818 13308 13942
rect 13372 13920 13400 14776
rect 13464 14482 13492 15982
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13372 13892 13492 13920
rect 13280 13790 13400 13818
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12728 13144 12848 13172
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12360 12022 12480 12050
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 9586 12388 11494
rect 12452 11354 12480 12022
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12544 11014 12572 12922
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12452 6118 12480 9998
rect 12544 9042 12572 10406
rect 12636 9654 12664 12582
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12728 8634 12756 11086
rect 12820 10810 12848 13144
rect 12898 13016 12954 13025
rect 12898 12951 12900 12960
rect 12952 12951 12954 12960
rect 13268 12980 13320 12986
rect 12900 12922 12952 12928
rect 13372 12968 13400 13790
rect 13464 13530 13492 13892
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13320 12940 13400 12968
rect 13268 12922 13320 12928
rect 13464 12900 13492 13466
rect 13372 12872 13492 12900
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12374 13400 12872
rect 13556 12866 13584 15302
rect 13648 14958 13676 16544
rect 13820 16526 13872 16532
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13740 15638 13768 15982
rect 13924 15638 13952 16050
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13912 15632 13964 15638
rect 13912 15574 13964 15580
rect 13740 15450 13768 15574
rect 13740 15422 13952 15450
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 12986 13676 13670
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13556 12838 13676 12866
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13556 12170 13584 12378
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13358 12064 13414 12073
rect 13004 11762 13032 12038
rect 13358 11999 13414 12008
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13372 11558 13400 11999
rect 13556 11898 13584 12106
rect 13648 11898 13676 12838
rect 13740 12442 13768 13126
rect 13832 12782 13860 15302
rect 13924 15162 13952 15422
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14016 14793 14044 17546
rect 14292 17270 14320 17575
rect 14280 17264 14332 17270
rect 14186 17232 14242 17241
rect 14280 17206 14332 17212
rect 14186 17167 14188 17176
rect 14240 17167 14242 17176
rect 14188 17138 14240 17144
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 16153 14228 16594
rect 14660 16522 14688 21898
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15198 21584 15254 21593
rect 15198 21519 15254 21528
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15016 20052 15068 20058
rect 14936 20012 15016 20040
rect 14936 18222 14964 20012
rect 15016 19994 15068 20000
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15028 18834 15056 19110
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 15028 18290 15056 18770
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14936 16794 14964 18158
rect 15028 17610 15056 18226
rect 15120 17882 15148 20402
rect 15212 19786 15240 21519
rect 15304 21486 15332 21830
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15396 19514 15424 22442
rect 15580 20602 15608 24074
rect 15764 23186 15792 26200
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15856 20602 15884 23190
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15658 19816 15714 19825
rect 15948 19802 15976 21286
rect 16040 20602 16068 24754
rect 16408 23662 16436 26200
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16224 21962 16252 22374
rect 17052 22166 17080 26200
rect 17696 24274 17724 26200
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17236 23594 17264 24074
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23662 18368 26200
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18892 24206 18920 24686
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17224 23588 17276 23594
rect 17224 23530 17276 23536
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 17144 22234 17172 22510
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17040 22160 17092 22166
rect 17040 22102 17092 22108
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16224 21622 16252 21898
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15658 19751 15714 19760
rect 15856 19774 15976 19802
rect 15672 19718 15700 19751
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15488 19514 15516 19654
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15198 19272 15254 19281
rect 15198 19207 15200 19216
rect 15252 19207 15254 19216
rect 15200 19178 15252 19184
rect 15660 18760 15712 18766
rect 15658 18728 15660 18737
rect 15712 18728 15714 18737
rect 15856 18714 15884 19774
rect 16132 19514 16160 20810
rect 16224 20806 16252 21558
rect 16580 21344 16632 21350
rect 16684 21332 16712 21898
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16632 21304 16712 21332
rect 16580 21286 16632 21292
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16028 19440 16080 19446
rect 15934 19408 15990 19417
rect 16028 19382 16080 19388
rect 15934 19343 15936 19352
rect 15988 19343 15990 19352
rect 15936 19314 15988 19320
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15948 18970 15976 19110
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15856 18686 15976 18714
rect 15658 18663 15714 18672
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15292 18080 15344 18086
rect 15344 18040 15424 18068
rect 15292 18022 15344 18028
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14186 16144 14242 16153
rect 14108 16102 14186 16130
rect 14002 14784 14058 14793
rect 14002 14719 14058 14728
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12820 2582 12848 10406
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13082 10160 13138 10169
rect 13082 10095 13138 10104
rect 13096 10062 13124 10095
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13372 5098 13400 11494
rect 13556 11354 13584 11834
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13464 10849 13492 11018
rect 13450 10840 13506 10849
rect 13450 10775 13506 10784
rect 13556 10062 13584 11290
rect 13634 10704 13690 10713
rect 13634 10639 13636 10648
rect 13688 10639 13690 10648
rect 13636 10610 13688 10616
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13740 9654 13768 12242
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13832 9178 13860 12582
rect 13924 11354 13952 14214
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14016 13297 14044 13466
rect 14108 13433 14136 16102
rect 14186 16079 14242 16088
rect 14292 16102 14504 16130
rect 14752 16114 14780 16662
rect 14936 16454 14964 16730
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14292 15978 14320 16102
rect 14476 15978 14504 16102
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14384 15094 14412 15642
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14414 14320 14894
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14476 14226 14504 15506
rect 14660 15473 14688 15982
rect 14646 15464 14702 15473
rect 14646 15399 14702 15408
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 14618 14596 15302
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14200 14198 14504 14226
rect 14094 13424 14150 13433
rect 14094 13359 14150 13368
rect 14002 13288 14058 13297
rect 14002 13223 14058 13232
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14016 12918 14044 13126
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 14108 12646 14136 13126
rect 14200 12646 14228 14198
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14096 12640 14148 12646
rect 14002 12608 14058 12617
rect 14096 12582 14148 12588
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14002 12543 14058 12552
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14016 10742 14044 12543
rect 14200 12442 14228 12582
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14292 11898 14320 14010
rect 14476 13802 14504 14198
rect 14660 13938 14688 15399
rect 14752 14958 14780 16050
rect 15028 15722 15056 17546
rect 15396 17202 15424 18040
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15120 16697 15148 17138
rect 15106 16688 15162 16697
rect 15106 16623 15162 16632
rect 14936 15706 15056 15722
rect 14924 15700 15056 15706
rect 14976 15694 15056 15700
rect 14924 15642 14976 15648
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14740 14952 14792 14958
rect 14738 14920 14740 14929
rect 14792 14920 14794 14929
rect 14738 14855 14794 14864
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14462 13424 14518 13433
rect 14462 13359 14518 13368
rect 14476 13326 14504 13359
rect 14464 13320 14516 13326
rect 14370 13288 14426 13297
rect 14464 13262 14516 13268
rect 14370 13223 14426 13232
rect 14384 12102 14412 13223
rect 14476 13161 14504 13262
rect 14462 13152 14518 13161
rect 14462 13087 14518 13096
rect 14752 13002 14780 14855
rect 14844 13394 14872 15506
rect 14936 14396 14964 15642
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 15028 15162 15056 15574
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 15120 15026 15148 15438
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15200 14952 15252 14958
rect 15120 14900 15200 14906
rect 15120 14894 15252 14900
rect 15120 14878 15240 14894
rect 15120 14498 15148 14878
rect 15120 14482 15240 14498
rect 15120 14476 15252 14482
rect 15120 14470 15200 14476
rect 14936 14368 15056 14396
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 13530 14964 14214
rect 15028 14006 15056 14368
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14476 12974 14780 13002
rect 14476 12170 14504 12974
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14568 12434 14596 12854
rect 14844 12458 14872 13330
rect 14924 13320 14976 13326
rect 15028 13297 15056 13942
rect 14924 13262 14976 13268
rect 15014 13288 15070 13297
rect 14936 12617 14964 13262
rect 15014 13223 15016 13232
rect 15068 13223 15070 13232
rect 15016 13194 15068 13200
rect 15016 12640 15068 12646
rect 14922 12608 14978 12617
rect 15016 12582 15068 12588
rect 14922 12543 14978 12552
rect 14568 12406 14688 12434
rect 14844 12430 14964 12458
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14660 11898 14688 12406
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14292 10577 14320 11630
rect 14384 10810 14412 11766
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14278 10568 14334 10577
rect 14278 10503 14334 10512
rect 14292 9926 14320 10503
rect 14476 9994 14504 11290
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 9674 14320 9862
rect 14200 9646 14320 9674
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14200 8566 14228 9646
rect 14370 8936 14426 8945
rect 14370 8871 14426 8880
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14384 7818 14412 8871
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 14568 4078 14596 11630
rect 14660 10606 14688 11834
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11218 14780 11698
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11218 14872 11494
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14740 11076 14792 11082
rect 14740 11018 14792 11024
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14752 10470 14780 11018
rect 14936 10606 14964 12430
rect 15028 10674 15056 12582
rect 15120 11218 15148 14470
rect 15200 14418 15252 14424
rect 15198 13016 15254 13025
rect 15198 12951 15200 12960
rect 15252 12951 15254 12960
rect 15200 12922 15252 12928
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15304 12306 15332 12650
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15396 11830 15424 17138
rect 15580 17066 15608 18566
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15856 16998 15884 18566
rect 15948 18154 15976 18686
rect 15936 18148 15988 18154
rect 15936 18090 15988 18096
rect 16040 17746 16068 19382
rect 16132 19242 16160 19450
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15856 16658 15884 16934
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15488 13394 15516 16390
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15580 13326 15608 15302
rect 15672 15094 15700 16390
rect 15764 16046 15792 16526
rect 15948 16250 15976 16934
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15842 16144 15898 16153
rect 15842 16079 15844 16088
rect 15896 16079 15898 16088
rect 15844 16050 15896 16056
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15764 15570 15792 15982
rect 15752 15564 15804 15570
rect 15804 15524 15884 15552
rect 15752 15506 15804 15512
rect 15750 15464 15806 15473
rect 15750 15399 15806 15408
rect 15764 15366 15792 15399
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15672 13172 15700 14010
rect 15856 13546 15884 15524
rect 15948 15502 15976 16186
rect 16040 15502 16068 17546
rect 16132 17134 16160 18906
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16224 16794 16252 20470
rect 16316 19922 16344 20742
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16500 20058 16528 20198
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16500 18970 16528 19722
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16592 18834 16620 21286
rect 16670 19816 16726 19825
rect 16670 19751 16726 19760
rect 16684 19378 16712 19751
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16776 18902 16804 21422
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16868 19514 16896 20266
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16960 19446 16988 21966
rect 17236 21962 17264 22918
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17236 21706 17264 21898
rect 17144 21678 17264 21706
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 17052 20942 17080 21354
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 17052 20466 17080 20878
rect 17144 20602 17172 21678
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 17052 19310 17080 20402
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17144 19378 17172 20198
rect 17236 19825 17264 21558
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 17328 19990 17356 20198
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17222 19816 17278 19825
rect 17222 19751 17278 19760
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16764 18896 16816 18902
rect 16764 18838 16816 18844
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16960 18737 16988 19110
rect 16946 18728 17002 18737
rect 16946 18663 17002 18672
rect 16960 18358 16988 18663
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 17038 18320 17094 18329
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 16454 16252 16730
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16040 13734 16068 15438
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 13938 16252 14758
rect 16316 13977 16344 18226
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16408 17270 16436 17682
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16500 17066 16528 17478
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16500 15638 16528 15846
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16302 13968 16358 13977
rect 16212 13932 16264 13938
rect 16302 13903 16358 13912
rect 16212 13874 16264 13880
rect 16500 13818 16528 15574
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16408 13790 16528 13818
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 15856 13518 15976 13546
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15580 13144 15700 13172
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14752 9926 14780 10134
rect 15028 9926 15056 10610
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 14660 8838 14688 9590
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14936 7886 14964 9318
rect 15120 9042 15148 9454
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15120 8430 15148 8978
rect 15212 8634 15240 9590
rect 15304 8906 15332 10950
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15396 8786 15424 11494
rect 15488 9042 15516 11562
rect 15580 11354 15608 13144
rect 15764 12850 15792 13330
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15764 12306 15792 12786
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 11694 15700 12038
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15856 11218 15884 13126
rect 15948 12782 15976 13518
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 16132 12442 16160 13670
rect 16316 13326 16344 13738
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16408 12918 16436 13790
rect 16486 13696 16542 13705
rect 16486 13631 16542 13640
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15672 8974 15700 10474
rect 15764 9178 15792 11154
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15856 9994 15884 10746
rect 16028 10600 16080 10606
rect 15934 10568 15990 10577
rect 16028 10542 16080 10548
rect 15934 10503 15936 10512
rect 15988 10503 15990 10512
rect 15936 10474 15988 10480
rect 16040 10266 16068 10542
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15856 9586 15884 9930
rect 16040 9654 16068 9998
rect 16132 9654 16160 12378
rect 16408 12374 16436 12650
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16224 11558 16252 12310
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16500 10674 16528 13631
rect 16592 12782 16620 17818
rect 16684 17678 16712 18090
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16670 16008 16726 16017
rect 16670 15943 16726 15952
rect 16684 12918 16712 15943
rect 16776 15706 16804 18294
rect 16960 16726 16988 18294
rect 17038 18255 17040 18264
rect 17092 18255 17094 18264
rect 17040 18226 17092 18232
rect 17052 17338 17080 18226
rect 17144 17728 17172 19314
rect 17236 17882 17264 19654
rect 17328 19514 17356 19654
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17420 19394 17448 20334
rect 17512 19417 17540 21286
rect 17328 19366 17448 19394
rect 17498 19408 17554 19417
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17328 17746 17356 19366
rect 17498 19343 17554 19352
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17420 18193 17448 18566
rect 17512 18358 17540 18566
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17406 18184 17462 18193
rect 17406 18119 17462 18128
rect 17316 17740 17368 17746
rect 17144 17700 17264 17728
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17144 16182 17172 16390
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16868 14278 16896 16050
rect 17236 16046 17264 17700
rect 17316 17682 17368 17688
rect 17512 17610 17540 18294
rect 17604 18057 17632 23122
rect 18248 23066 18276 23122
rect 18248 23038 18368 23066
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18340 22438 18368 23038
rect 18512 23044 18564 23050
rect 18512 22986 18564 22992
rect 18524 22710 18552 22986
rect 18512 22704 18564 22710
rect 18512 22646 18564 22652
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18328 22432 18380 22438
rect 18328 22374 18380 22380
rect 17866 21992 17922 22001
rect 17866 21927 17922 21936
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17590 18048 17646 18057
rect 17590 17983 17646 17992
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17512 16590 17540 16662
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17406 16280 17462 16289
rect 17406 16215 17408 16224
rect 17460 16215 17462 16224
rect 17408 16186 17460 16192
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15348 16988 15846
rect 17132 15360 17184 15366
rect 16960 15320 17132 15348
rect 17132 15302 17184 15308
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16856 14272 16908 14278
rect 16854 14240 16856 14249
rect 16908 14240 16910 14249
rect 16854 14175 16910 14184
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16776 13938 16804 14010
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16776 12850 16804 13194
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16670 12744 16726 12753
rect 16670 12679 16726 12688
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16592 10130 16620 12582
rect 16684 11354 16712 12679
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16684 10470 16712 11018
rect 16776 10742 16804 12038
rect 16868 11150 16896 14010
rect 17052 13870 17080 14418
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17144 13569 17172 15302
rect 17236 14890 17264 15982
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17130 13560 17186 13569
rect 17130 13495 17186 13504
rect 17130 13288 17186 13297
rect 16960 13232 17130 13240
rect 16960 13212 17132 13232
rect 16960 12850 16988 13212
rect 17184 13223 17186 13232
rect 17132 13194 17184 13200
rect 17236 13138 17264 14826
rect 17144 13110 17264 13138
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16960 12306 16988 12786
rect 17052 12646 17080 12854
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16960 11830 16988 12242
rect 17052 12238 17080 12582
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 17144 11014 17172 13110
rect 17328 12850 17356 15846
rect 17420 15570 17448 16050
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17420 14414 17448 14894
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17420 13734 17448 14350
rect 17512 14074 17540 14554
rect 17604 14074 17632 15914
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17420 12374 17448 13670
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17512 12306 17540 13806
rect 17696 13297 17724 19722
rect 17774 18456 17830 18465
rect 17774 18391 17830 18400
rect 17788 17678 17816 18391
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17880 15706 17908 21927
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18340 20058 18368 21490
rect 18432 20806 18460 22510
rect 18524 22030 18552 22646
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 16674 18368 19382
rect 18432 19378 18460 19994
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18524 18766 18552 20946
rect 18616 19854 18644 24006
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18800 22982 18828 23462
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 21622 18828 22918
rect 18892 22778 18920 23054
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18984 22098 19012 26200
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 19076 23186 19104 24346
rect 19628 24342 19656 26200
rect 20272 24342 20300 26200
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 19616 24336 19668 24342
rect 19616 24278 19668 24284
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19260 23186 19288 23734
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19260 22710 19288 23122
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19352 22642 19380 22714
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18984 21486 19012 21830
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18892 20602 18920 21422
rect 19352 21350 19380 22578
rect 19444 22030 19472 24006
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19628 23254 19656 23802
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20364 23254 20392 23734
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 20352 23248 20404 23254
rect 20352 23190 20404 23196
rect 19524 23044 19576 23050
rect 19524 22986 19576 22992
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19444 21350 19472 21558
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19352 20942 19380 21286
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19444 20806 19472 21286
rect 19432 20800 19484 20806
rect 19338 20768 19394 20777
rect 19432 20742 19484 20748
rect 19338 20703 19394 20712
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18892 19990 18920 20538
rect 18880 19984 18932 19990
rect 18694 19952 18750 19961
rect 18880 19926 18932 19932
rect 19352 19922 19380 20703
rect 19444 20466 19472 20742
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 18694 19887 18750 19896
rect 19340 19916 19392 19922
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18248 16658 18368 16674
rect 18236 16652 18368 16658
rect 18288 16646 18368 16652
rect 18236 16594 18288 16600
rect 18340 16454 18368 16646
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17880 15366 17908 15642
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18052 14884 18104 14890
rect 18052 14826 18104 14832
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17682 13288 17738 13297
rect 17682 13223 17738 13232
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17224 12096 17276 12102
rect 17222 12064 17224 12073
rect 17276 12064 17278 12073
rect 17222 11999 17278 12008
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 10266 16712 10406
rect 17236 10266 17264 10950
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17328 10198 17356 10950
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16486 9616 16542 9625
rect 15844 9580 15896 9586
rect 16486 9551 16488 9560
rect 15844 9522 15896 9528
rect 16540 9551 16542 9560
rect 16488 9522 16540 9528
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15304 8758 15424 8786
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15212 8498 15240 8570
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13372 3058 13400 3878
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14844 3126 14872 3334
rect 15212 3194 15240 8434
rect 15304 3602 15332 8758
rect 15856 6254 15884 9046
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 16040 5574 16068 9318
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16500 8498 16528 8978
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16592 8566 16620 8842
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16408 7954 16436 8366
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15764 4049 15792 4082
rect 15750 4040 15806 4049
rect 15750 3975 15806 3984
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 13832 800 13860 2450
rect 14476 2446 14504 2926
rect 15304 2514 15332 3538
rect 15856 3534 15884 4490
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 16592 3126 16620 8502
rect 16684 8362 16712 9658
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16776 7954 16804 8502
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16868 6798 16896 9046
rect 16960 7954 16988 9862
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17144 8566 17172 9114
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17236 8430 17264 9862
rect 17420 9178 17448 11154
rect 17498 10840 17554 10849
rect 17498 10775 17500 10784
rect 17552 10775 17554 10784
rect 17500 10746 17552 10752
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17604 10470 17632 10678
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17512 10198 17540 10406
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17512 8634 17540 9522
rect 17604 9518 17632 10406
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 17696 3670 17724 11154
rect 17788 10724 17816 14758
rect 18064 14414 18092 14826
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 13870 17908 14214
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 14074 18368 16186
rect 18432 15910 18460 17614
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18524 15609 18552 18226
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 17610 18644 18022
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17202 18644 17546
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18616 16425 18644 16594
rect 18602 16416 18658 16425
rect 18602 16351 18658 16360
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18510 15600 18566 15609
rect 18510 15535 18566 15544
rect 18616 15502 18644 16186
rect 18708 15706 18736 19887
rect 19340 19858 19392 19864
rect 19338 19680 19394 19689
rect 19338 19615 19394 19624
rect 19352 18698 19380 19615
rect 19444 19310 19472 20402
rect 19536 19718 19564 22986
rect 19812 22234 19840 22986
rect 19800 22228 19852 22234
rect 19800 22170 19852 22176
rect 19708 22160 19760 22166
rect 19708 22102 19760 22108
rect 19720 21010 19748 22102
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19628 20262 19656 20742
rect 19720 20602 19748 20946
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19524 19440 19576 19446
rect 19524 19382 19576 19388
rect 19432 19304 19484 19310
rect 19430 19272 19432 19281
rect 19484 19272 19486 19281
rect 19430 19207 19486 19216
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18800 16425 18828 17478
rect 19168 17338 19196 18294
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18892 16658 18920 17206
rect 18984 16794 19012 17206
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19076 16794 19104 17138
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 18786 16416 18842 16425
rect 18786 16351 18842 16360
rect 18800 15994 18828 16351
rect 18892 16114 18920 16594
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18800 15966 18920 15994
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18800 15706 18828 15846
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18432 14618 18460 15438
rect 18604 15088 18656 15094
rect 18708 15076 18736 15642
rect 18800 15609 18828 15642
rect 18786 15600 18842 15609
rect 18786 15535 18842 15544
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18656 15048 18736 15076
rect 18604 15030 18656 15036
rect 18800 15008 18828 15098
rect 18708 14980 18828 15008
rect 18708 14940 18736 14980
rect 18616 14912 18736 14940
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18420 14408 18472 14414
rect 18616 14396 18644 14912
rect 18786 14648 18842 14657
rect 18786 14583 18842 14592
rect 18800 14414 18828 14583
rect 18472 14368 18644 14396
rect 18788 14408 18840 14414
rect 18420 14350 18472 14356
rect 18788 14350 18840 14356
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18050 13968 18106 13977
rect 18050 13903 18106 13912
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 12442 17908 13806
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17972 13530 18000 13738
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18064 13326 18092 13903
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17880 11880 17908 12378
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17960 11892 18012 11898
rect 17880 11852 17960 11880
rect 17960 11834 18012 11840
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 17788 10696 18000 10724
rect 17788 9625 17816 10696
rect 17972 10606 18000 10696
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17774 9616 17830 9625
rect 17774 9551 17830 9560
rect 17880 8906 17908 10066
rect 18156 9976 18184 10746
rect 18340 10266 18368 13466
rect 18432 12889 18460 14350
rect 18512 14272 18564 14278
rect 18604 14272 18656 14278
rect 18512 14214 18564 14220
rect 18602 14240 18604 14249
rect 18656 14240 18658 14249
rect 18524 13308 18552 14214
rect 18602 14175 18658 14184
rect 18616 13938 18644 14175
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18892 13870 18920 15966
rect 18984 15502 19012 16390
rect 19076 15978 19104 16730
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 19156 15904 19208 15910
rect 19154 15872 19156 15881
rect 19208 15872 19210 15881
rect 19154 15807 19210 15816
rect 19352 15706 19380 18634
rect 19430 18048 19486 18057
rect 19430 17983 19486 17992
rect 19444 17882 19472 17983
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19536 17814 19564 19382
rect 19628 19174 19656 20198
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19628 18698 19656 19110
rect 19720 18834 19748 20538
rect 19812 19310 19840 20946
rect 20364 20777 20392 23190
rect 20640 21622 20668 24210
rect 20824 24206 20852 24550
rect 20916 24274 20944 26200
rect 21560 24886 21588 26200
rect 21548 24880 21600 24886
rect 21548 24822 21600 24828
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21468 23866 21496 24142
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 20824 23186 20852 23462
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20824 22642 20852 23122
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 21008 21690 21036 23462
rect 21744 23186 21772 23598
rect 22204 23225 22232 26200
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22190 23216 22246 23225
rect 21732 23180 21784 23186
rect 22190 23151 22246 23160
rect 21732 23122 21784 23128
rect 21548 23044 21600 23050
rect 21548 22986 21600 22992
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20350 20768 20406 20777
rect 20350 20703 20406 20712
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19904 20058 19932 20538
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19904 18970 19932 19450
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 19628 18222 19656 18634
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19628 17882 19656 18158
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 19076 15026 19104 15642
rect 19246 15192 19302 15201
rect 19246 15127 19248 15136
rect 19300 15127 19302 15136
rect 19248 15098 19300 15104
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19168 15014 19380 15042
rect 18970 14920 19026 14929
rect 18970 14855 18972 14864
rect 19024 14855 19026 14864
rect 18972 14826 19024 14832
rect 19168 14793 19196 15014
rect 19248 14816 19300 14822
rect 19154 14784 19210 14793
rect 19248 14758 19300 14764
rect 19154 14719 19210 14728
rect 19260 14550 19288 14758
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18984 13394 19012 13806
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18524 13280 18644 13308
rect 18510 13016 18566 13025
rect 18510 12951 18566 12960
rect 18418 12880 18474 12889
rect 18418 12815 18474 12824
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18340 10130 18368 10202
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18156 9948 18368 9976
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17880 7426 17908 8570
rect 18340 7886 18368 9948
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18432 7750 18460 11222
rect 18524 11082 18552 12951
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10062 18552 11018
rect 18616 10130 18644 13280
rect 18984 12918 19012 13330
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18892 12170 18920 12786
rect 19352 12442 19380 15014
rect 19444 14074 19472 16390
rect 19904 15706 19932 17070
rect 19996 16046 20024 20198
rect 20088 20058 20116 20266
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20456 19718 20484 20334
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20628 19780 20680 19786
rect 20628 19722 20680 19728
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20456 18834 20484 19654
rect 20534 19272 20590 19281
rect 20534 19207 20590 19216
rect 20548 19174 20576 19207
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20548 18340 20576 19110
rect 20640 18873 20668 19722
rect 20732 18902 20760 19790
rect 20916 19174 20944 19790
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20720 18896 20772 18902
rect 20626 18864 20682 18873
rect 20720 18838 20772 18844
rect 21192 18834 21220 22714
rect 21560 22642 21588 22986
rect 21744 22642 21772 23122
rect 21824 23044 21876 23050
rect 21824 22986 21876 22992
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21836 22778 21864 22986
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21560 22420 21588 22578
rect 21836 22506 21864 22714
rect 21824 22500 21876 22506
rect 21824 22442 21876 22448
rect 21640 22432 21692 22438
rect 21560 22392 21640 22420
rect 21640 22374 21692 22380
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21364 21412 21416 21418
rect 21364 21354 21416 21360
rect 21376 19718 21404 21354
rect 21468 19922 21496 21830
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21560 20398 21588 21558
rect 21652 21350 21680 22374
rect 21928 22094 21956 22986
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22020 22778 22048 22918
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22008 22636 22060 22642
rect 22060 22596 22140 22624
rect 22008 22578 22060 22584
rect 21836 22066 21956 22094
rect 21836 21978 21864 22066
rect 21744 21962 21864 21978
rect 21732 21956 21864 21962
rect 21784 21950 21864 21956
rect 21732 21898 21784 21904
rect 22112 21434 22140 22596
rect 22572 22137 22600 23598
rect 22664 23066 22692 24074
rect 22744 23588 22796 23594
rect 22744 23530 22796 23536
rect 22756 23254 22784 23530
rect 22744 23248 22796 23254
rect 22744 23190 22796 23196
rect 22664 23038 22784 23066
rect 22558 22128 22614 22137
rect 22558 22063 22614 22072
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22192 21480 22244 21486
rect 22112 21428 22192 21434
rect 22112 21422 22244 21428
rect 22112 21406 22232 21422
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21822 21040 21878 21049
rect 21822 20975 21878 20984
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 20626 18799 20682 18808
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20628 18352 20680 18358
rect 20548 18312 20628 18340
rect 20680 18312 20760 18340
rect 20628 18294 20680 18300
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19536 14006 19564 14214
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19628 13938 19656 14350
rect 19720 14278 19748 15302
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19720 13734 19748 14214
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19444 12306 19472 13466
rect 19812 13190 19840 14282
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13394 20024 13670
rect 20088 13530 20116 14418
rect 20180 14074 20208 14486
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18708 11558 18736 11698
rect 18800 11694 18828 12106
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18800 11234 18828 11630
rect 18892 11354 18920 12106
rect 19076 11694 19104 12174
rect 19064 11688 19116 11694
rect 18984 11648 19064 11676
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18800 11206 18920 11234
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18616 9602 18644 10066
rect 18524 9574 18644 9602
rect 18524 8090 18552 9574
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 8634 18644 9454
rect 18708 8974 18736 10610
rect 18800 9382 18828 11018
rect 18892 9518 18920 11206
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18892 9042 18920 9454
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18616 7954 18644 8570
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17880 7410 18000 7426
rect 17880 7404 18012 7410
rect 17880 7398 17960 7404
rect 17960 7346 18012 7352
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 4214 18368 6190
rect 18892 5234 18920 7958
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18328 4208 18380 4214
rect 18328 4150 18380 4156
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 18984 3466 19012 11648
rect 19064 11630 19116 11636
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19168 11286 19196 11494
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19444 11218 19472 12242
rect 19536 12170 19564 12718
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19076 8634 19104 11086
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19168 10266 19196 10542
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19628 10130 19656 12786
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19720 10810 19748 12718
rect 19812 11762 19840 12786
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19812 10674 19840 10950
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19812 10198 19840 10610
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19444 9042 19472 10066
rect 19800 9988 19852 9994
rect 19800 9930 19852 9936
rect 19708 9648 19760 9654
rect 19812 9636 19840 9930
rect 19760 9608 19840 9636
rect 19708 9590 19760 9596
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19628 9178 19656 9454
rect 19812 9382 19840 9608
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19444 8090 19472 8978
rect 19812 8974 19840 9318
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19812 8566 19840 8910
rect 19904 8634 19932 12242
rect 19996 11898 20024 13126
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20088 11218 20116 12106
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20180 11082 20208 14010
rect 20272 13530 20300 15302
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20364 13462 20392 17614
rect 20732 17610 20760 18312
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20536 17264 20588 17270
rect 20732 17252 20760 17546
rect 20588 17224 20760 17252
rect 20536 17206 20588 17212
rect 20732 16590 20760 17224
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20732 16454 20760 16526
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 16182 20760 16390
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20732 15858 20760 15914
rect 20640 15830 20760 15858
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14346 20576 14758
rect 20640 14482 20668 15830
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20626 14376 20682 14385
rect 20536 14340 20588 14346
rect 20626 14311 20682 14320
rect 20536 14282 20588 14288
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20272 10674 20300 12718
rect 20456 11830 20484 12718
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20548 11830 20576 12174
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 11286 20392 11630
rect 20456 11286 20484 11766
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20272 10266 20300 10610
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20456 9994 20484 11018
rect 20640 10538 20668 14311
rect 20732 11898 20760 15030
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20824 11762 20852 15982
rect 20916 15706 20944 18702
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21192 17882 21220 18022
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20916 13530 20944 14962
rect 21008 14958 21036 16662
rect 21100 14958 21128 17818
rect 21284 17270 21312 18226
rect 21272 17264 21324 17270
rect 21272 17206 21324 17212
rect 21284 16726 21312 17206
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21376 16572 21404 18566
rect 21456 18080 21508 18086
rect 21560 18068 21588 20334
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21508 18040 21588 18068
rect 21456 18022 21508 18028
rect 21192 16544 21404 16572
rect 21192 15178 21220 16544
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15366 21312 15846
rect 21468 15570 21496 18022
rect 21652 17898 21680 18566
rect 21560 17870 21680 17898
rect 21560 17270 21588 17870
rect 21744 17746 21772 19654
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21652 17610 21680 17682
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21652 16182 21680 17002
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21652 15910 21680 16118
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21192 15150 21312 15178
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 20994 14512 21050 14521
rect 21100 14482 21128 14894
rect 20994 14447 21050 14456
rect 21088 14476 21140 14482
rect 21008 13841 21036 14447
rect 21088 14418 21140 14424
rect 20994 13832 21050 13841
rect 20994 13767 21050 13776
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21008 13394 21036 13767
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 20902 13288 20958 13297
rect 21008 13258 21036 13330
rect 20902 13223 20958 13232
rect 20996 13252 21048 13258
rect 20916 12986 20944 13223
rect 20996 13194 21048 13200
rect 21284 13190 21312 15150
rect 21376 14482 21404 15506
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21376 14074 21404 14418
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21008 12714 21036 12786
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 20994 12608 21050 12617
rect 20994 12543 21050 12552
rect 21008 12306 21036 12543
rect 21284 12374 21312 13126
rect 21468 12714 21496 15302
rect 21560 14958 21588 15438
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21560 13394 21588 14554
rect 21652 14346 21680 15846
rect 21744 14906 21772 17206
rect 21836 15094 21864 20975
rect 22112 20466 22140 21406
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22204 20874 22232 21286
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22296 20754 22324 21966
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22374 21720 22430 21729
rect 22374 21655 22430 21664
rect 22388 21457 22416 21655
rect 22374 21448 22430 21457
rect 22374 21383 22430 21392
rect 22480 21350 22508 21830
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22466 21040 22522 21049
rect 22572 21010 22600 21830
rect 22664 21010 22692 22034
rect 22466 20975 22522 20984
rect 22560 21004 22612 21010
rect 22480 20777 22508 20975
rect 22560 20946 22612 20952
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22466 20768 22522 20777
rect 22296 20726 22416 20754
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22190 20496 22246 20505
rect 22100 20460 22152 20466
rect 22190 20431 22246 20440
rect 22100 20402 22152 20408
rect 22112 19446 22140 20402
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22112 17746 22140 19382
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 22112 17270 22140 17682
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21744 14878 21864 14906
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21744 14482 21772 14758
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21836 14385 21864 14878
rect 21822 14376 21878 14385
rect 21640 14340 21692 14346
rect 21822 14311 21878 14320
rect 21640 14282 21692 14288
rect 21652 13938 21680 14282
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21928 13870 21956 15982
rect 22204 15978 22232 20431
rect 22296 19922 22324 20538
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22296 19242 22324 19722
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22296 18970 22324 19178
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22296 17678 22324 18702
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22296 17066 22324 17614
rect 22388 17241 22416 20726
rect 22466 20703 22522 20712
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22374 17232 22430 17241
rect 22374 17167 22430 17176
rect 22374 17096 22430 17105
rect 22284 17060 22336 17066
rect 22374 17031 22430 17040
rect 22284 17002 22336 17008
rect 22388 16998 22416 17031
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22480 16658 22508 18022
rect 22572 17542 22600 20334
rect 22756 20330 22784 23038
rect 22848 22681 22876 26200
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23492 23798 23520 26200
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23294 23080 23350 23089
rect 23294 23015 23350 23024
rect 23308 22982 23336 23015
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 22834 22672 22890 22681
rect 22834 22607 22890 22616
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22940 21894 22968 21966
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22848 21486 22876 21626
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 21078 23336 22510
rect 23388 22500 23440 22506
rect 23388 22442 23440 22448
rect 23400 22098 23428 22442
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 22166 23520 22374
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23584 21962 23612 23666
rect 23756 23656 23808 23662
rect 23756 23598 23808 23604
rect 23664 23588 23716 23594
rect 23664 23530 23716 23536
rect 23676 23322 23704 23530
rect 23768 23322 23796 23598
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22574 23704 22918
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23386 21448 23442 21457
rect 23386 21383 23442 21392
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22940 20602 22968 20878
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22742 20224 22798 20233
rect 22742 20159 22798 20168
rect 22756 19718 22784 20159
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23400 19961 23428 21383
rect 23492 21078 23520 21898
rect 23664 21888 23716 21894
rect 23768 21865 23796 22578
rect 23664 21830 23716 21836
rect 23754 21856 23810 21865
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23676 20913 23704 21830
rect 23754 21791 23810 21800
rect 23860 21706 23888 23462
rect 23952 22710 23980 24006
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23952 22545 23980 22646
rect 23938 22536 23994 22545
rect 23938 22471 23994 22480
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23768 21678 23888 21706
rect 23662 20904 23718 20913
rect 23572 20868 23624 20874
rect 23662 20839 23718 20848
rect 23572 20810 23624 20816
rect 23386 19952 23442 19961
rect 23386 19887 23442 19896
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 22664 19446 22692 19654
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22664 18358 22692 19382
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22756 18290 22784 18906
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23308 17882 23336 19314
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22112 14074 22140 15506
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 21916 13864 21968 13870
rect 22112 13818 22140 14010
rect 22204 14006 22232 14758
rect 22480 14618 22508 16594
rect 22572 15706 22600 17274
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 22756 16658 22784 17206
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23400 16794 23428 18226
rect 23492 17678 23520 18634
rect 23584 17882 23612 20810
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23676 18154 23704 20470
rect 23768 20466 23796 21678
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23952 19922 23980 21966
rect 24044 20534 24072 22374
rect 24122 21856 24178 21865
rect 24122 21791 24178 21800
rect 24136 21622 24164 21791
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24136 20874 24164 21558
rect 24320 21146 24348 26302
rect 24766 26200 24822 27000
rect 25410 26200 25466 27000
rect 26054 26200 26110 27000
rect 26698 26330 26754 27000
rect 26698 26302 27016 26330
rect 26698 26200 26754 26302
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 24504 24342 24532 24754
rect 24780 24682 24808 26200
rect 24768 24676 24820 24682
rect 24768 24618 24820 24624
rect 24492 24336 24544 24342
rect 24492 24278 24544 24284
rect 25424 24206 25452 26200
rect 25964 24880 26016 24886
rect 25964 24822 26016 24828
rect 25780 24336 25832 24342
rect 25778 24304 25780 24313
rect 25832 24304 25834 24313
rect 25778 24239 25834 24248
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24872 23662 24900 24006
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 23186 24900 23462
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24596 21729 24624 22374
rect 24688 22273 24716 22986
rect 24780 22681 24808 22986
rect 24766 22672 24822 22681
rect 24964 22642 24992 23666
rect 25332 22982 25360 24074
rect 25424 23254 25452 24142
rect 25872 23792 25924 23798
rect 25872 23734 25924 23740
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25412 23248 25464 23254
rect 25412 23190 25464 23196
rect 25320 22976 25372 22982
rect 25318 22944 25320 22953
rect 25372 22944 25374 22953
rect 25318 22879 25374 22888
rect 24766 22607 24822 22616
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24860 22500 24912 22506
rect 24674 22264 24730 22273
rect 24674 22199 24730 22208
rect 24780 21894 24808 22471
rect 24860 22442 24912 22448
rect 24872 22166 24900 22442
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 24860 22160 24912 22166
rect 24860 22102 24912 22108
rect 25148 22098 25176 22374
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 25608 22030 25636 23598
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24582 21720 24638 21729
rect 24582 21655 24638 21664
rect 24596 21486 24624 21655
rect 24584 21480 24636 21486
rect 24584 21422 24636 21428
rect 24308 21140 24360 21146
rect 24308 21082 24360 21088
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24320 20942 24348 21082
rect 24780 20942 24808 21082
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24124 20868 24176 20874
rect 24676 20868 24728 20874
rect 24124 20810 24176 20816
rect 24596 20828 24676 20856
rect 24596 20534 24624 20828
rect 24676 20810 24728 20816
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 24584 20528 24636 20534
rect 24584 20470 24636 20476
rect 23940 19916 23992 19922
rect 23940 19858 23992 19864
rect 24228 19718 24256 20470
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 23768 19553 23796 19654
rect 23754 19544 23810 19553
rect 23754 19479 23810 19488
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23860 18698 23888 19110
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 24136 18358 24164 18702
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 23664 18148 23716 18154
rect 23664 18090 23716 18096
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23492 17338 23520 17614
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 22742 15736 22798 15745
rect 22560 15700 22612 15706
rect 22742 15671 22798 15680
rect 22560 15642 22612 15648
rect 22756 14890 22784 15671
rect 22848 15162 22876 16390
rect 23308 16250 23336 16390
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22560 14544 22612 14550
rect 22560 14486 22612 14492
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 21916 13806 21968 13812
rect 22020 13802 22140 13818
rect 22008 13796 22140 13802
rect 22060 13790 22140 13796
rect 22008 13738 22060 13744
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 21180 12232 21232 12238
rect 21232 12180 21496 12186
rect 21180 12174 21496 12180
rect 21192 12170 21496 12174
rect 21192 12164 21508 12170
rect 21192 12158 21456 12164
rect 21456 12106 21508 12112
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20916 11370 20944 12038
rect 21192 11694 21220 12038
rect 21560 11694 21588 13330
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21652 11558 21680 13194
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21744 12238 21772 12378
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 20732 11342 20944 11370
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19812 7886 19840 8502
rect 19904 7954 19932 8570
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19628 6798 19656 7754
rect 19812 7410 19840 7822
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 20732 7274 20760 11342
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 21100 10130 21128 10542
rect 21284 10470 21312 11494
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21100 9722 21128 10066
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21468 8974 21496 9862
rect 21548 9648 21600 9654
rect 21546 9616 21548 9625
rect 21600 9616 21602 9625
rect 21546 9551 21602 9560
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21468 8430 21496 8910
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4758 19104 5102
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 19076 3126 19104 4694
rect 19260 4690 19288 6598
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19352 3194 19380 3402
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15948 800 15976 2314
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 2926
rect 19444 2446 19472 6054
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 3738 20024 4558
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19996 2514 20024 3674
rect 20640 3058 20668 4966
rect 21008 3534 21036 7754
rect 21192 7478 21220 8366
rect 21468 7886 21496 8366
rect 21928 8090 21956 12786
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 22020 11898 22048 12718
rect 22374 12336 22430 12345
rect 22374 12271 22376 12280
rect 22428 12271 22430 12280
rect 22376 12242 22428 12248
rect 22388 11898 22416 12242
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 10690 22048 11494
rect 22204 11150 22232 11766
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22480 11558 22508 11698
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 11354 22508 11494
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22284 10736 22336 10742
rect 22020 10662 22232 10690
rect 22284 10678 22336 10684
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10062 22048 10542
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22020 8906 22048 9318
rect 22112 9178 22140 10406
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 22020 8498 22048 8842
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22112 8430 22140 9114
rect 22204 8922 22232 10662
rect 22296 9382 22324 10678
rect 22480 9994 22508 11290
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22480 9178 22508 9930
rect 22572 9654 22600 14486
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 13530 22784 13670
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22848 13025 22876 14350
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23216 14074 23244 14214
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22834 13016 22890 13025
rect 22834 12951 22890 12960
rect 22744 12776 22796 12782
rect 22848 12764 22876 12951
rect 22796 12736 22876 12764
rect 22928 12776 22980 12782
rect 22926 12744 22928 12753
rect 22980 12744 22982 12753
rect 22744 12718 22796 12724
rect 22756 12617 22784 12718
rect 22926 12679 22982 12688
rect 22940 12646 22968 12679
rect 22928 12640 22980 12646
rect 22742 12608 22798 12617
rect 22928 12582 22980 12588
rect 22742 12543 22798 12552
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11354 23336 14962
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23400 12102 23428 13194
rect 23492 12986 23520 15914
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23584 12866 23612 16050
rect 23676 13530 23704 16390
rect 23768 15162 23796 17682
rect 24136 17270 24164 18294
rect 24124 17264 24176 17270
rect 24124 17206 24176 17212
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 24136 15026 24164 15302
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23860 13326 23888 14214
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23676 12986 23704 13126
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23860 12918 23888 13126
rect 23848 12912 23900 12918
rect 23584 12838 23796 12866
rect 23848 12854 23900 12860
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23584 12617 23612 12718
rect 23570 12608 23626 12617
rect 23570 12543 23626 12552
rect 23676 12306 23704 12718
rect 23768 12374 23796 12838
rect 23756 12368 23808 12374
rect 23756 12310 23808 12316
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23492 11694 23520 12242
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22664 10810 22692 11086
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 23584 10538 23612 11018
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22204 8894 22324 8922
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22204 7886 22232 8774
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21284 7546 21312 7754
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21468 7342 21496 7686
rect 22296 7546 22324 8894
rect 23400 8838 23428 9522
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 22468 8356 22520 8362
rect 22520 8316 22600 8344
rect 22468 8298 22520 8304
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22572 7342 22600 8316
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21928 4690 21956 6598
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23400 4826 23428 8774
rect 23584 7954 23612 10474
rect 23768 10266 23796 11154
rect 23952 11082 23980 13806
rect 24044 13546 24072 14894
rect 24136 14822 24164 14962
rect 24228 14958 24256 19654
rect 24492 19440 24544 19446
rect 24596 19428 24624 20470
rect 24544 19400 24624 19428
rect 24492 19382 24544 19388
rect 24596 19009 24624 19400
rect 24582 19000 24638 19009
rect 24582 18935 24638 18944
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24504 17134 24532 18294
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24504 16046 24532 17070
rect 24596 16590 24624 18935
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24688 17649 24716 18226
rect 24674 17640 24730 17649
rect 24674 17575 24730 17584
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24596 16182 24624 16526
rect 24584 16176 24636 16182
rect 24584 16118 24636 16124
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24688 15978 24716 17478
rect 24780 17218 24808 18566
rect 24872 17338 24900 21966
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25148 21350 25176 21490
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 24964 20058 24992 21082
rect 25148 20777 25176 21286
rect 25240 21185 25268 21422
rect 25226 21176 25282 21185
rect 25226 21111 25282 21120
rect 25134 20768 25190 20777
rect 25134 20703 25190 20712
rect 25226 20496 25282 20505
rect 25226 20431 25282 20440
rect 25240 20058 25268 20431
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24964 17746 24992 19246
rect 25056 18630 25084 19994
rect 25332 19938 25360 21830
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25424 21486 25452 21626
rect 25412 21480 25464 21486
rect 25412 21422 25464 21428
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25594 20768 25650 20777
rect 25148 19910 25360 19938
rect 25148 18630 25176 19910
rect 25320 19780 25372 19786
rect 25320 19722 25372 19728
rect 25228 19236 25280 19242
rect 25228 19178 25280 19184
rect 25240 18834 25268 19178
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25134 18320 25190 18329
rect 25134 18255 25136 18264
rect 25188 18255 25190 18264
rect 25136 18226 25188 18232
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17746 25084 18022
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25148 17610 25176 18226
rect 25332 18222 25360 19722
rect 25424 19514 25452 20742
rect 25594 20703 25650 20712
rect 25608 20398 25636 20703
rect 25700 20602 25728 23054
rect 25884 22710 25912 23734
rect 25872 22704 25924 22710
rect 25872 22646 25924 22652
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25792 20874 25820 21830
rect 25872 21344 25924 21350
rect 25870 21312 25872 21321
rect 25924 21312 25926 21321
rect 25870 21247 25926 21256
rect 25976 20913 26004 24822
rect 26068 24206 26096 26200
rect 26332 24812 26384 24818
rect 26332 24754 26384 24760
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 26344 24342 26372 24754
rect 26436 24410 26464 24754
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26332 24336 26384 24342
rect 26332 24278 26384 24284
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26436 24138 26464 24346
rect 26606 24304 26662 24313
rect 26606 24239 26608 24248
rect 26660 24239 26662 24248
rect 26608 24210 26660 24216
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 26988 24070 27016 26302
rect 27342 26200 27398 27000
rect 27986 26330 28042 27000
rect 27986 26302 28488 26330
rect 27986 26200 28042 26302
rect 27356 24274 27384 26200
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27252 24132 27304 24138
rect 27252 24074 27304 24080
rect 27344 24132 27396 24138
rect 27344 24074 27396 24080
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 26344 22438 26372 23122
rect 26620 22574 26648 23598
rect 27264 23050 27292 24074
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 27264 22778 27292 22986
rect 27356 22778 27384 24074
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 27712 23792 27764 23798
rect 27712 23734 27764 23740
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 27436 22976 27488 22982
rect 27436 22918 27488 22924
rect 27448 22778 27476 22918
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27264 22642 27292 22714
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 26608 22568 26660 22574
rect 26608 22510 26660 22516
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 27068 22228 27120 22234
rect 27068 22170 27120 22176
rect 26608 22160 26660 22166
rect 26422 22128 26478 22137
rect 26608 22102 26660 22108
rect 26422 22063 26478 22072
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 26068 21486 26096 21898
rect 26056 21480 26108 21486
rect 26054 21448 26056 21457
rect 26108 21448 26110 21457
rect 26054 21383 26110 21392
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 26068 21078 26096 21286
rect 26146 21176 26202 21185
rect 26146 21111 26202 21120
rect 26056 21072 26108 21078
rect 26056 21014 26108 21020
rect 25962 20904 26018 20913
rect 25780 20868 25832 20874
rect 25962 20839 26018 20848
rect 25780 20810 25832 20816
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25516 20058 25544 20198
rect 25504 20052 25556 20058
rect 25504 19994 25556 20000
rect 25504 19848 25556 19854
rect 25504 19790 25556 19796
rect 25516 19514 25544 19790
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25608 19310 25636 20334
rect 25700 19378 25728 20538
rect 25872 20528 25924 20534
rect 25872 20470 25924 20476
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25700 18834 25728 19314
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25792 18426 25820 19110
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25228 17604 25280 17610
rect 25228 17546 25280 17552
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 25056 17218 25084 17478
rect 24780 17190 25084 17218
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24780 15858 24808 17190
rect 24688 15830 24808 15858
rect 24308 15564 24360 15570
rect 24308 15506 24360 15512
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24320 13802 24348 15506
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24044 13518 24164 13546
rect 24136 12714 24164 13518
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 24124 12708 24176 12714
rect 24124 12650 24176 12656
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24136 11830 24164 12174
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 24228 10810 24256 13194
rect 24216 10804 24268 10810
rect 24216 10746 24268 10752
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23768 10169 23796 10202
rect 23754 10160 23810 10169
rect 23754 10095 23810 10104
rect 23860 9994 23888 10678
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23860 9586 23888 9930
rect 23952 9926 23980 10542
rect 24320 10266 24348 13398
rect 24412 12986 24440 14214
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24504 13308 24532 13874
rect 24596 13433 24624 14962
rect 24582 13424 24638 13433
rect 24582 13359 24638 13368
rect 24504 13280 24624 13308
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24504 12617 24532 13126
rect 24596 12986 24624 13280
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24490 12608 24546 12617
rect 24490 12543 24546 12552
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24504 11898 24532 12242
rect 24596 12238 24624 12922
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24504 11218 24532 11834
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24596 11150 24624 12174
rect 24688 11558 24716 15830
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 24860 15632 24912 15638
rect 24860 15574 24912 15580
rect 24872 14929 24900 15574
rect 25044 15428 25096 15434
rect 25044 15370 25096 15376
rect 24858 14920 24914 14929
rect 24858 14855 24914 14864
rect 25056 14550 25084 15370
rect 25148 15366 25176 15642
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25148 15162 25176 15302
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25044 14544 25096 14550
rect 25044 14486 25096 14492
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25148 13326 25176 14214
rect 25240 13462 25268 17546
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25332 14074 25360 15506
rect 25516 14618 25544 17070
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25516 14074 25544 14554
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25228 13456 25280 13462
rect 25228 13398 25280 13404
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25332 12918 25360 14010
rect 25608 13530 25636 17138
rect 25884 16658 25912 20470
rect 25976 20466 26004 20839
rect 26160 20618 26188 21111
rect 26436 21010 26464 22063
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 26424 21004 26476 21010
rect 26424 20946 26476 20952
rect 26252 20777 26280 20946
rect 26516 20936 26568 20942
rect 26514 20904 26516 20913
rect 26568 20904 26570 20913
rect 26514 20839 26570 20848
rect 26238 20768 26294 20777
rect 26238 20703 26294 20712
rect 26160 20590 26556 20618
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 26056 20324 26108 20330
rect 26056 20266 26108 20272
rect 26148 20324 26200 20330
rect 26148 20266 26200 20272
rect 26068 20058 26096 20266
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 25976 19938 26004 19994
rect 26054 19952 26110 19961
rect 25976 19910 26054 19938
rect 26054 19887 26056 19896
rect 26108 19887 26110 19896
rect 26056 19858 26108 19864
rect 26160 19446 26188 20266
rect 26424 20256 26476 20262
rect 26424 20198 26476 20204
rect 26148 19440 26200 19446
rect 26146 19408 26148 19417
rect 26200 19408 26202 19417
rect 26436 19378 26464 20198
rect 26146 19343 26202 19352
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26146 19000 26202 19009
rect 26146 18935 26202 18944
rect 26160 18698 26188 18935
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 25962 18320 26018 18329
rect 25962 18255 26018 18264
rect 25976 17270 26004 18255
rect 26056 18148 26108 18154
rect 26056 18090 26108 18096
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 26068 16726 26096 18090
rect 26344 18086 26372 19246
rect 26332 18080 26384 18086
rect 26332 18022 26384 18028
rect 26330 17912 26386 17921
rect 26330 17847 26386 17856
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26056 16720 26108 16726
rect 26056 16662 26108 16668
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 26160 15706 26188 17682
rect 26240 17672 26292 17678
rect 26238 17640 26240 17649
rect 26292 17640 26294 17649
rect 26238 17575 26294 17584
rect 26252 16969 26280 17575
rect 26238 16960 26294 16969
rect 26238 16895 26294 16904
rect 26344 16794 26372 17847
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26240 15700 26292 15706
rect 26240 15642 26292 15648
rect 25686 15464 25742 15473
rect 26252 15434 26280 15642
rect 25686 15399 25688 15408
rect 25740 15399 25742 15408
rect 26240 15428 26292 15434
rect 25688 15370 25740 15376
rect 26240 15370 26292 15376
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 25700 15162 25728 15370
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25884 15094 25912 15302
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25688 14340 25740 14346
rect 25688 14282 25740 14288
rect 25700 14006 25728 14282
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 24872 12646 24900 12854
rect 24952 12776 25004 12782
rect 25228 12776 25280 12782
rect 24952 12718 25004 12724
rect 25226 12744 25228 12753
rect 25280 12744 25282 12753
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24964 12306 24992 12718
rect 25226 12679 25282 12688
rect 25332 12434 25360 12854
rect 25700 12646 25728 13942
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25240 12406 25360 12434
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24584 11144 24636 11150
rect 24636 11104 24716 11132
rect 24584 11086 24636 11092
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23768 9382 23796 9454
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 9042 23796 9318
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23952 6322 23980 9862
rect 24044 9042 24072 9998
rect 24320 9518 24348 10202
rect 24688 9654 24716 11104
rect 24780 10538 24808 11494
rect 25240 11354 25268 12406
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25608 11014 25636 11766
rect 25700 11762 25728 12582
rect 25792 11762 25820 14418
rect 25884 13258 25912 14758
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 26068 13394 26096 14418
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 26056 13184 26108 13190
rect 26056 13126 26108 13132
rect 25976 12986 26004 13126
rect 25964 12980 26016 12986
rect 25964 12922 26016 12928
rect 25964 12640 26016 12646
rect 25964 12582 26016 12588
rect 25976 12374 26004 12582
rect 26068 12442 26096 13126
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 25964 12368 26016 12374
rect 25964 12310 26016 12316
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 26160 11626 26188 14826
rect 26252 12918 26280 15370
rect 26344 15065 26372 15370
rect 26330 15056 26386 15065
rect 26330 14991 26386 15000
rect 26436 14618 26464 19314
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26528 14074 26556 20590
rect 26620 19242 26648 22102
rect 26884 21956 26936 21962
rect 26884 21898 26936 21904
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 26608 19236 26660 19242
rect 26608 19178 26660 19184
rect 26712 18834 26740 21830
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26804 19718 26832 20810
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26792 19236 26844 19242
rect 26792 19178 26844 19184
rect 26700 18828 26752 18834
rect 26700 18770 26752 18776
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26606 17776 26662 17785
rect 26606 17711 26662 17720
rect 26620 17542 26648 17711
rect 26608 17536 26660 17542
rect 26608 17478 26660 17484
rect 26620 16114 26648 17478
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26712 15638 26740 18158
rect 26804 16046 26832 19178
rect 26896 17270 26924 21898
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26988 18986 27016 21490
rect 27080 21185 27108 22170
rect 27172 22166 27200 22578
rect 27528 22500 27580 22506
rect 27528 22442 27580 22448
rect 27160 22160 27212 22166
rect 27160 22102 27212 22108
rect 27540 21706 27568 22442
rect 27632 22234 27660 22986
rect 27724 22506 27752 23734
rect 27816 23730 27844 24006
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27712 22500 27764 22506
rect 27712 22442 27764 22448
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 27816 21962 27844 23462
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28080 22500 28132 22506
rect 28080 22442 28132 22448
rect 28092 22098 28120 22442
rect 28080 22092 28132 22098
rect 28276 22094 28304 22578
rect 28368 22522 28396 24006
rect 28460 23662 28488 26302
rect 28630 26200 28686 27000
rect 29274 26330 29330 27000
rect 29274 26302 29592 26330
rect 29274 26200 29330 26302
rect 28644 24342 28672 26200
rect 29564 24750 29592 26302
rect 29918 26200 29974 27000
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26330 33838 27000
rect 34060 26376 34112 26382
rect 33782 26324 34060 26330
rect 34426 26330 34482 27000
rect 33782 26318 34112 26324
rect 33782 26302 34100 26318
rect 34256 26302 34482 26330
rect 33782 26200 33838 26302
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29748 24410 29776 24550
rect 29736 24404 29788 24410
rect 29736 24346 29788 24352
rect 28632 24336 28684 24342
rect 28632 24278 28684 24284
rect 28632 24064 28684 24070
rect 28632 24006 28684 24012
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28448 23656 28500 23662
rect 28448 23598 28500 23604
rect 28552 23322 28580 23666
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28368 22494 28488 22522
rect 28276 22066 28396 22094
rect 28080 22034 28132 22040
rect 27804 21956 27856 21962
rect 27804 21898 27856 21904
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27540 21690 27660 21706
rect 27540 21684 27672 21690
rect 27540 21678 27620 21684
rect 27620 21626 27672 21632
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27066 21176 27122 21185
rect 27066 21111 27122 21120
rect 27264 21078 27292 21286
rect 27252 21072 27304 21078
rect 27252 21014 27304 21020
rect 27160 21004 27212 21010
rect 27160 20946 27212 20952
rect 27172 19854 27200 20946
rect 27356 20913 27384 21422
rect 27908 21010 27936 21490
rect 27896 21004 27948 21010
rect 27896 20946 27948 20952
rect 27342 20904 27398 20913
rect 27342 20839 27344 20848
rect 27396 20839 27398 20848
rect 27344 20810 27396 20816
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28264 20528 28316 20534
rect 28368 20482 28396 22066
rect 28316 20476 28396 20482
rect 28264 20470 28396 20476
rect 28276 20454 28396 20470
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27356 19922 27384 20198
rect 27804 19984 27856 19990
rect 27804 19926 27856 19932
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 27160 19848 27212 19854
rect 27212 19808 27292 19836
rect 27160 19790 27212 19796
rect 27160 19712 27212 19718
rect 27158 19680 27160 19689
rect 27212 19680 27214 19689
rect 27158 19615 27214 19624
rect 27264 19334 27292 19808
rect 27264 19306 27384 19334
rect 27540 19310 27568 19858
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 26988 18958 27108 18986
rect 27080 18902 27108 18958
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 27264 18426 27292 19110
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 26884 17264 26936 17270
rect 26884 17206 26936 17212
rect 26976 17128 27028 17134
rect 26974 17096 26976 17105
rect 27028 17096 27030 17105
rect 26974 17031 27030 17040
rect 27080 16658 27108 17478
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27066 16144 27122 16153
rect 27066 16079 27122 16088
rect 26792 16040 26844 16046
rect 26792 15982 26844 15988
rect 26700 15632 26752 15638
rect 26700 15574 26752 15580
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26344 11694 26372 12378
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26148 11620 26200 11626
rect 26148 11562 26200 11568
rect 26620 11354 26648 15506
rect 26804 15366 26832 15982
rect 26976 15972 27028 15978
rect 26976 15914 27028 15920
rect 26884 15904 26936 15910
rect 26884 15846 26936 15852
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26700 13252 26752 13258
rect 26700 13194 26752 13200
rect 26712 12374 26740 13194
rect 26804 13025 26832 15302
rect 26790 13016 26846 13025
rect 26790 12951 26846 12960
rect 26700 12368 26752 12374
rect 26700 12310 26752 12316
rect 26896 12170 26924 15846
rect 26988 12442 27016 15914
rect 27080 15706 27108 16079
rect 27068 15700 27120 15706
rect 27068 15642 27120 15648
rect 27066 15600 27122 15609
rect 27066 15535 27122 15544
rect 27080 15348 27108 15535
rect 27172 15502 27200 18022
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27160 15360 27212 15366
rect 27080 15320 27160 15348
rect 27080 15094 27108 15320
rect 27160 15302 27212 15308
rect 27068 15088 27120 15094
rect 27068 15030 27120 15036
rect 27158 13016 27214 13025
rect 27068 12980 27120 12986
rect 27158 12951 27214 12960
rect 27068 12922 27120 12928
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 27080 12170 27108 12922
rect 27172 12918 27200 12951
rect 27160 12912 27212 12918
rect 27160 12854 27212 12860
rect 27264 12434 27292 17002
rect 27356 15910 27384 19306
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27434 19000 27490 19009
rect 27632 18970 27660 19654
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27724 19174 27752 19246
rect 27712 19168 27764 19174
rect 27712 19110 27764 19116
rect 27434 18935 27490 18944
rect 27620 18964 27672 18970
rect 27448 18766 27476 18935
rect 27620 18906 27672 18912
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27448 17678 27476 18702
rect 27724 18426 27752 18906
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27448 16658 27476 17614
rect 27816 17338 27844 19926
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 28172 19304 28224 19310
rect 28172 19246 28224 19252
rect 28184 18766 28212 19246
rect 28276 19242 28304 19450
rect 28354 19408 28410 19417
rect 28354 19343 28356 19352
rect 28408 19343 28410 19352
rect 28356 19314 28408 19320
rect 28264 19236 28316 19242
rect 28264 19178 28316 19184
rect 28172 18760 28224 18766
rect 28172 18702 28224 18708
rect 28368 18630 28396 19314
rect 28460 19174 28488 22494
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 28552 20398 28580 21898
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28540 20052 28592 20058
rect 28540 19994 28592 20000
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 28354 18184 28410 18193
rect 28354 18119 28410 18128
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28276 17542 28304 18022
rect 28264 17536 28316 17542
rect 28264 17478 28316 17484
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27804 17332 27856 17338
rect 27804 17274 27856 17280
rect 27618 17232 27674 17241
rect 28170 17232 28226 17241
rect 27618 17167 27620 17176
rect 27672 17167 27674 17176
rect 27988 17196 28040 17202
rect 27620 17138 27672 17144
rect 28170 17167 28226 17176
rect 27988 17138 28040 17144
rect 27896 17128 27948 17134
rect 27724 17088 27896 17116
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27448 16046 27476 16594
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27540 16114 27568 16390
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27342 15056 27398 15065
rect 27342 14991 27344 15000
rect 27396 14991 27398 15000
rect 27344 14962 27396 14968
rect 27344 14408 27396 14414
rect 27344 14350 27396 14356
rect 27356 13870 27384 14350
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27172 12406 27292 12434
rect 27172 12306 27200 12406
rect 27356 12306 27384 13806
rect 27448 13734 27476 15302
rect 27632 14074 27660 16730
rect 27724 14464 27752 17088
rect 28000 17105 28028 17138
rect 27896 17070 27948 17076
rect 27986 17096 28042 17105
rect 27986 17031 28042 17040
rect 28000 16726 28028 17031
rect 27988 16720 28040 16726
rect 27988 16662 28040 16668
rect 28184 16454 28212 17167
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 16232 28396 18119
rect 28460 17610 28488 18770
rect 28448 17604 28500 17610
rect 28448 17546 28500 17552
rect 28552 17082 28580 19994
rect 28644 19990 28672 24006
rect 29184 23656 29236 23662
rect 29184 23598 29236 23604
rect 29196 23322 29224 23598
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29828 23588 29880 23594
rect 29828 23530 29880 23536
rect 29276 23520 29328 23526
rect 29276 23462 29328 23468
rect 29184 23316 29236 23322
rect 29184 23258 29236 23264
rect 29196 22658 29224 23258
rect 28920 22630 29224 22658
rect 28920 22574 28948 22630
rect 28908 22568 28960 22574
rect 28908 22510 28960 22516
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 28724 21956 28776 21962
rect 28724 21898 28776 21904
rect 28736 21690 28764 21898
rect 28724 21684 28776 21690
rect 28724 21626 28776 21632
rect 28920 21486 28948 22034
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28828 21049 28856 21422
rect 28814 21040 28870 21049
rect 28814 20975 28870 20984
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28632 19984 28684 19990
rect 28632 19926 28684 19932
rect 28630 19544 28686 19553
rect 28736 19514 28764 20878
rect 28828 20874 28856 20975
rect 28816 20868 28868 20874
rect 28816 20810 28868 20816
rect 29092 20392 29144 20398
rect 29092 20334 29144 20340
rect 29104 20074 29132 20334
rect 29012 20046 29132 20074
rect 28630 19479 28686 19488
rect 28724 19508 28776 19514
rect 28644 19446 28672 19479
rect 28724 19450 28776 19456
rect 28632 19440 28684 19446
rect 28632 19382 28684 19388
rect 29012 19334 29040 20046
rect 29092 19916 29144 19922
rect 29092 19858 29144 19864
rect 28632 19304 28684 19310
rect 28632 19246 28684 19252
rect 28966 19306 29040 19334
rect 28644 18630 28672 19246
rect 28966 18986 28994 19306
rect 29104 19258 29132 19858
rect 29182 19272 29238 19281
rect 29104 19230 29182 19258
rect 29182 19207 29238 19216
rect 29092 19168 29144 19174
rect 29092 19110 29144 19116
rect 28736 18958 28994 18986
rect 28632 18624 28684 18630
rect 28632 18566 28684 18572
rect 28460 17054 28580 17082
rect 28460 16522 28488 17054
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 28184 16204 28396 16232
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27816 15026 27844 16118
rect 28184 15502 28212 16204
rect 28264 16108 28316 16114
rect 28460 16096 28488 16458
rect 28316 16068 28488 16096
rect 28264 16050 28316 16056
rect 28552 16028 28580 16730
rect 28644 16130 28672 18566
rect 28736 16794 28764 18958
rect 28920 18834 29040 18850
rect 28908 18828 29040 18834
rect 28960 18822 29040 18828
rect 28908 18770 28960 18776
rect 29012 18737 29040 18822
rect 28998 18728 29054 18737
rect 28998 18663 29054 18672
rect 29104 18601 29132 19110
rect 29182 18864 29238 18873
rect 29182 18799 29238 18808
rect 29196 18630 29224 18799
rect 29184 18624 29236 18630
rect 29090 18592 29146 18601
rect 29184 18566 29236 18572
rect 29090 18527 29146 18536
rect 28908 18216 28960 18222
rect 28908 18158 28960 18164
rect 28920 18086 28948 18158
rect 29288 18154 29316 23462
rect 29748 23322 29776 23530
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 29380 21865 29408 22918
rect 29460 22704 29512 22710
rect 29460 22646 29512 22652
rect 29366 21856 29422 21865
rect 29366 21791 29422 21800
rect 29472 21536 29500 22646
rect 29734 22264 29790 22273
rect 29734 22199 29790 22208
rect 29748 22166 29776 22199
rect 29736 22160 29788 22166
rect 29736 22102 29788 22108
rect 29550 21992 29606 22001
rect 29550 21927 29606 21936
rect 29380 21508 29500 21536
rect 29380 20330 29408 21508
rect 29460 21412 29512 21418
rect 29460 21354 29512 21360
rect 29472 20398 29500 21354
rect 29460 20392 29512 20398
rect 29460 20334 29512 20340
rect 29368 20324 29420 20330
rect 29368 20266 29420 20272
rect 29564 20074 29592 21927
rect 29644 21888 29696 21894
rect 29644 21830 29696 21836
rect 29656 20534 29684 21830
rect 29840 21622 29868 23530
rect 29932 23322 29960 26200
rect 30576 24682 30604 26200
rect 30380 24676 30432 24682
rect 30380 24618 30432 24624
rect 30564 24676 30616 24682
rect 30564 24618 30616 24624
rect 30196 24404 30248 24410
rect 30196 24346 30248 24352
rect 29920 23316 29972 23322
rect 29920 23258 29972 23264
rect 30208 23186 30236 24346
rect 30392 24290 30420 24618
rect 30564 24336 30616 24342
rect 30392 24284 30564 24290
rect 30392 24278 30616 24284
rect 30392 24262 30604 24278
rect 30392 24206 30420 24262
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23186 30328 23462
rect 30196 23180 30248 23186
rect 30196 23122 30248 23128
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30012 22704 30064 22710
rect 30012 22646 30064 22652
rect 30024 22506 30052 22646
rect 30012 22500 30064 22506
rect 30012 22442 30064 22448
rect 29918 22128 29974 22137
rect 29918 22063 29974 22072
rect 29932 22030 29960 22063
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29828 21616 29880 21622
rect 29828 21558 29880 21564
rect 29734 21176 29790 21185
rect 29734 21111 29736 21120
rect 29788 21111 29790 21120
rect 29736 21082 29788 21088
rect 29644 20528 29696 20534
rect 29644 20470 29696 20476
rect 29472 20046 29592 20074
rect 29472 19990 29500 20046
rect 29460 19984 29512 19990
rect 29380 19944 29460 19972
rect 29380 19310 29408 19944
rect 29460 19926 29512 19932
rect 29550 19952 29606 19961
rect 29550 19887 29606 19896
rect 29564 19357 29592 19887
rect 29644 19712 29696 19718
rect 29644 19654 29696 19660
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29550 19348 29606 19357
rect 29368 19304 29420 19310
rect 29550 19283 29606 19292
rect 29368 19246 29420 19252
rect 29656 19242 29684 19654
rect 29748 19357 29776 19654
rect 29734 19348 29790 19357
rect 29734 19283 29790 19292
rect 29460 19236 29512 19242
rect 29460 19178 29512 19184
rect 29644 19236 29696 19242
rect 29840 19224 29868 21558
rect 30116 21078 30144 22918
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30208 22098 30236 22374
rect 30196 22092 30248 22098
rect 30196 22034 30248 22040
rect 30392 22030 30420 22510
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 30380 22024 30432 22030
rect 30380 21966 30432 21972
rect 30484 21962 30512 22374
rect 30472 21956 30524 21962
rect 30472 21898 30524 21904
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30288 21480 30340 21486
rect 30288 21422 30340 21428
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30104 21072 30156 21078
rect 30104 21014 30156 21020
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29932 19334 29960 20878
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30024 19718 30052 20742
rect 30116 20398 30144 20742
rect 30104 20392 30156 20398
rect 30104 20334 30156 20340
rect 30104 19848 30156 19854
rect 30102 19816 30104 19825
rect 30156 19816 30158 19825
rect 30102 19751 30158 19760
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 30208 19394 30236 21286
rect 30300 20330 30328 21422
rect 30392 20856 30420 21830
rect 30576 21690 30604 24006
rect 31024 23792 31076 23798
rect 31024 23734 31076 23740
rect 31036 23662 31064 23734
rect 31024 23656 31076 23662
rect 31024 23598 31076 23604
rect 31036 23186 31064 23598
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 30748 22976 30800 22982
rect 30748 22918 30800 22924
rect 30760 22642 30788 22918
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30748 22636 30800 22642
rect 30748 22578 30800 22584
rect 30668 22545 30696 22578
rect 30654 22536 30710 22545
rect 30654 22471 30710 22480
rect 30656 22228 30708 22234
rect 30656 22170 30708 22176
rect 30564 21684 30616 21690
rect 30564 21626 30616 21632
rect 30564 21412 30616 21418
rect 30564 21354 30616 21360
rect 30576 20913 30604 21354
rect 30668 21146 30696 22170
rect 30760 21894 30788 22578
rect 30852 22438 30880 22714
rect 30840 22432 30892 22438
rect 30840 22374 30892 22380
rect 30840 22024 30892 22030
rect 30840 21966 30892 21972
rect 30748 21888 30800 21894
rect 30748 21830 30800 21836
rect 30748 21480 30800 21486
rect 30748 21422 30800 21428
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30562 20904 30618 20913
rect 30472 20868 30524 20874
rect 30392 20828 30472 20856
rect 30562 20839 30618 20848
rect 30472 20810 30524 20816
rect 30288 20324 30340 20330
rect 30288 20266 30340 20272
rect 30378 19816 30434 19825
rect 30484 19786 30512 20810
rect 30656 20392 30708 20398
rect 30656 20334 30708 20340
rect 30564 20256 30616 20262
rect 30564 20198 30616 20204
rect 30378 19751 30380 19760
rect 30432 19751 30434 19760
rect 30472 19780 30524 19786
rect 30380 19722 30432 19728
rect 30472 19722 30524 19728
rect 30288 19712 30340 19718
rect 30288 19654 30340 19660
rect 30116 19366 30236 19394
rect 30300 19378 30328 19654
rect 30288 19372 30340 19378
rect 29932 19315 30052 19334
rect 29932 19306 30066 19315
rect 30010 19241 30066 19250
rect 29840 19196 29960 19224
rect 29644 19178 29696 19184
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29000 18148 29052 18154
rect 29000 18090 29052 18096
rect 29276 18148 29328 18154
rect 29276 18090 29328 18096
rect 28908 18080 28960 18086
rect 28908 18022 28960 18028
rect 28906 17912 28962 17921
rect 28906 17847 28962 17856
rect 28920 17814 28948 17847
rect 28908 17808 28960 17814
rect 28908 17750 28960 17756
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28814 16960 28870 16969
rect 28814 16895 28870 16904
rect 28724 16788 28776 16794
rect 28724 16730 28776 16736
rect 28644 16102 28764 16130
rect 28632 16040 28684 16046
rect 28552 16000 28632 16028
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 27804 14476 27856 14482
rect 27724 14436 27804 14464
rect 27804 14418 27856 14424
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27436 13728 27488 13734
rect 27436 13670 27488 13676
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 26884 12164 26936 12170
rect 26884 12106 26936 12112
rect 27068 12164 27120 12170
rect 27068 12106 27120 12112
rect 26976 11824 27028 11830
rect 26976 11766 27028 11772
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 25596 11008 25648 11014
rect 25596 10950 25648 10956
rect 26332 10804 26384 10810
rect 26332 10746 26384 10752
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 26068 9994 26096 10406
rect 26344 10266 26372 10746
rect 26620 10606 26648 11290
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26712 10674 26740 11018
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26620 10198 26648 10542
rect 26712 10470 26740 10610
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26608 10192 26660 10198
rect 26608 10134 26660 10140
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 25056 9178 25084 9862
rect 26068 9722 26096 9930
rect 26712 9926 26740 10406
rect 26896 10130 26924 11086
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 26712 9722 26740 9862
rect 26056 9716 26108 9722
rect 26056 9658 26108 9664
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24044 8498 24072 8978
rect 25792 8838 25820 9386
rect 25976 8974 26004 9454
rect 25964 8968 26016 8974
rect 25962 8936 25964 8945
rect 26016 8936 26018 8945
rect 25962 8871 26018 8880
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24872 8362 24900 8774
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 25792 7750 25820 8774
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 25792 4826 25820 7686
rect 26988 6254 27016 11766
rect 27172 11082 27200 12242
rect 27632 12238 27660 14010
rect 27724 13190 27752 14282
rect 27816 14074 27844 14418
rect 28092 14414 28120 14758
rect 28552 14550 28580 16000
rect 28632 15982 28684 15988
rect 28540 14544 28592 14550
rect 28540 14486 28592 14492
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 28448 13796 28500 13802
rect 28448 13738 28500 13744
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27528 12164 27580 12170
rect 27528 12106 27580 12112
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27356 11898 27384 12038
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 27068 10804 27120 10810
rect 27068 10746 27120 10752
rect 27080 6322 27108 10746
rect 27172 9518 27200 11018
rect 27264 9994 27292 11494
rect 27344 10736 27396 10742
rect 27344 10678 27396 10684
rect 27356 10606 27384 10678
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27448 10470 27476 11630
rect 27436 10464 27488 10470
rect 27436 10406 27488 10412
rect 27252 9988 27304 9994
rect 27252 9930 27304 9936
rect 27264 9654 27292 9930
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 27540 8022 27568 12106
rect 27724 10169 27752 13126
rect 27816 11626 27844 13262
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27804 11620 27856 11626
rect 27804 11562 27856 11568
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27710 10160 27766 10169
rect 27710 10095 27766 10104
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27816 6390 27844 8774
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27068 6316 27120 6322
rect 27068 6258 27120 6264
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 28368 6186 28396 13466
rect 28460 13258 28488 13738
rect 28448 13252 28500 13258
rect 28448 13194 28500 13200
rect 28460 12918 28488 13194
rect 28552 13190 28580 14486
rect 28632 14408 28684 14414
rect 28736 14396 28764 16102
rect 28828 15706 28856 16895
rect 28920 16590 28948 17614
rect 29012 16590 29040 18090
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29184 17808 29236 17814
rect 29184 17750 29236 17756
rect 29196 17610 29224 17750
rect 29184 17604 29236 17610
rect 29184 17546 29236 17552
rect 29092 17536 29144 17542
rect 29092 17478 29144 17484
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 29000 16584 29052 16590
rect 29000 16526 29052 16532
rect 28920 16182 28948 16526
rect 29104 16182 29132 17478
rect 28908 16176 28960 16182
rect 28908 16118 28960 16124
rect 29092 16176 29144 16182
rect 29092 16118 29144 16124
rect 29104 15706 29132 16118
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 28828 15434 28856 15642
rect 28816 15428 28868 15434
rect 28816 15370 28868 15376
rect 29000 15088 29052 15094
rect 29104 15076 29132 15642
rect 29052 15048 29132 15076
rect 29000 15030 29052 15036
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28684 14368 28764 14396
rect 28632 14350 28684 14356
rect 28540 13184 28592 13190
rect 28538 13152 28540 13161
rect 28592 13152 28594 13161
rect 28538 13087 28594 13096
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28448 12912 28500 12918
rect 28448 12854 28500 12860
rect 28460 11830 28488 12854
rect 28448 11824 28500 11830
rect 28448 11766 28500 11772
rect 28552 11354 28580 12922
rect 28644 12753 28672 14350
rect 28828 14006 28856 14758
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28816 14000 28868 14006
rect 28816 13942 28868 13948
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 28920 13530 28948 13874
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 29012 13326 29040 14214
rect 29104 13802 29132 15048
rect 29288 14890 29316 17818
rect 29380 16794 29408 18634
rect 29368 16788 29420 16794
rect 29472 16776 29500 19178
rect 29550 19136 29606 19145
rect 29550 19071 29606 19080
rect 29564 17882 29592 19071
rect 29642 19000 29698 19009
rect 29932 18952 29960 19196
rect 29642 18935 29698 18944
rect 29656 18834 29684 18935
rect 29840 18924 29960 18952
rect 30012 18964 30064 18970
rect 29644 18828 29696 18834
rect 29644 18770 29696 18776
rect 29642 18728 29698 18737
rect 29840 18698 29868 18924
rect 30012 18906 30064 18912
rect 29920 18828 29972 18834
rect 29920 18770 29972 18776
rect 29642 18663 29698 18672
rect 29828 18692 29880 18698
rect 29656 18630 29684 18663
rect 29828 18634 29880 18640
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29644 18080 29696 18086
rect 29644 18022 29696 18028
rect 29552 17876 29604 17882
rect 29552 17818 29604 17824
rect 29564 17270 29592 17818
rect 29552 17264 29604 17270
rect 29552 17206 29604 17212
rect 29472 16748 29592 16776
rect 29368 16730 29420 16736
rect 29460 16652 29512 16658
rect 29460 16594 29512 16600
rect 29368 16448 29420 16454
rect 29368 16390 29420 16396
rect 29380 16017 29408 16390
rect 29366 16008 29422 16017
rect 29366 15943 29422 15952
rect 29276 14884 29328 14890
rect 29276 14826 29328 14832
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 29092 13796 29144 13802
rect 29092 13738 29144 13744
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28814 13152 28870 13161
rect 28630 12744 28686 12753
rect 28630 12679 28686 12688
rect 28632 11892 28684 11898
rect 28736 11880 28764 13126
rect 28814 13087 28870 13096
rect 28828 12646 28856 13087
rect 28816 12640 28868 12646
rect 28816 12582 28868 12588
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28684 11852 28764 11880
rect 28632 11834 28684 11840
rect 28828 11694 28856 12174
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 28828 11354 28856 11630
rect 28908 11620 28960 11626
rect 28908 11562 28960 11568
rect 28540 11348 28592 11354
rect 28816 11348 28868 11354
rect 28540 11290 28592 11296
rect 28736 11308 28816 11336
rect 28540 11076 28592 11082
rect 28540 11018 28592 11024
rect 28552 9994 28580 11018
rect 28736 10810 28764 11308
rect 28816 11290 28868 11296
rect 28920 11098 28948 11562
rect 29288 11132 29316 14418
rect 29380 14278 29408 15943
rect 29368 14272 29420 14278
rect 29368 14214 29420 14220
rect 29380 12918 29408 14214
rect 29368 12912 29420 12918
rect 29368 12854 29420 12860
rect 29472 11200 29500 16594
rect 29564 15706 29592 16748
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29552 15020 29604 15026
rect 29552 14962 29604 14968
rect 29564 14822 29592 14962
rect 29552 14816 29604 14822
rect 29552 14758 29604 14764
rect 29656 14482 29684 18022
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 29748 14958 29776 17070
rect 29828 16040 29880 16046
rect 29828 15982 29880 15988
rect 29840 15162 29868 15982
rect 29828 15156 29880 15162
rect 29828 15098 29880 15104
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29644 14476 29696 14482
rect 29644 14418 29696 14424
rect 29748 13258 29776 14894
rect 29840 14226 29868 15098
rect 29932 14958 29960 18770
rect 30024 18154 30052 18906
rect 30116 18290 30144 19366
rect 30288 19314 30340 19320
rect 30380 19304 30432 19310
rect 30380 19246 30432 19252
rect 30288 19236 30340 19242
rect 30288 19178 30340 19184
rect 30194 19136 30250 19145
rect 30194 19071 30250 19080
rect 30208 18426 30236 19071
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30104 18284 30156 18290
rect 30104 18226 30156 18232
rect 30300 18222 30328 19178
rect 30288 18216 30340 18222
rect 30288 18158 30340 18164
rect 30012 18148 30064 18154
rect 30012 18090 30064 18096
rect 30024 16658 30052 18090
rect 30392 17610 30420 19246
rect 30472 18624 30524 18630
rect 30472 18566 30524 18572
rect 30104 17604 30156 17610
rect 30104 17546 30156 17552
rect 30380 17604 30432 17610
rect 30380 17546 30432 17552
rect 30116 17513 30144 17546
rect 30102 17504 30158 17513
rect 30102 17439 30158 17448
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30116 16794 30144 17070
rect 30288 17060 30340 17066
rect 30288 17002 30340 17008
rect 30196 16992 30248 16998
rect 30196 16934 30248 16940
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30208 16697 30236 16934
rect 30194 16688 30250 16697
rect 30012 16652 30064 16658
rect 30194 16623 30250 16632
rect 30012 16594 30064 16600
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 30012 15360 30064 15366
rect 30012 15302 30064 15308
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 30024 14414 30052 15302
rect 30012 14408 30064 14414
rect 30012 14350 30064 14356
rect 30116 14278 30144 15438
rect 30300 15366 30328 17002
rect 30392 16250 30420 17070
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30484 15586 30512 18566
rect 30576 17202 30604 20198
rect 30668 17338 30696 20334
rect 30760 19009 30788 21422
rect 30852 20602 30880 21966
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 30944 20874 30972 21490
rect 31036 21146 31064 23122
rect 31024 21140 31076 21146
rect 31024 21082 31076 21088
rect 31128 21026 31156 24006
rect 31220 22982 31248 26200
rect 31864 24614 31892 26200
rect 32508 24721 32536 26200
rect 32864 24744 32916 24750
rect 32494 24712 32550 24721
rect 32864 24686 32916 24692
rect 32494 24647 32550 24656
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31300 24336 31352 24342
rect 31300 24278 31352 24284
rect 31312 23254 31340 24278
rect 31576 24268 31628 24274
rect 31576 24210 31628 24216
rect 32772 24268 32824 24274
rect 32772 24210 32824 24216
rect 31392 23792 31444 23798
rect 31588 23780 31616 24210
rect 32312 24064 32364 24070
rect 32312 24006 32364 24012
rect 31444 23752 31616 23780
rect 31392 23734 31444 23740
rect 31760 23656 31812 23662
rect 31760 23598 31812 23604
rect 31300 23248 31352 23254
rect 31300 23190 31352 23196
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 31312 22624 31340 23190
rect 31772 23186 31800 23598
rect 32324 23526 32352 24006
rect 32496 23792 32548 23798
rect 32496 23734 32548 23740
rect 32312 23520 32364 23526
rect 32312 23462 32364 23468
rect 31668 23180 31720 23186
rect 31588 23140 31668 23168
rect 31482 22672 31538 22681
rect 31312 22596 31432 22624
rect 31482 22607 31538 22616
rect 31208 22500 31260 22506
rect 31208 22442 31260 22448
rect 31220 22001 31248 22442
rect 31404 22250 31432 22596
rect 31496 22438 31524 22607
rect 31484 22432 31536 22438
rect 31484 22374 31536 22380
rect 31404 22234 31524 22250
rect 31404 22228 31536 22234
rect 31404 22222 31484 22228
rect 31484 22170 31536 22176
rect 31588 22098 31616 23140
rect 31668 23122 31720 23128
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 31668 22228 31720 22234
rect 31668 22170 31720 22176
rect 31576 22092 31628 22098
rect 31576 22034 31628 22040
rect 31588 22003 31616 22034
rect 31206 21992 31262 22001
rect 31206 21927 31208 21936
rect 31260 21927 31262 21936
rect 31208 21898 31260 21904
rect 31206 21720 31262 21729
rect 31206 21655 31208 21664
rect 31260 21655 31262 21664
rect 31208 21626 31260 21632
rect 31036 20998 31156 21026
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 31036 20754 31064 20998
rect 31390 20904 31446 20913
rect 31390 20839 31446 20848
rect 30944 20726 31064 20754
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30746 19000 30802 19009
rect 30746 18935 30802 18944
rect 30746 18864 30802 18873
rect 30746 18799 30802 18808
rect 30760 18698 30788 18799
rect 30748 18692 30800 18698
rect 30748 18634 30800 18640
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30656 17332 30708 17338
rect 30656 17274 30708 17280
rect 30760 17218 30788 18022
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30668 17190 30788 17218
rect 30564 16720 30616 16726
rect 30564 16662 30616 16668
rect 30576 16028 30604 16662
rect 30668 16182 30696 17190
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 30656 16176 30708 16182
rect 30656 16118 30708 16124
rect 30576 16000 30696 16028
rect 30392 15558 30512 15586
rect 30288 15360 30340 15366
rect 30288 15302 30340 15308
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30104 14272 30156 14278
rect 29840 14198 29960 14226
rect 30104 14214 30156 14220
rect 29932 13462 29960 14198
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 29920 13456 29972 13462
rect 29920 13398 29972 13404
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29736 13252 29788 13258
rect 29736 13194 29788 13200
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29656 11370 29684 12718
rect 29748 11801 29776 12854
rect 29734 11792 29790 11801
rect 29734 11727 29790 11736
rect 29656 11342 29776 11370
rect 29472 11172 29684 11200
rect 29368 11144 29420 11150
rect 29288 11104 29368 11132
rect 28920 11082 29040 11098
rect 29368 11086 29420 11092
rect 28908 11076 29040 11082
rect 28960 11070 29040 11076
rect 28908 11018 28960 11024
rect 29012 11014 29040 11070
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 29012 10198 29040 10950
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29000 10192 29052 10198
rect 28630 10160 28686 10169
rect 29000 10134 29052 10140
rect 28630 10095 28686 10104
rect 28540 9988 28592 9994
rect 28540 9930 28592 9936
rect 28644 7274 28672 10095
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28736 9722 28764 9930
rect 28724 9716 28776 9722
rect 28724 9658 28776 9664
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28828 8430 28856 9318
rect 29104 8566 29132 10202
rect 29380 10198 29408 11086
rect 29460 11076 29512 11082
rect 29460 11018 29512 11024
rect 29472 10606 29500 11018
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29564 10606 29592 10678
rect 29460 10600 29512 10606
rect 29460 10542 29512 10548
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29368 10192 29420 10198
rect 29368 10134 29420 10140
rect 29564 10130 29592 10542
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 29564 9518 29592 10066
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29288 9382 29316 9454
rect 29656 9450 29684 11172
rect 29748 10674 29776 11342
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29840 10606 29868 13330
rect 29932 12170 29960 13398
rect 30024 12850 30052 14010
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 30024 12306 30052 12786
rect 30116 12345 30144 14214
rect 30208 13326 30236 14758
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30300 13172 30328 14894
rect 30392 13394 30420 15558
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30484 15162 30512 15370
rect 30472 15156 30524 15162
rect 30472 15098 30524 15104
rect 30484 14822 30512 15098
rect 30472 14816 30524 14822
rect 30472 14758 30524 14764
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30576 14278 30604 14554
rect 30668 14482 30696 16000
rect 30760 15910 30788 17070
rect 30852 16182 30880 20198
rect 30944 20058 30972 20726
rect 31022 20496 31078 20505
rect 31022 20431 31078 20440
rect 30932 20052 30984 20058
rect 30932 19994 30984 20000
rect 31036 19854 31064 20431
rect 30932 19848 30984 19854
rect 30932 19790 30984 19796
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 30944 18970 30972 19790
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 30944 18465 30972 18906
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 30930 18456 30986 18465
rect 30930 18391 30986 18400
rect 31036 16590 31064 18566
rect 31220 18426 31248 20742
rect 31300 19712 31352 19718
rect 31300 19654 31352 19660
rect 31312 18630 31340 19654
rect 31404 19514 31432 20839
rect 31680 20618 31708 22170
rect 32220 22024 32272 22030
rect 31850 21992 31906 22001
rect 31772 21950 31850 21978
rect 31772 20874 31800 21950
rect 32220 21966 32272 21972
rect 31850 21927 31906 21936
rect 31760 20868 31812 20874
rect 31760 20810 31812 20816
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31484 20596 31536 20602
rect 31484 20538 31536 20544
rect 31588 20590 31708 20618
rect 31392 19508 31444 19514
rect 31392 19450 31444 19456
rect 31496 19446 31524 20538
rect 31588 20534 31616 20590
rect 31576 20528 31628 20534
rect 31668 20528 31720 20534
rect 31576 20470 31628 20476
rect 31666 20496 31668 20505
rect 31720 20496 31722 20505
rect 31666 20431 31722 20440
rect 31576 20052 31628 20058
rect 31576 19994 31628 20000
rect 31484 19440 31536 19446
rect 31484 19382 31536 19388
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31484 17740 31536 17746
rect 31484 17682 31536 17688
rect 31392 17672 31444 17678
rect 31114 17640 31170 17649
rect 31392 17614 31444 17620
rect 31114 17575 31170 17584
rect 31128 16658 31156 17575
rect 31404 17338 31432 17614
rect 31392 17332 31444 17338
rect 31392 17274 31444 17280
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30760 15434 30788 15846
rect 31116 15564 31168 15570
rect 31116 15506 31168 15512
rect 30748 15428 30800 15434
rect 30748 15370 30800 15376
rect 30656 14476 30708 14482
rect 30760 14464 30788 15370
rect 30840 14476 30892 14482
rect 30760 14436 30840 14464
rect 30656 14418 30708 14424
rect 30840 14418 30892 14424
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 31128 14074 31156 15506
rect 31312 15162 31340 16390
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31404 14618 31432 15846
rect 31392 14612 31444 14618
rect 31392 14554 31444 14560
rect 31496 14482 31524 17682
rect 31588 17592 31616 19994
rect 31772 19446 31800 20810
rect 31864 20398 31892 20810
rect 32232 20806 32260 21966
rect 32508 21894 32536 23734
rect 32784 23730 32812 24210
rect 32876 24206 32904 24686
rect 33152 24596 33180 26200
rect 33152 24568 33456 24596
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 33048 24336 33100 24342
rect 33048 24278 33100 24284
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32772 23724 32824 23730
rect 32772 23666 32824 23672
rect 32692 21894 32720 23666
rect 32784 23118 32812 23666
rect 32876 23254 32904 24142
rect 33060 23798 33088 24278
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 33048 23792 33100 23798
rect 33048 23734 33100 23740
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33336 23322 33364 24142
rect 33428 23361 33456 24568
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33598 23488 33654 23497
rect 33598 23423 33654 23432
rect 33414 23352 33470 23361
rect 33324 23316 33376 23322
rect 33414 23287 33470 23296
rect 33324 23258 33376 23264
rect 32864 23248 32916 23254
rect 32864 23190 32916 23196
rect 33324 23180 33376 23186
rect 33324 23122 33376 23128
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 33232 23044 33284 23050
rect 33232 22986 33284 22992
rect 33244 22778 33272 22986
rect 33232 22772 33284 22778
rect 33232 22714 33284 22720
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32772 22092 32824 22098
rect 32772 22034 32824 22040
rect 32496 21888 32548 21894
rect 32416 21848 32496 21876
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 32232 20534 32260 20742
rect 32220 20528 32272 20534
rect 32220 20470 32272 20476
rect 32324 20398 32352 20946
rect 32416 20942 32444 21848
rect 32496 21830 32548 21836
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32588 21616 32640 21622
rect 32588 21558 32640 21564
rect 32404 20936 32456 20942
rect 32404 20878 32456 20884
rect 32496 20936 32548 20942
rect 32496 20878 32548 20884
rect 32508 20602 32536 20878
rect 32496 20596 32548 20602
rect 32496 20538 32548 20544
rect 32600 20398 32628 21558
rect 31852 20392 31904 20398
rect 31944 20392 31996 20398
rect 31852 20334 31904 20340
rect 31942 20360 31944 20369
rect 32312 20392 32364 20398
rect 31996 20360 31998 20369
rect 32312 20334 32364 20340
rect 32588 20392 32640 20398
rect 32588 20334 32640 20340
rect 31942 20295 31998 20304
rect 32784 20058 32812 22034
rect 32862 21856 32918 21865
rect 32862 21791 32918 21800
rect 33230 21856 33286 21865
rect 33230 21791 33286 21800
rect 32876 21049 32904 21791
rect 33244 21593 33272 21791
rect 33230 21584 33286 21593
rect 33230 21519 33286 21528
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32862 21040 32918 21049
rect 32862 20975 32918 20984
rect 32876 20874 32904 20975
rect 32864 20868 32916 20874
rect 32864 20810 32916 20816
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32772 20052 32824 20058
rect 32772 19994 32824 20000
rect 32772 19916 32824 19922
rect 32772 19858 32824 19864
rect 32784 19802 32812 19858
rect 32312 19780 32364 19786
rect 32692 19774 32812 19802
rect 32692 19768 32720 19774
rect 32364 19740 32720 19768
rect 32312 19722 32364 19728
rect 33336 19718 33364 23122
rect 33612 22710 33640 23423
rect 33888 23202 33916 24142
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 34072 23633 34100 24006
rect 34058 23624 34114 23633
rect 34058 23559 34114 23568
rect 34256 23225 34284 26302
rect 34426 26200 34482 26302
rect 35070 26200 35126 27000
rect 35714 26330 35770 27000
rect 35714 26302 35848 26330
rect 35714 26200 35770 26302
rect 34980 24744 35032 24750
rect 34980 24686 35032 24692
rect 34992 24274 35020 24686
rect 34336 24268 34388 24274
rect 34336 24210 34388 24216
rect 34980 24268 35032 24274
rect 34980 24210 35032 24216
rect 33796 23186 33916 23202
rect 33784 23180 33916 23186
rect 33836 23174 33916 23180
rect 33784 23122 33836 23128
rect 33784 22976 33836 22982
rect 33784 22918 33836 22924
rect 33600 22704 33652 22710
rect 33600 22646 33652 22652
rect 33692 22500 33744 22506
rect 33692 22442 33744 22448
rect 33704 22409 33732 22442
rect 33690 22400 33746 22409
rect 33690 22335 33746 22344
rect 33692 21956 33744 21962
rect 33692 21898 33744 21904
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33428 21690 33456 21830
rect 33598 21720 33654 21729
rect 33416 21684 33468 21690
rect 33598 21655 33600 21664
rect 33416 21626 33468 21632
rect 33652 21655 33654 21664
rect 33600 21626 33652 21632
rect 33506 21584 33562 21593
rect 33704 21554 33732 21898
rect 33506 21519 33508 21528
rect 33560 21519 33562 21528
rect 33692 21548 33744 21554
rect 33508 21490 33560 21496
rect 33692 21490 33744 21496
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 33416 20392 33468 20398
rect 33416 20334 33468 20340
rect 32128 19712 32180 19718
rect 32128 19654 32180 19660
rect 33324 19712 33376 19718
rect 33324 19654 33376 19660
rect 31760 19440 31812 19446
rect 31760 19382 31812 19388
rect 31760 19168 31812 19174
rect 31760 19110 31812 19116
rect 31772 17678 31800 19110
rect 31852 18624 31904 18630
rect 31852 18566 31904 18572
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31668 17604 31720 17610
rect 31588 17564 31668 17592
rect 31668 17546 31720 17552
rect 31576 17060 31628 17066
rect 31576 17002 31628 17008
rect 31208 14476 31260 14482
rect 31208 14418 31260 14424
rect 31484 14476 31536 14482
rect 31484 14418 31536 14424
rect 31116 14068 31168 14074
rect 31116 14010 31168 14016
rect 31128 13938 31156 14010
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 30840 13728 30892 13734
rect 30840 13670 30892 13676
rect 30380 13388 30432 13394
rect 30380 13330 30432 13336
rect 30208 13144 30328 13172
rect 30102 12336 30158 12345
rect 30012 12300 30064 12306
rect 30102 12271 30158 12280
rect 30012 12242 30064 12248
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 30116 11778 30144 12271
rect 30024 11750 30144 11778
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 29828 10600 29880 10606
rect 29828 10542 29880 10548
rect 29840 10266 29868 10542
rect 29828 10260 29880 10266
rect 29828 10202 29880 10208
rect 29644 9444 29696 9450
rect 29644 9386 29696 9392
rect 29276 9376 29328 9382
rect 29276 9318 29328 9324
rect 29656 9110 29684 9386
rect 29644 9104 29696 9110
rect 29644 9046 29696 9052
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 28632 7268 28684 7274
rect 28632 7210 28684 7216
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 26148 4752 26200 4758
rect 26148 4694 26200 4700
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 21008 2990 21036 3470
rect 21284 3058 21312 4422
rect 22112 4214 22140 4558
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22112 3618 22140 4150
rect 23216 4146 23244 4558
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22112 3590 22232 3618
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 22204 2922 22232 3590
rect 22848 3534 22876 3878
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23308 3738 23336 4014
rect 23584 3738 23612 4626
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24780 4214 24808 4422
rect 24768 4208 24820 4214
rect 24768 4150 24820 4156
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20180 800 20208 2450
rect 22112 2446 22140 2858
rect 22296 2854 22324 3334
rect 22756 2922 22784 3334
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 23308 2854 23336 3674
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23768 3058 23796 3470
rect 24584 3188 24636 3194
rect 24584 3130 24636 3136
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22296 800 22324 2450
rect 24412 800 24440 2450
rect 24596 2446 24624 3130
rect 24872 2582 24900 4014
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 25976 3194 26004 3674
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 26160 3058 26188 4694
rect 28724 4548 28776 4554
rect 28724 4490 28776 4496
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27804 4072 27856 4078
rect 27896 4072 27948 4078
rect 27804 4014 27856 4020
rect 27894 4040 27896 4049
rect 27948 4040 27950 4049
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26528 3398 26556 3470
rect 26516 3392 26568 3398
rect 26516 3334 26568 3340
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 26528 2990 26556 3334
rect 27540 3194 27568 3878
rect 27816 3194 27844 4014
rect 27894 3975 27950 3984
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 28368 3398 28396 3538
rect 28356 3392 28408 3398
rect 28356 3334 28408 3340
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 28368 3058 28396 3334
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 28736 2990 28764 4490
rect 28828 3058 28856 8366
rect 29932 7954 29960 10746
rect 30024 10198 30052 11750
rect 30208 11558 30236 13144
rect 30562 12880 30618 12889
rect 30562 12815 30618 12824
rect 30288 11688 30340 11694
rect 30288 11630 30340 11636
rect 30470 11656 30526 11665
rect 30196 11552 30248 11558
rect 30196 11494 30248 11500
rect 30196 11212 30248 11218
rect 30196 11154 30248 11160
rect 30012 10192 30064 10198
rect 30012 10134 30064 10140
rect 30208 9722 30236 11154
rect 30300 11150 30328 11630
rect 30470 11591 30526 11600
rect 30484 11354 30512 11591
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30300 10742 30328 11086
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30392 10266 30420 11018
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30380 10260 30432 10266
rect 30380 10202 30432 10208
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 30116 9518 30144 9590
rect 30104 9512 30156 9518
rect 30104 9454 30156 9460
rect 30484 9382 30512 10542
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30196 9036 30248 9042
rect 30196 8978 30248 8984
rect 30208 8838 30236 8978
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 30484 7750 30512 8570
rect 30576 8090 30604 12815
rect 30852 11694 30880 13670
rect 31024 12368 31076 12374
rect 31024 12310 31076 12316
rect 30840 11688 30892 11694
rect 30840 11630 30892 11636
rect 31036 11286 31064 12310
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31128 11898 31156 12174
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 31024 11280 31076 11286
rect 31024 11222 31076 11228
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 30668 10130 30696 10610
rect 30746 10568 30802 10577
rect 30746 10503 30802 10512
rect 30760 10470 30788 10503
rect 30748 10464 30800 10470
rect 30748 10406 30800 10412
rect 30656 10124 30708 10130
rect 30656 10066 30708 10072
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30760 9654 30788 9998
rect 30748 9648 30800 9654
rect 30748 9590 30800 9596
rect 30760 8838 30788 9590
rect 30748 8832 30800 8838
rect 30748 8774 30800 8780
rect 30760 8566 30788 8774
rect 30748 8560 30800 8566
rect 30748 8502 30800 8508
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 30576 7886 30604 8026
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30760 7818 30788 8502
rect 30748 7812 30800 7818
rect 30748 7754 30800 7760
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30484 7410 30512 7686
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30484 7002 30512 7346
rect 30472 6996 30524 7002
rect 30472 6938 30524 6944
rect 30852 6390 30880 10950
rect 31128 10810 31156 11698
rect 31220 11098 31248 14418
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31496 13326 31524 13874
rect 31588 13394 31616 17002
rect 31760 16992 31812 16998
rect 31760 16934 31812 16940
rect 31772 16250 31800 16934
rect 31864 16454 31892 18566
rect 32140 18358 32168 19654
rect 32864 19508 32916 19514
rect 32864 19450 32916 19456
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 32680 19304 32732 19310
rect 32680 19246 32732 19252
rect 32770 19272 32826 19281
rect 32128 18352 32180 18358
rect 32128 18294 32180 18300
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 32048 17524 32076 18226
rect 32128 17536 32180 17542
rect 32048 17496 32128 17524
rect 32048 17270 32076 17496
rect 32128 17478 32180 17484
rect 32036 17264 32088 17270
rect 32036 17206 32088 17212
rect 31944 16584 31996 16590
rect 31944 16526 31996 16532
rect 31852 16448 31904 16454
rect 31852 16390 31904 16396
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 31956 16046 31984 16526
rect 31944 16040 31996 16046
rect 31944 15982 31996 15988
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31772 15434 31800 15846
rect 31760 15428 31812 15434
rect 31760 15370 31812 15376
rect 31668 15360 31720 15366
rect 31668 15302 31720 15308
rect 31576 13388 31628 13394
rect 31576 13330 31628 13336
rect 31484 13320 31536 13326
rect 31484 13262 31536 13268
rect 31680 13274 31708 15302
rect 31772 13938 31800 15370
rect 31852 14952 31904 14958
rect 31852 14894 31904 14900
rect 31760 13932 31812 13938
rect 31760 13874 31812 13880
rect 31392 12844 31444 12850
rect 31496 12832 31524 13262
rect 31680 13246 31800 13274
rect 31668 13184 31720 13190
rect 31668 13126 31720 13132
rect 31444 12804 31524 12832
rect 31392 12786 31444 12792
rect 31496 12306 31524 12804
rect 31484 12300 31536 12306
rect 31484 12242 31536 12248
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31404 11830 31432 12038
rect 31392 11824 31444 11830
rect 31392 11766 31444 11772
rect 31392 11620 31444 11626
rect 31392 11562 31444 11568
rect 31404 11354 31432 11562
rect 31496 11558 31524 12242
rect 31484 11552 31536 11558
rect 31484 11494 31536 11500
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 31220 11082 31340 11098
rect 31496 11082 31524 11494
rect 31220 11076 31352 11082
rect 31220 11070 31300 11076
rect 31300 11018 31352 11024
rect 31484 11076 31536 11082
rect 31484 11018 31536 11024
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 31496 10742 31524 11018
rect 31576 11008 31628 11014
rect 31576 10950 31628 10956
rect 31484 10736 31536 10742
rect 31484 10678 31536 10684
rect 31588 9722 31616 10950
rect 31576 9716 31628 9722
rect 31576 9658 31628 9664
rect 31484 9648 31536 9654
rect 31484 9590 31536 9596
rect 30930 9072 30986 9081
rect 31496 9042 31524 9590
rect 31588 9466 31616 9658
rect 31680 9586 31708 13126
rect 31772 12986 31800 13246
rect 31760 12980 31812 12986
rect 31760 12922 31812 12928
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31772 12442 31800 12786
rect 31760 12436 31812 12442
rect 31760 12378 31812 12384
rect 31864 11898 31892 14894
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 31760 11688 31812 11694
rect 31760 11630 31812 11636
rect 31772 11506 31800 11630
rect 31772 11478 31892 11506
rect 31864 10470 31892 11478
rect 31760 10464 31812 10470
rect 31760 10406 31812 10412
rect 31852 10464 31904 10470
rect 31852 10406 31904 10412
rect 31772 9761 31800 10406
rect 31758 9752 31814 9761
rect 31864 9722 31892 10406
rect 31956 10248 31984 15982
rect 32048 15366 32076 17206
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 32232 16658 32260 17138
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 32128 16516 32180 16522
rect 32128 16458 32180 16464
rect 32036 15360 32088 15366
rect 32036 15302 32088 15308
rect 32140 12918 32168 16458
rect 32220 16040 32272 16046
rect 32324 16028 32352 19246
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32508 18222 32536 19110
rect 32692 18902 32720 19246
rect 32770 19207 32826 19216
rect 32680 18896 32732 18902
rect 32680 18838 32732 18844
rect 32680 18760 32732 18766
rect 32784 18737 32812 19207
rect 32680 18702 32732 18708
rect 32770 18728 32826 18737
rect 32586 18592 32642 18601
rect 32586 18527 32642 18536
rect 32600 18426 32628 18527
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 32496 18216 32548 18222
rect 32496 18158 32548 18164
rect 32404 17604 32456 17610
rect 32404 17546 32456 17552
rect 32272 16000 32352 16028
rect 32220 15982 32272 15988
rect 32036 12912 32088 12918
rect 32036 12854 32088 12860
rect 32128 12912 32180 12918
rect 32128 12854 32180 12860
rect 32048 12782 32076 12854
rect 32036 12776 32088 12782
rect 32036 12718 32088 12724
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32140 11218 32168 12174
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 32036 10260 32088 10266
rect 31956 10220 32036 10248
rect 32036 10202 32088 10208
rect 31944 9988 31996 9994
rect 31944 9930 31996 9936
rect 31758 9687 31814 9696
rect 31852 9716 31904 9722
rect 31852 9658 31904 9664
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 31956 9518 31984 9930
rect 32048 9926 32076 10202
rect 32140 10130 32168 11154
rect 32232 10606 32260 15982
rect 32312 14476 32364 14482
rect 32312 14418 32364 14424
rect 32324 12646 32352 14418
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32312 12164 32364 12170
rect 32312 12106 32364 12112
rect 32324 11778 32352 12106
rect 32416 11898 32444 17546
rect 32508 17218 32536 18158
rect 32692 17814 32720 18702
rect 32770 18663 32826 18672
rect 32772 18624 32824 18630
rect 32772 18566 32824 18572
rect 32784 18426 32812 18566
rect 32772 18420 32824 18426
rect 32772 18362 32824 18368
rect 32680 17808 32732 17814
rect 32680 17750 32732 17756
rect 32508 17190 32720 17218
rect 32508 16658 32536 17190
rect 32692 17134 32720 17190
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 32680 17128 32732 17134
rect 32680 17070 32732 17076
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32600 16028 32628 17070
rect 32772 16040 32824 16046
rect 32600 16000 32772 16028
rect 32600 15638 32628 16000
rect 32772 15982 32824 15988
rect 32588 15632 32640 15638
rect 32588 15574 32640 15580
rect 32496 14952 32548 14958
rect 32496 14894 32548 14900
rect 32508 13870 32536 14894
rect 32876 14414 32904 19450
rect 33428 19334 33456 20334
rect 33244 19306 33456 19334
rect 33244 19224 33272 19306
rect 33244 19196 33364 19224
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32956 18964 33008 18970
rect 32956 18906 33008 18912
rect 32968 18630 32996 18906
rect 33232 18896 33284 18902
rect 33232 18838 33284 18844
rect 32956 18624 33008 18630
rect 32956 18566 33008 18572
rect 33138 18592 33194 18601
rect 32968 18086 32996 18566
rect 33138 18527 33194 18536
rect 33152 18290 33180 18527
rect 33244 18358 33272 18838
rect 33232 18352 33284 18358
rect 33232 18294 33284 18300
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 32956 18080 33008 18086
rect 32956 18022 33008 18028
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 33336 17746 33364 19196
rect 33416 19168 33468 19174
rect 33520 19156 33548 21286
rect 33692 20800 33744 20806
rect 33692 20742 33744 20748
rect 33704 20398 33732 20742
rect 33692 20392 33744 20398
rect 33692 20334 33744 20340
rect 33600 19916 33652 19922
rect 33600 19858 33652 19864
rect 33612 19718 33640 19858
rect 33600 19712 33652 19718
rect 33600 19654 33652 19660
rect 33600 19304 33652 19310
rect 33600 19246 33652 19252
rect 33468 19128 33548 19156
rect 33416 19110 33468 19116
rect 33612 19009 33640 19246
rect 33704 19174 33732 20334
rect 33796 19854 33824 22918
rect 33888 22710 33916 23174
rect 34242 23216 34298 23225
rect 34242 23151 34298 23160
rect 34244 23112 34296 23118
rect 34244 23054 34296 23060
rect 33876 22704 33928 22710
rect 33876 22646 33928 22652
rect 33968 22432 34020 22438
rect 33968 22374 34020 22380
rect 33980 22098 34008 22374
rect 34256 22234 34284 23054
rect 34348 23050 34376 24210
rect 34428 24132 34480 24138
rect 34428 24074 34480 24080
rect 34336 23044 34388 23050
rect 34336 22986 34388 22992
rect 34440 22574 34468 24074
rect 34980 23656 35032 23662
rect 34980 23598 35032 23604
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34532 23186 34560 23462
rect 34520 23180 34572 23186
rect 34520 23122 34572 23128
rect 34992 23118 35020 23598
rect 35084 23322 35112 26200
rect 35164 24812 35216 24818
rect 35164 24754 35216 24760
rect 35176 24274 35204 24754
rect 35532 24744 35584 24750
rect 35532 24686 35584 24692
rect 35164 24268 35216 24274
rect 35164 24210 35216 24216
rect 35256 24064 35308 24070
rect 35256 24006 35308 24012
rect 35268 23769 35296 24006
rect 35254 23760 35310 23769
rect 35254 23695 35310 23704
rect 35440 23520 35492 23526
rect 35440 23462 35492 23468
rect 35072 23316 35124 23322
rect 35072 23258 35124 23264
rect 34980 23112 35032 23118
rect 34980 23054 35032 23060
rect 34520 22976 34572 22982
rect 34612 22976 34664 22982
rect 34520 22918 34572 22924
rect 34610 22944 34612 22953
rect 34796 22976 34848 22982
rect 34664 22944 34666 22953
rect 34428 22568 34480 22574
rect 34428 22510 34480 22516
rect 34532 22438 34560 22918
rect 34796 22918 34848 22924
rect 34610 22879 34666 22888
rect 34624 22710 34652 22879
rect 34612 22704 34664 22710
rect 34612 22646 34664 22652
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34244 22228 34296 22234
rect 34244 22170 34296 22176
rect 33968 22092 34020 22098
rect 33968 22034 34020 22040
rect 34624 21962 34652 22646
rect 34808 22545 34836 22918
rect 34992 22778 35020 23054
rect 35452 22778 35480 23462
rect 35544 22930 35572 24686
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35636 23798 35664 24006
rect 35624 23792 35676 23798
rect 35624 23734 35676 23740
rect 35716 23180 35768 23186
rect 35716 23122 35768 23128
rect 35728 23066 35756 23122
rect 35636 23050 35756 23066
rect 35624 23044 35756 23050
rect 35676 23038 35756 23044
rect 35624 22986 35676 22992
rect 35544 22902 35664 22930
rect 34980 22772 35032 22778
rect 34980 22714 35032 22720
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 34794 22536 34850 22545
rect 34794 22471 34850 22480
rect 34612 21956 34664 21962
rect 34612 21898 34664 21904
rect 34426 21720 34482 21729
rect 34426 21655 34482 21664
rect 34244 21412 34296 21418
rect 34244 21354 34296 21360
rect 34060 21072 34112 21078
rect 34060 21014 34112 21020
rect 33968 21004 34020 21010
rect 33968 20946 34020 20952
rect 33784 19848 33836 19854
rect 33784 19790 33836 19796
rect 33782 19544 33838 19553
rect 33782 19479 33838 19488
rect 33796 19446 33824 19479
rect 33784 19440 33836 19446
rect 33784 19382 33836 19388
rect 33876 19372 33928 19378
rect 33876 19314 33928 19320
rect 33692 19168 33744 19174
rect 33692 19110 33744 19116
rect 33784 19168 33836 19174
rect 33784 19110 33836 19116
rect 33598 19000 33654 19009
rect 33598 18935 33654 18944
rect 33692 18896 33744 18902
rect 33428 18856 33692 18884
rect 33428 18154 33456 18856
rect 33692 18838 33744 18844
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 33416 18148 33468 18154
rect 33416 18090 33468 18096
rect 33416 17876 33468 17882
rect 33416 17818 33468 17824
rect 33324 17740 33376 17746
rect 33324 17682 33376 17688
rect 33428 17542 33456 17818
rect 33416 17536 33468 17542
rect 33416 17478 33468 17484
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 33060 14958 33088 15302
rect 33048 14952 33100 14958
rect 33048 14894 33100 14900
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32864 14408 32916 14414
rect 32864 14350 32916 14356
rect 33336 14346 33364 16050
rect 33428 15978 33456 17478
rect 33416 15972 33468 15978
rect 33416 15914 33468 15920
rect 33416 14952 33468 14958
rect 33416 14894 33468 14900
rect 33324 14340 33376 14346
rect 33324 14282 33376 14288
rect 33428 14278 33456 14894
rect 32588 14272 32640 14278
rect 32588 14214 32640 14220
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 32600 13870 32628 14214
rect 32496 13864 32548 13870
rect 32496 13806 32548 13812
rect 32588 13864 32640 13870
rect 32588 13806 32640 13812
rect 32784 13376 32812 14214
rect 33416 13864 33468 13870
rect 33416 13806 33468 13812
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32692 13348 32812 13376
rect 32588 12640 32640 12646
rect 32588 12582 32640 12588
rect 32404 11892 32456 11898
rect 32404 11834 32456 11840
rect 32600 11778 32628 12582
rect 32692 11898 32720 13348
rect 33428 13190 33456 13806
rect 33416 13184 33468 13190
rect 33416 13126 33468 13132
rect 33428 12918 33456 13126
rect 32772 12912 32824 12918
rect 32772 12854 32824 12860
rect 33416 12912 33468 12918
rect 33416 12854 33468 12860
rect 32680 11892 32732 11898
rect 32680 11834 32732 11840
rect 32324 11750 32628 11778
rect 32324 10606 32352 11750
rect 32220 10600 32272 10606
rect 32220 10542 32272 10548
rect 32312 10600 32364 10606
rect 32312 10542 32364 10548
rect 32232 10470 32260 10542
rect 32220 10464 32272 10470
rect 32220 10406 32272 10412
rect 32784 10130 32812 12854
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 32864 12640 32916 12646
rect 32864 12582 32916 12588
rect 32876 12170 32904 12582
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32864 12164 32916 12170
rect 32864 12106 32916 12112
rect 32864 11688 32916 11694
rect 32864 11630 32916 11636
rect 32876 11286 32904 11630
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 33336 11354 33364 12786
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 32864 11280 32916 11286
rect 32864 11222 32916 11228
rect 32128 10124 32180 10130
rect 32128 10066 32180 10072
rect 32220 10124 32272 10130
rect 32220 10066 32272 10072
rect 32772 10124 32824 10130
rect 32772 10066 32824 10072
rect 32036 9920 32088 9926
rect 32036 9862 32088 9868
rect 32036 9716 32088 9722
rect 32036 9658 32088 9664
rect 31760 9512 31812 9518
rect 31588 9460 31760 9466
rect 31588 9454 31812 9460
rect 31944 9512 31996 9518
rect 31944 9454 31996 9460
rect 31588 9438 31800 9454
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31772 9194 31800 9318
rect 31680 9166 31800 9194
rect 30930 9007 30986 9016
rect 31484 9036 31536 9042
rect 30944 8974 30972 9007
rect 31484 8978 31536 8984
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 31128 7546 31156 8434
rect 31680 7818 31708 9166
rect 31772 8906 31800 9166
rect 31760 8900 31812 8906
rect 31760 8842 31812 8848
rect 31852 8424 31904 8430
rect 31852 8366 31904 8372
rect 31668 7812 31720 7818
rect 31668 7754 31720 7760
rect 31760 7812 31812 7818
rect 31760 7754 31812 7760
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31404 7546 31432 7686
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 30840 6384 30892 6390
rect 30840 6326 30892 6332
rect 31772 3534 31800 7754
rect 31864 7478 31892 8366
rect 31956 8362 31984 9454
rect 31944 8356 31996 8362
rect 31944 8298 31996 8304
rect 32048 8294 32076 9658
rect 32232 9450 32260 10066
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32404 9920 32456 9926
rect 32404 9862 32456 9868
rect 32310 9752 32366 9761
rect 32310 9687 32312 9696
rect 32364 9687 32366 9696
rect 32312 9658 32364 9664
rect 32220 9444 32272 9450
rect 32220 9386 32272 9392
rect 32416 9178 32444 9862
rect 32508 9654 32536 9998
rect 32680 9988 32732 9994
rect 32680 9930 32732 9936
rect 32496 9648 32548 9654
rect 32496 9590 32548 9596
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32508 9042 32536 9590
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32600 9178 32628 9318
rect 32588 9172 32640 9178
rect 32588 9114 32640 9120
rect 32496 9036 32548 9042
rect 32496 8978 32548 8984
rect 32508 8922 32536 8978
rect 32324 8894 32536 8922
rect 32128 8832 32180 8838
rect 32128 8774 32180 8780
rect 32140 8634 32168 8774
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 32324 8498 32352 8894
rect 32600 8650 32628 9114
rect 32508 8634 32628 8650
rect 32496 8628 32628 8634
rect 32548 8622 32628 8628
rect 32496 8570 32548 8576
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32036 8288 32088 8294
rect 32036 8230 32088 8236
rect 32232 7954 32260 8366
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32600 7750 32628 8502
rect 32692 7886 32720 9930
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32784 9042 32812 9454
rect 32876 9058 32904 11222
rect 33336 11150 33364 11290
rect 33324 11144 33376 11150
rect 33324 11086 33376 11092
rect 33324 10736 33376 10742
rect 33324 10678 33376 10684
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33336 9674 33364 10678
rect 33520 10062 33548 18702
rect 33796 18630 33824 19110
rect 33888 18766 33916 19314
rect 33876 18760 33928 18766
rect 33876 18702 33928 18708
rect 33784 18624 33836 18630
rect 33876 18624 33928 18630
rect 33784 18566 33836 18572
rect 33874 18592 33876 18601
rect 33928 18592 33930 18601
rect 33874 18527 33930 18536
rect 33980 18358 34008 20946
rect 33968 18352 34020 18358
rect 33968 18294 34020 18300
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33612 17338 33640 18158
rect 33888 17649 33916 18158
rect 33874 17640 33930 17649
rect 33874 17575 33930 17584
rect 33692 17536 33744 17542
rect 33692 17478 33744 17484
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 33704 16289 33732 17478
rect 33876 17060 33928 17066
rect 33876 17002 33928 17008
rect 33888 16794 33916 17002
rect 33876 16788 33928 16794
rect 33876 16730 33928 16736
rect 33968 16448 34020 16454
rect 33968 16390 34020 16396
rect 33690 16280 33746 16289
rect 33690 16215 33746 16224
rect 33692 15904 33744 15910
rect 33692 15846 33744 15852
rect 33600 14612 33652 14618
rect 33600 14554 33652 14560
rect 33612 11744 33640 14554
rect 33704 14414 33732 15846
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33888 15162 33916 15302
rect 33876 15156 33928 15162
rect 33876 15098 33928 15104
rect 33784 14952 33836 14958
rect 33784 14894 33836 14900
rect 33796 14550 33824 14894
rect 33980 14890 34008 16390
rect 34072 15094 34100 21014
rect 34256 21010 34284 21354
rect 34244 21004 34296 21010
rect 34244 20946 34296 20952
rect 34244 19780 34296 19786
rect 34244 19722 34296 19728
rect 34256 19514 34284 19722
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 34244 19508 34296 19514
rect 34244 19450 34296 19456
rect 34150 18864 34206 18873
rect 34150 18799 34152 18808
rect 34204 18799 34206 18808
rect 34152 18770 34204 18776
rect 34348 16454 34376 19654
rect 34440 19310 34468 21655
rect 34624 20942 34652 21898
rect 34808 21690 34836 22471
rect 35346 22400 35402 22409
rect 35346 22335 35402 22344
rect 35164 21888 35216 21894
rect 35084 21848 35164 21876
rect 35084 21690 35112 21848
rect 35256 21888 35308 21894
rect 35164 21830 35216 21836
rect 35254 21856 35256 21865
rect 35308 21856 35310 21865
rect 35254 21791 35310 21800
rect 34796 21684 34848 21690
rect 34796 21626 34848 21632
rect 35072 21684 35124 21690
rect 35072 21626 35124 21632
rect 34980 21344 35032 21350
rect 34980 21286 35032 21292
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34610 20496 34666 20505
rect 34610 20431 34666 20440
rect 34888 20460 34940 20466
rect 34520 20392 34572 20398
rect 34520 20334 34572 20340
rect 34428 19304 34480 19310
rect 34428 19246 34480 19252
rect 34532 18834 34560 20334
rect 34624 19446 34652 20431
rect 34888 20402 34940 20408
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34704 19984 34756 19990
rect 34704 19926 34756 19932
rect 34612 19440 34664 19446
rect 34612 19382 34664 19388
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 34624 18766 34652 19382
rect 34612 18760 34664 18766
rect 34612 18702 34664 18708
rect 34428 17536 34480 17542
rect 34428 17478 34480 17484
rect 34440 17270 34468 17478
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 34440 16794 34468 17206
rect 34428 16788 34480 16794
rect 34428 16730 34480 16736
rect 34440 16590 34468 16730
rect 34428 16584 34480 16590
rect 34428 16526 34480 16532
rect 34336 16448 34388 16454
rect 34336 16390 34388 16396
rect 34152 15904 34204 15910
rect 34152 15846 34204 15852
rect 34060 15088 34112 15094
rect 34060 15030 34112 15036
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 33784 14544 33836 14550
rect 33784 14486 33836 14492
rect 33692 14408 33744 14414
rect 33692 14350 33744 14356
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 33784 13524 33836 13530
rect 33784 13466 33836 13472
rect 33692 13388 33744 13394
rect 33692 13330 33744 13336
rect 33704 12782 33732 13330
rect 33692 12776 33744 12782
rect 33692 12718 33744 12724
rect 33796 11898 33824 13466
rect 34072 13326 34100 13806
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 33968 13252 34020 13258
rect 33968 13194 34020 13200
rect 33980 12832 34008 13194
rect 34072 12986 34100 13262
rect 34164 13190 34192 15846
rect 34348 15502 34376 16390
rect 34440 15706 34468 16526
rect 34428 15700 34480 15706
rect 34428 15642 34480 15648
rect 34336 15496 34388 15502
rect 34336 15438 34388 15444
rect 34612 14884 34664 14890
rect 34612 14826 34664 14832
rect 34244 14816 34296 14822
rect 34244 14758 34296 14764
rect 34256 14618 34284 14758
rect 34244 14612 34296 14618
rect 34244 14554 34296 14560
rect 34244 14272 34296 14278
rect 34244 14214 34296 14220
rect 34152 13184 34204 13190
rect 34152 13126 34204 13132
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 33888 12804 34008 12832
rect 33888 12306 33916 12804
rect 33876 12300 33928 12306
rect 33876 12242 33928 12248
rect 34164 12238 34192 13126
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 33784 11892 33836 11898
rect 33784 11834 33836 11840
rect 33692 11756 33744 11762
rect 33612 11716 33692 11744
rect 33692 11698 33744 11704
rect 33968 11688 34020 11694
rect 33968 11630 34020 11636
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33244 9646 33364 9674
rect 33244 9382 33272 9646
rect 33520 9489 33548 9998
rect 33506 9480 33562 9489
rect 33506 9415 33562 9424
rect 33232 9376 33284 9382
rect 33232 9318 33284 9324
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 33324 9104 33376 9110
rect 32772 9036 32824 9042
rect 32876 9030 32996 9058
rect 33324 9046 33376 9052
rect 32772 8978 32824 8984
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 31852 7472 31904 7478
rect 31852 7414 31904 7420
rect 32600 7206 32628 7686
rect 32784 7478 32812 8978
rect 32968 8430 32996 9030
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 33060 8430 33088 8978
rect 33336 8634 33364 9046
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33324 8628 33376 8634
rect 33324 8570 33376 8576
rect 33888 8566 33916 8910
rect 33876 8560 33928 8566
rect 33876 8502 33928 8508
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32772 7472 32824 7478
rect 32772 7414 32824 7420
rect 32588 7200 32640 7206
rect 32588 7142 32640 7148
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 33980 3602 34008 11630
rect 33968 3596 34020 3602
rect 33968 3538 34020 3544
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 29000 3460 29052 3466
rect 29000 3402 29052 3408
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 26332 2984 26384 2990
rect 26332 2926 26384 2932
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 26344 2650 26372 2926
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 24860 2576 24912 2582
rect 24860 2518 24912 2524
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 26528 800 26556 2450
rect 27172 2446 27200 2790
rect 29012 2650 29040 3402
rect 29552 3392 29604 3398
rect 29552 3334 29604 3340
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 29564 2514 29592 3334
rect 31312 3194 31340 3402
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31772 3126 31800 3470
rect 31760 3120 31812 3126
rect 31760 3062 31812 3068
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 31404 2650 31432 2994
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33704 2650 33732 2994
rect 31392 2644 31444 2650
rect 31392 2586 31444 2592
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 34164 2582 34192 12174
rect 34256 11694 34284 14214
rect 34428 13456 34480 13462
rect 34428 13398 34480 13404
rect 34440 12918 34468 13398
rect 34428 12912 34480 12918
rect 34428 12854 34480 12860
rect 34336 12096 34388 12102
rect 34336 12038 34388 12044
rect 34348 11898 34376 12038
rect 34336 11892 34388 11898
rect 34336 11834 34388 11840
rect 34440 11744 34468 12854
rect 34624 12850 34652 14826
rect 34716 14006 34744 19926
rect 34808 19378 34836 20334
rect 34900 19514 34928 20402
rect 34888 19508 34940 19514
rect 34888 19450 34940 19456
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 34808 19145 34836 19314
rect 34794 19136 34850 19145
rect 34794 19071 34850 19080
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34808 16250 34836 17070
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 34808 15570 34836 16186
rect 34900 15609 34928 19450
rect 34992 19446 35020 21286
rect 35084 21078 35112 21626
rect 35164 21344 35216 21350
rect 35164 21286 35216 21292
rect 35072 21072 35124 21078
rect 35072 21014 35124 21020
rect 35072 20392 35124 20398
rect 35072 20334 35124 20340
rect 35084 19922 35112 20334
rect 35072 19916 35124 19922
rect 35072 19858 35124 19864
rect 34980 19440 35032 19446
rect 34980 19382 35032 19388
rect 34980 18964 35032 18970
rect 34980 18906 35032 18912
rect 34886 15600 34942 15609
rect 34796 15564 34848 15570
rect 34886 15535 34942 15544
rect 34796 15506 34848 15512
rect 34808 14482 34836 15506
rect 34888 15428 34940 15434
rect 34888 15370 34940 15376
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 34796 14340 34848 14346
rect 34796 14282 34848 14288
rect 34704 14000 34756 14006
rect 34704 13942 34756 13948
rect 34704 13796 34756 13802
rect 34704 13738 34756 13744
rect 34612 12844 34664 12850
rect 34612 12786 34664 12792
rect 34520 12708 34572 12714
rect 34520 12650 34572 12656
rect 34348 11716 34468 11744
rect 34244 11688 34296 11694
rect 34244 11630 34296 11636
rect 34244 11552 34296 11558
rect 34244 11494 34296 11500
rect 34256 11286 34284 11494
rect 34244 11280 34296 11286
rect 34244 11222 34296 11228
rect 34244 9988 34296 9994
rect 34244 9930 34296 9936
rect 34256 9042 34284 9930
rect 34244 9036 34296 9042
rect 34244 8978 34296 8984
rect 34256 8838 34284 8978
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34348 8566 34376 11716
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 34440 11354 34468 11494
rect 34428 11348 34480 11354
rect 34428 11290 34480 11296
rect 34428 10192 34480 10198
rect 34428 10134 34480 10140
rect 34336 8560 34388 8566
rect 34336 8502 34388 8508
rect 34440 7478 34468 10134
rect 34532 8974 34560 12650
rect 34612 12164 34664 12170
rect 34612 12106 34664 12112
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34624 7954 34652 12106
rect 34716 10606 34744 13738
rect 34808 11082 34836 14282
rect 34900 14006 34928 15370
rect 34888 14000 34940 14006
rect 34888 13942 34940 13948
rect 34888 13320 34940 13326
rect 34888 13262 34940 13268
rect 34900 12918 34928 13262
rect 34992 12986 35020 18906
rect 35084 17814 35112 19858
rect 35072 17808 35124 17814
rect 35072 17750 35124 17756
rect 35072 17536 35124 17542
rect 35072 17478 35124 17484
rect 35084 17338 35112 17478
rect 35072 17332 35124 17338
rect 35072 17274 35124 17280
rect 35176 17202 35204 21286
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 35268 20777 35296 20878
rect 35254 20768 35310 20777
rect 35254 20703 35310 20712
rect 35268 20262 35296 20703
rect 35256 20256 35308 20262
rect 35256 20198 35308 20204
rect 35268 18290 35296 20198
rect 35360 19922 35388 22335
rect 35452 22166 35480 22714
rect 35532 22636 35584 22642
rect 35532 22578 35584 22584
rect 35440 22160 35492 22166
rect 35440 22102 35492 22108
rect 35348 19916 35400 19922
rect 35348 19858 35400 19864
rect 35544 18766 35572 22578
rect 35636 21622 35664 22902
rect 35820 22681 35848 26302
rect 36358 26200 36414 27000
rect 37002 26330 37058 27000
rect 37002 26302 37228 26330
rect 37002 26200 37058 26302
rect 35900 24404 35952 24410
rect 35900 24346 35952 24352
rect 35912 23594 35940 24346
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 35900 23588 35952 23594
rect 35900 23530 35952 23536
rect 36096 23497 36124 24006
rect 36176 23656 36228 23662
rect 36176 23598 36228 23604
rect 36082 23488 36138 23497
rect 36082 23423 36138 23432
rect 35898 23080 35954 23089
rect 35898 23015 35954 23024
rect 35992 23044 36044 23050
rect 35912 22778 35940 23015
rect 35992 22986 36044 22992
rect 36004 22953 36032 22986
rect 35990 22944 36046 22953
rect 35990 22879 36046 22888
rect 35900 22772 35952 22778
rect 35900 22714 35952 22720
rect 35806 22672 35862 22681
rect 35806 22607 35862 22616
rect 35808 22432 35860 22438
rect 35808 22374 35860 22380
rect 35624 21616 35676 21622
rect 35624 21558 35676 21564
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35728 21146 35756 21286
rect 35716 21140 35768 21146
rect 35716 21082 35768 21088
rect 35820 21026 35848 22374
rect 35912 22098 35940 22714
rect 36082 22128 36138 22137
rect 35900 22092 35952 22098
rect 36082 22063 36138 22072
rect 35900 22034 35952 22040
rect 35992 21480 36044 21486
rect 35992 21422 36044 21428
rect 36004 21350 36032 21422
rect 35992 21344 36044 21350
rect 35992 21286 36044 21292
rect 35728 20998 35848 21026
rect 35900 21004 35952 21010
rect 35728 19854 35756 20998
rect 35900 20946 35952 20952
rect 35912 20534 35940 20946
rect 35900 20528 35952 20534
rect 35900 20470 35952 20476
rect 36096 20262 36124 22063
rect 36188 21894 36216 23598
rect 36372 22710 36400 26200
rect 36452 24336 36504 24342
rect 36452 24278 36504 24284
rect 36464 23662 36492 24278
rect 36728 24268 36780 24274
rect 36728 24210 36780 24216
rect 36452 23656 36504 23662
rect 36452 23598 36504 23604
rect 36544 23656 36596 23662
rect 36544 23598 36596 23604
rect 36556 23526 36584 23598
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36636 23316 36688 23322
rect 36636 23258 36688 23264
rect 36360 22704 36412 22710
rect 36360 22646 36412 22652
rect 36452 22500 36504 22506
rect 36452 22442 36504 22448
rect 36176 21888 36228 21894
rect 36176 21830 36228 21836
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36268 21480 36320 21486
rect 36268 21422 36320 21428
rect 36188 20602 36216 21422
rect 36280 20806 36308 21422
rect 36268 20800 36320 20806
rect 36268 20742 36320 20748
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36084 20256 36136 20262
rect 36084 20198 36136 20204
rect 36176 19916 36228 19922
rect 36176 19858 36228 19864
rect 35716 19848 35768 19854
rect 35716 19790 35768 19796
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 36084 19712 36136 19718
rect 36084 19654 36136 19660
rect 35532 18760 35584 18766
rect 35532 18702 35584 18708
rect 35348 18692 35400 18698
rect 35348 18634 35400 18640
rect 35360 18426 35388 18634
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35256 18284 35308 18290
rect 35256 18226 35308 18232
rect 35532 17876 35584 17882
rect 35532 17818 35584 17824
rect 35256 17808 35308 17814
rect 35256 17750 35308 17756
rect 35164 17196 35216 17202
rect 35164 17138 35216 17144
rect 35164 15904 35216 15910
rect 35164 15846 35216 15852
rect 35176 14346 35204 15846
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 35176 14006 35204 14282
rect 35268 14056 35296 17750
rect 35544 17649 35572 17818
rect 35530 17640 35586 17649
rect 35530 17575 35586 17584
rect 35714 17640 35770 17649
rect 35714 17575 35770 17584
rect 35544 17542 35572 17575
rect 35440 17536 35492 17542
rect 35438 17504 35440 17513
rect 35532 17536 35584 17542
rect 35492 17504 35494 17513
rect 35532 17478 35584 17484
rect 35438 17439 35494 17448
rect 35452 17270 35480 17439
rect 35440 17264 35492 17270
rect 35440 17206 35492 17212
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 35360 14890 35388 16934
rect 35452 16590 35480 17206
rect 35440 16584 35492 16590
rect 35440 16526 35492 16532
rect 35532 16448 35584 16454
rect 35532 16390 35584 16396
rect 35348 14884 35400 14890
rect 35348 14826 35400 14832
rect 35440 14816 35492 14822
rect 35440 14758 35492 14764
rect 35452 14278 35480 14758
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35268 14028 35388 14056
rect 35164 14000 35216 14006
rect 35164 13942 35216 13948
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 35164 13184 35216 13190
rect 35164 13126 35216 13132
rect 34980 12980 35032 12986
rect 34980 12922 35032 12928
rect 34888 12912 34940 12918
rect 35176 12889 35204 13126
rect 34888 12854 34940 12860
rect 35162 12880 35218 12889
rect 34900 12238 34928 12854
rect 35162 12815 35218 12824
rect 35164 12776 35216 12782
rect 35164 12718 35216 12724
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 34900 11694 34928 12174
rect 35176 12170 35204 12718
rect 35164 12164 35216 12170
rect 35164 12106 35216 12112
rect 35268 11898 35296 13874
rect 35360 12782 35388 14028
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 35256 11892 35308 11898
rect 35256 11834 35308 11840
rect 35072 11824 35124 11830
rect 35072 11766 35124 11772
rect 34888 11688 34940 11694
rect 34888 11630 34940 11636
rect 34796 11076 34848 11082
rect 34796 11018 34848 11024
rect 34704 10600 34756 10606
rect 34704 10542 34756 10548
rect 34716 10130 34744 10542
rect 34704 10124 34756 10130
rect 34704 10066 34756 10072
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 34900 9722 34928 9998
rect 34888 9716 34940 9722
rect 34888 9658 34940 9664
rect 35084 9042 35112 11766
rect 35544 11082 35572 16390
rect 35728 16153 35756 17575
rect 35714 16144 35770 16153
rect 35714 16079 35770 16088
rect 35714 16008 35770 16017
rect 35714 15943 35770 15952
rect 35728 14521 35756 15943
rect 35820 15094 35848 19654
rect 35900 19372 35952 19378
rect 35900 19314 35952 19320
rect 35912 18086 35940 19314
rect 35992 19304 36044 19310
rect 35992 19246 36044 19252
rect 35900 18080 35952 18086
rect 35900 18022 35952 18028
rect 36004 17184 36032 19246
rect 36096 19009 36124 19654
rect 36082 19000 36138 19009
rect 36082 18935 36138 18944
rect 36084 18624 36136 18630
rect 36084 18566 36136 18572
rect 36096 18358 36124 18566
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 36096 17660 36124 18294
rect 36188 17882 36216 19858
rect 36372 19786 36400 21830
rect 36360 19780 36412 19786
rect 36360 19722 36412 19728
rect 36464 19174 36492 22442
rect 36544 21956 36596 21962
rect 36544 21898 36596 21904
rect 36556 21418 36584 21898
rect 36648 21418 36676 23258
rect 36544 21412 36596 21418
rect 36544 21354 36596 21360
rect 36636 21412 36688 21418
rect 36636 21354 36688 21360
rect 36740 21146 36768 24210
rect 36820 24064 36872 24070
rect 36820 24006 36872 24012
rect 36832 22166 36860 24006
rect 37004 23044 37056 23050
rect 37004 22986 37056 22992
rect 36912 22976 36964 22982
rect 37016 22953 37044 22986
rect 36912 22918 36964 22924
rect 37002 22944 37058 22953
rect 36924 22438 36952 22918
rect 37002 22879 37058 22888
rect 36912 22432 36964 22438
rect 36912 22374 36964 22380
rect 36820 22160 36872 22166
rect 36820 22102 36872 22108
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36924 21010 36952 22374
rect 37200 22114 37228 26302
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 37752 26302 38346 26330
rect 37556 24404 37608 24410
rect 37556 24346 37608 24352
rect 37464 24268 37516 24274
rect 37464 24210 37516 24216
rect 37370 23488 37426 23497
rect 37370 23423 37426 23432
rect 37384 23118 37412 23423
rect 37372 23112 37424 23118
rect 37372 23054 37424 23060
rect 37280 22704 37332 22710
rect 37280 22646 37332 22652
rect 37292 22545 37320 22646
rect 37278 22536 37334 22545
rect 37278 22471 37334 22480
rect 37278 22128 37334 22137
rect 37096 22092 37148 22098
rect 37200 22086 37278 22114
rect 37278 22063 37334 22072
rect 37096 22034 37148 22040
rect 37004 21344 37056 21350
rect 37004 21286 37056 21292
rect 36912 21004 36964 21010
rect 36912 20946 36964 20952
rect 36912 20800 36964 20806
rect 36912 20742 36964 20748
rect 36924 20602 36952 20742
rect 36912 20596 36964 20602
rect 36912 20538 36964 20544
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36556 19514 36584 19654
rect 36924 19514 36952 20538
rect 36544 19508 36596 19514
rect 36544 19450 36596 19456
rect 36912 19508 36964 19514
rect 36912 19450 36964 19456
rect 36452 19168 36504 19174
rect 36452 19110 36504 19116
rect 36636 19168 36688 19174
rect 36912 19168 36964 19174
rect 36636 19110 36688 19116
rect 36910 19136 36912 19145
rect 36964 19136 36966 19145
rect 36268 18284 36320 18290
rect 36268 18226 36320 18232
rect 36176 17876 36228 17882
rect 36176 17818 36228 17824
rect 36176 17672 36228 17678
rect 36096 17632 36176 17660
rect 36176 17614 36228 17620
rect 35912 17156 36032 17184
rect 35912 16522 35940 17156
rect 36188 16794 36216 17614
rect 36176 16788 36228 16794
rect 36176 16730 36228 16736
rect 35900 16516 35952 16522
rect 35900 16458 35952 16464
rect 35912 15570 35940 16458
rect 36188 16182 36216 16730
rect 36176 16176 36228 16182
rect 36176 16118 36228 16124
rect 36188 15570 36216 16118
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 36176 15564 36228 15570
rect 36176 15506 36228 15512
rect 35900 15360 35952 15366
rect 35900 15302 35952 15308
rect 35808 15088 35860 15094
rect 35808 15030 35860 15036
rect 35714 14512 35770 14521
rect 35714 14447 35770 14456
rect 35624 13932 35676 13938
rect 35624 13874 35676 13880
rect 35636 11665 35664 13874
rect 35912 13258 35940 15302
rect 35992 14816 36044 14822
rect 35992 14758 36044 14764
rect 35900 13252 35952 13258
rect 35900 13194 35952 13200
rect 35716 13184 35768 13190
rect 35716 13126 35768 13132
rect 35728 11830 35756 13126
rect 35808 12776 35860 12782
rect 35808 12718 35860 12724
rect 35820 12646 35848 12718
rect 35808 12640 35860 12646
rect 35808 12582 35860 12588
rect 35716 11824 35768 11830
rect 35716 11766 35768 11772
rect 35622 11656 35678 11665
rect 35622 11591 35678 11600
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35532 11076 35584 11082
rect 35532 11018 35584 11024
rect 35636 10674 35664 11494
rect 35728 11218 35756 11766
rect 35716 11212 35768 11218
rect 35716 11154 35768 11160
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35624 10532 35676 10538
rect 35624 10474 35676 10480
rect 35636 10248 35664 10474
rect 35452 10220 35664 10248
rect 35164 10124 35216 10130
rect 35164 10066 35216 10072
rect 35176 9722 35204 10066
rect 35452 9994 35480 10220
rect 35728 9994 35756 11154
rect 35900 11076 35952 11082
rect 35900 11018 35952 11024
rect 35440 9988 35492 9994
rect 35440 9930 35492 9936
rect 35716 9988 35768 9994
rect 35716 9930 35768 9936
rect 35728 9722 35756 9930
rect 35164 9716 35216 9722
rect 35164 9658 35216 9664
rect 35716 9716 35768 9722
rect 35716 9658 35768 9664
rect 35912 9518 35940 11018
rect 35900 9512 35952 9518
rect 35900 9454 35952 9460
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35544 9042 35572 9318
rect 36004 9110 36032 14758
rect 36176 13932 36228 13938
rect 36176 13874 36228 13880
rect 36188 13734 36216 13874
rect 36176 13728 36228 13734
rect 36176 13670 36228 13676
rect 36280 13530 36308 18226
rect 36648 17542 36676 19110
rect 36910 19071 36966 19080
rect 36820 18624 36872 18630
rect 36820 18566 36872 18572
rect 36728 18080 36780 18086
rect 36728 18022 36780 18028
rect 36636 17536 36688 17542
rect 36636 17478 36688 17484
rect 36360 17196 36412 17202
rect 36360 17138 36412 17144
rect 36372 16794 36400 17138
rect 36544 17128 36596 17134
rect 36544 17070 36596 17076
rect 36360 16788 36412 16794
rect 36360 16730 36412 16736
rect 36358 16280 36414 16289
rect 36358 16215 36414 16224
rect 36372 15094 36400 16215
rect 36452 15564 36504 15570
rect 36452 15506 36504 15512
rect 36360 15088 36412 15094
rect 36360 15030 36412 15036
rect 36464 14346 36492 15506
rect 36556 15042 36584 17070
rect 36636 16992 36688 16998
rect 36636 16934 36688 16940
rect 36648 16794 36676 16934
rect 36636 16788 36688 16794
rect 36636 16730 36688 16736
rect 36634 16688 36690 16697
rect 36634 16623 36690 16632
rect 36648 16590 36676 16623
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 36740 16454 36768 18022
rect 36728 16448 36780 16454
rect 36728 16390 36780 16396
rect 36556 15014 36676 15042
rect 36544 14884 36596 14890
rect 36544 14826 36596 14832
rect 36452 14340 36504 14346
rect 36452 14282 36504 14288
rect 36464 13802 36492 14282
rect 36452 13796 36504 13802
rect 36452 13738 36504 13744
rect 36268 13524 36320 13530
rect 36268 13466 36320 13472
rect 36450 12880 36506 12889
rect 36450 12815 36506 12824
rect 36464 12782 36492 12815
rect 36452 12776 36504 12782
rect 36452 12718 36504 12724
rect 36556 12102 36584 14826
rect 36648 14618 36676 15014
rect 36636 14612 36688 14618
rect 36636 14554 36688 14560
rect 36648 13870 36676 14554
rect 36636 13864 36688 13870
rect 36636 13806 36688 13812
rect 36648 13258 36676 13806
rect 36740 13546 36768 16390
rect 36832 14278 36860 18566
rect 36912 18284 36964 18290
rect 36912 18226 36964 18232
rect 36924 16266 36952 18226
rect 37016 18154 37044 21286
rect 37108 20602 37136 22034
rect 37372 21888 37424 21894
rect 37278 21856 37334 21865
rect 37476 21876 37504 24210
rect 37568 22506 37596 24346
rect 37660 22574 37688 26200
rect 37648 22568 37700 22574
rect 37648 22510 37700 22516
rect 37556 22500 37608 22506
rect 37556 22442 37608 22448
rect 37648 22092 37700 22098
rect 37648 22034 37700 22040
rect 37424 21848 37504 21876
rect 37372 21830 37424 21836
rect 37278 21791 37334 21800
rect 37292 21622 37320 21791
rect 37384 21729 37412 21830
rect 37370 21720 37426 21729
rect 37370 21655 37426 21664
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 37188 21480 37240 21486
rect 37186 21448 37188 21457
rect 37240 21448 37242 21457
rect 37186 21383 37242 21392
rect 37280 21344 37332 21350
rect 37280 21286 37332 21292
rect 37292 20806 37320 21286
rect 37384 21078 37412 21655
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37568 21185 37596 21490
rect 37660 21350 37688 22034
rect 37648 21344 37700 21350
rect 37648 21286 37700 21292
rect 37554 21176 37610 21185
rect 37752 21146 37780 26302
rect 38290 26200 38346 26302
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43352 26376 43404 26382
rect 43352 26318 43404 26324
rect 38844 24676 38896 24682
rect 38844 24618 38896 24624
rect 38660 24336 38712 24342
rect 38712 24296 38792 24324
rect 38660 24278 38712 24284
rect 37832 24064 37884 24070
rect 37832 24006 37884 24012
rect 38384 24064 38436 24070
rect 38384 24006 38436 24012
rect 37844 23769 37872 24006
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 37830 23760 37886 23769
rect 37830 23695 37886 23704
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37832 22636 37884 22642
rect 37832 22578 37884 22584
rect 37844 22098 37872 22578
rect 37832 22092 37884 22098
rect 37832 22034 37884 22040
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37832 21616 37884 21622
rect 37832 21558 37884 21564
rect 37554 21111 37610 21120
rect 37648 21140 37700 21146
rect 37648 21082 37700 21088
rect 37740 21140 37792 21146
rect 37740 21082 37792 21088
rect 37372 21072 37424 21078
rect 37372 21014 37424 21020
rect 37556 20868 37608 20874
rect 37556 20810 37608 20816
rect 37280 20800 37332 20806
rect 37278 20768 37280 20777
rect 37332 20768 37334 20777
rect 37278 20703 37334 20712
rect 37096 20596 37148 20602
rect 37096 20538 37148 20544
rect 37188 20528 37240 20534
rect 37188 20470 37240 20476
rect 37094 19000 37150 19009
rect 37094 18935 37150 18944
rect 37108 18193 37136 18935
rect 37200 18426 37228 20470
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37280 20392 37332 20398
rect 37280 20334 37332 20340
rect 37292 18834 37320 20334
rect 37372 19916 37424 19922
rect 37372 19858 37424 19864
rect 37280 18828 37332 18834
rect 37280 18770 37332 18776
rect 37188 18420 37240 18426
rect 37188 18362 37240 18368
rect 37292 18358 37320 18770
rect 37280 18352 37332 18358
rect 37280 18294 37332 18300
rect 37094 18184 37150 18193
rect 37004 18148 37056 18154
rect 37094 18119 37150 18128
rect 37004 18090 37056 18096
rect 37016 16640 37044 18090
rect 37280 16992 37332 16998
rect 37280 16934 37332 16940
rect 37096 16652 37148 16658
rect 37016 16612 37096 16640
rect 37096 16594 37148 16600
rect 36924 16250 37044 16266
rect 36924 16244 37056 16250
rect 36924 16238 37004 16244
rect 37004 16186 37056 16192
rect 37108 16130 37136 16594
rect 37016 16102 37136 16130
rect 36820 14272 36872 14278
rect 36820 14214 36872 14220
rect 37016 14006 37044 16102
rect 37188 15904 37240 15910
rect 37188 15846 37240 15852
rect 37200 14521 37228 15846
rect 37186 14512 37242 14521
rect 37096 14476 37148 14482
rect 37186 14447 37242 14456
rect 37096 14418 37148 14424
rect 37004 14000 37056 14006
rect 37004 13942 37056 13948
rect 36740 13518 36952 13546
rect 36728 13388 36780 13394
rect 36728 13330 36780 13336
rect 36636 13252 36688 13258
rect 36636 13194 36688 13200
rect 36740 12986 36768 13330
rect 36728 12980 36780 12986
rect 36728 12922 36780 12928
rect 36924 12918 36952 13518
rect 36912 12912 36964 12918
rect 36912 12854 36964 12860
rect 36924 12646 36952 12854
rect 36912 12640 36964 12646
rect 36912 12582 36964 12588
rect 36924 12434 36952 12582
rect 36924 12406 37044 12434
rect 36544 12096 36596 12102
rect 36464 12056 36544 12084
rect 36464 11694 36492 12056
rect 36544 12038 36596 12044
rect 36728 12096 36780 12102
rect 36728 12038 36780 12044
rect 36740 11830 36768 12038
rect 36728 11824 36780 11830
rect 36728 11766 36780 11772
rect 36820 11756 36872 11762
rect 36820 11698 36872 11704
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 36648 10742 36676 11630
rect 36832 10810 36860 11698
rect 36820 10804 36872 10810
rect 36820 10746 36872 10752
rect 36636 10736 36688 10742
rect 36636 10678 36688 10684
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36084 9648 36136 9654
rect 36084 9590 36136 9596
rect 35992 9104 36044 9110
rect 35990 9072 35992 9081
rect 36044 9072 36046 9081
rect 34980 9036 35032 9042
rect 34980 8978 35032 8984
rect 35072 9036 35124 9042
rect 35072 8978 35124 8984
rect 35532 9036 35584 9042
rect 35990 9007 36046 9016
rect 35532 8978 35584 8984
rect 34992 8634 35020 8978
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 35624 8832 35676 8838
rect 35624 8774 35676 8780
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 35268 8090 35296 8774
rect 35636 8566 35664 8774
rect 35624 8560 35676 8566
rect 35624 8502 35676 8508
rect 36096 8498 36124 9590
rect 36372 9178 36400 10542
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 36464 8906 36492 10610
rect 36542 10568 36598 10577
rect 36542 10503 36544 10512
rect 36596 10503 36598 10512
rect 36544 10474 36596 10480
rect 36648 10266 36676 10678
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36636 10260 36688 10266
rect 36636 10202 36688 10208
rect 36924 9926 36952 10406
rect 36820 9920 36872 9926
rect 36820 9862 36872 9868
rect 36912 9920 36964 9926
rect 36912 9862 36964 9868
rect 36452 8900 36504 8906
rect 36452 8842 36504 8848
rect 36832 8498 36860 9862
rect 36924 9722 36952 9862
rect 36912 9716 36964 9722
rect 36912 9658 36964 9664
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 35256 8084 35308 8090
rect 35256 8026 35308 8032
rect 34612 7948 34664 7954
rect 34612 7890 34664 7896
rect 34428 7472 34480 7478
rect 34428 7414 34480 7420
rect 37016 6322 37044 12406
rect 37108 12238 37136 14418
rect 37188 14272 37240 14278
rect 37188 14214 37240 14220
rect 37200 13938 37228 14214
rect 37292 14006 37320 16934
rect 37384 16266 37412 19858
rect 37476 16998 37504 20402
rect 37568 19718 37596 20810
rect 37660 20398 37688 21082
rect 37740 20800 37792 20806
rect 37740 20742 37792 20748
rect 37752 20534 37780 20742
rect 37740 20528 37792 20534
rect 37740 20470 37792 20476
rect 37648 20392 37700 20398
rect 37648 20334 37700 20340
rect 37648 20256 37700 20262
rect 37648 20198 37700 20204
rect 37740 20256 37792 20262
rect 37740 20198 37792 20204
rect 37556 19712 37608 19718
rect 37556 19654 37608 19660
rect 37568 18630 37596 19654
rect 37660 19145 37688 20198
rect 37752 19242 37780 20198
rect 37844 19854 37872 21558
rect 37924 21480 37976 21486
rect 38292 21480 38344 21486
rect 37924 21422 37976 21428
rect 38212 21440 38292 21468
rect 37936 21010 37964 21422
rect 38108 21072 38160 21078
rect 38212 21060 38240 21440
rect 38292 21422 38344 21428
rect 38160 21032 38240 21060
rect 38108 21014 38160 21020
rect 37924 21004 37976 21010
rect 37924 20946 37976 20952
rect 38396 20913 38424 24006
rect 38568 23520 38620 23526
rect 38568 23462 38620 23468
rect 38580 23202 38608 23462
rect 38580 23186 38700 23202
rect 38580 23180 38712 23186
rect 38580 23174 38660 23180
rect 38660 23122 38712 23128
rect 38660 23044 38712 23050
rect 38660 22986 38712 22992
rect 38672 22778 38700 22986
rect 38660 22772 38712 22778
rect 38660 22714 38712 22720
rect 38566 21856 38622 21865
rect 38566 21791 38622 21800
rect 38580 21622 38608 21791
rect 38568 21616 38620 21622
rect 38568 21558 38620 21564
rect 38382 20904 38438 20913
rect 38382 20839 38438 20848
rect 38764 20806 38792 24296
rect 38856 24206 38884 24618
rect 38844 24200 38896 24206
rect 38844 24142 38896 24148
rect 38856 23730 38884 24142
rect 38844 23724 38896 23730
rect 38844 23666 38896 23672
rect 38948 22778 38976 26200
rect 39212 24744 39264 24750
rect 39212 24686 39264 24692
rect 39224 23798 39252 24686
rect 39592 24682 39620 26200
rect 39396 24676 39448 24682
rect 39396 24618 39448 24624
rect 39580 24676 39632 24682
rect 39580 24618 39632 24624
rect 39408 24410 39436 24618
rect 39488 24608 39540 24614
rect 39488 24550 39540 24556
rect 39396 24404 39448 24410
rect 39396 24346 39448 24352
rect 39500 24206 39528 24550
rect 40132 24268 40184 24274
rect 40132 24210 40184 24216
rect 39488 24200 39540 24206
rect 39488 24142 39540 24148
rect 39212 23792 39264 23798
rect 39212 23734 39264 23740
rect 39302 23760 39358 23769
rect 39302 23695 39358 23704
rect 39316 23322 39344 23695
rect 39500 23594 39528 24142
rect 40040 24064 40092 24070
rect 40040 24006 40092 24012
rect 40052 23866 40080 24006
rect 40040 23860 40092 23866
rect 40040 23802 40092 23808
rect 39764 23656 39816 23662
rect 39764 23598 39816 23604
rect 39946 23624 40002 23633
rect 39488 23588 39540 23594
rect 39488 23530 39540 23536
rect 39396 23520 39448 23526
rect 39396 23462 39448 23468
rect 39028 23316 39080 23322
rect 39028 23258 39080 23264
rect 39304 23316 39356 23322
rect 39304 23258 39356 23264
rect 38936 22772 38988 22778
rect 38936 22714 38988 22720
rect 38844 22704 38896 22710
rect 38844 22646 38896 22652
rect 38856 22574 38884 22646
rect 38844 22568 38896 22574
rect 38844 22510 38896 22516
rect 38844 21956 38896 21962
rect 38844 21898 38896 21904
rect 38856 21706 38884 21898
rect 39040 21706 39068 23258
rect 39212 23180 39264 23186
rect 39212 23122 39264 23128
rect 39224 22642 39252 23122
rect 39408 23089 39436 23462
rect 39394 23080 39450 23089
rect 39394 23015 39450 23024
rect 39776 22982 39804 23598
rect 39946 23559 40002 23568
rect 39960 22982 39988 23559
rect 39764 22976 39816 22982
rect 39764 22918 39816 22924
rect 39948 22976 40000 22982
rect 39948 22918 40000 22924
rect 39776 22642 39804 22918
rect 39212 22636 39264 22642
rect 39212 22578 39264 22584
rect 39764 22636 39816 22642
rect 39764 22578 39816 22584
rect 39224 22234 39252 22578
rect 39304 22500 39356 22506
rect 39304 22442 39356 22448
rect 39488 22500 39540 22506
rect 39488 22442 39540 22448
rect 39120 22228 39172 22234
rect 39120 22170 39172 22176
rect 39212 22228 39264 22234
rect 39212 22170 39264 22176
rect 38856 21678 39068 21706
rect 39132 20874 39160 22170
rect 39316 21894 39344 22442
rect 39500 22001 39528 22442
rect 39580 22228 39632 22234
rect 39580 22170 39632 22176
rect 39486 21992 39542 22001
rect 39486 21927 39542 21936
rect 39304 21888 39356 21894
rect 39304 21830 39356 21836
rect 39592 21570 39620 22170
rect 39776 22114 39804 22578
rect 40040 22432 40092 22438
rect 40040 22374 40092 22380
rect 39856 22160 39908 22166
rect 39776 22108 39856 22114
rect 39776 22102 39908 22108
rect 39776 22086 39896 22102
rect 39776 21622 39804 22086
rect 40052 21690 40080 22374
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 39500 21542 39620 21570
rect 39764 21616 39816 21622
rect 39764 21558 39816 21564
rect 39500 21418 39528 21542
rect 39580 21480 39632 21486
rect 39580 21422 39632 21428
rect 39764 21480 39816 21486
rect 39764 21422 39816 21428
rect 39488 21412 39540 21418
rect 39488 21354 39540 21360
rect 39500 21010 39528 21354
rect 39592 21146 39620 21422
rect 39580 21140 39632 21146
rect 39580 21082 39632 21088
rect 39776 21010 39804 21422
rect 40038 21312 40094 21321
rect 40038 21247 40094 21256
rect 39488 21004 39540 21010
rect 39488 20946 39540 20952
rect 39764 21004 39816 21010
rect 39764 20946 39816 20952
rect 39120 20868 39172 20874
rect 39120 20810 39172 20816
rect 38752 20800 38804 20806
rect 38474 20768 38530 20777
rect 38752 20742 38804 20748
rect 37950 20700 38258 20709
rect 38474 20703 38530 20712
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37924 20528 37976 20534
rect 37924 20470 37976 20476
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37936 19700 37964 20470
rect 38200 20052 38252 20058
rect 38200 19994 38252 20000
rect 38292 20052 38344 20058
rect 38292 19994 38344 20000
rect 38212 19854 38240 19994
rect 38200 19848 38252 19854
rect 38200 19790 38252 19796
rect 37844 19672 37964 19700
rect 37844 19310 37872 19672
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 38304 19378 38332 19994
rect 38384 19712 38436 19718
rect 38384 19654 38436 19660
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 37832 19304 37884 19310
rect 37832 19246 37884 19252
rect 37740 19236 37792 19242
rect 37740 19178 37792 19184
rect 37646 19136 37702 19145
rect 37646 19071 37702 19080
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37568 18154 37596 18566
rect 37752 18306 37780 19178
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 37660 18278 37780 18306
rect 37556 18148 37608 18154
rect 37556 18090 37608 18096
rect 37568 17678 37596 18090
rect 37660 17882 37688 18278
rect 37844 18222 37872 19110
rect 38014 18728 38070 18737
rect 38014 18663 38070 18672
rect 38028 18630 38056 18663
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 38396 18442 38424 19654
rect 38488 19514 38516 20703
rect 39500 20466 39528 20946
rect 39776 20874 39804 20946
rect 39764 20868 39816 20874
rect 39764 20810 39816 20816
rect 40052 20777 40080 21247
rect 40144 20874 40172 24210
rect 40236 21554 40264 26200
rect 40592 24812 40644 24818
rect 40592 24754 40644 24760
rect 40408 24608 40460 24614
rect 40408 24550 40460 24556
rect 40420 24206 40448 24550
rect 40604 24274 40632 24754
rect 42168 24274 42196 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 42892 24336 42944 24342
rect 42892 24278 42944 24284
rect 43364 24290 43392 26318
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26200 45430 27000
rect 46018 26330 46074 27000
rect 46018 26302 46336 26330
rect 46018 26200 46074 26302
rect 43904 24744 43956 24750
rect 43534 24712 43590 24721
rect 43904 24686 43956 24692
rect 43534 24647 43590 24656
rect 43548 24342 43576 24647
rect 43536 24336 43588 24342
rect 40592 24268 40644 24274
rect 40592 24210 40644 24216
rect 42156 24268 42208 24274
rect 42156 24210 42208 24216
rect 40408 24200 40460 24206
rect 40408 24142 40460 24148
rect 42156 24132 42208 24138
rect 42156 24074 42208 24080
rect 40960 24064 41012 24070
rect 40960 24006 41012 24012
rect 40682 23216 40738 23225
rect 40682 23151 40738 23160
rect 40500 22976 40552 22982
rect 40500 22918 40552 22924
rect 40408 22636 40460 22642
rect 40408 22578 40460 22584
rect 40316 22432 40368 22438
rect 40314 22400 40316 22409
rect 40368 22400 40370 22409
rect 40314 22335 40370 22344
rect 40316 22092 40368 22098
rect 40316 22034 40368 22040
rect 40224 21548 40276 21554
rect 40224 21490 40276 21496
rect 40328 21185 40356 22034
rect 40314 21176 40370 21185
rect 40314 21111 40370 21120
rect 40132 20868 40184 20874
rect 40132 20810 40184 20816
rect 40038 20768 40094 20777
rect 40038 20703 40094 20712
rect 39488 20460 39540 20466
rect 39488 20402 39540 20408
rect 39764 20460 39816 20466
rect 39764 20402 39816 20408
rect 39396 19916 39448 19922
rect 39396 19858 39448 19864
rect 38476 19508 38528 19514
rect 38476 19450 38528 19456
rect 39408 19310 39436 19858
rect 39776 19825 39804 20402
rect 40132 20392 40184 20398
rect 40132 20334 40184 20340
rect 39856 19848 39908 19854
rect 39762 19816 39818 19825
rect 39856 19790 39908 19796
rect 39762 19751 39818 19760
rect 39396 19304 39448 19310
rect 39396 19246 39448 19252
rect 39672 19304 39724 19310
rect 39672 19246 39724 19252
rect 39408 18970 39436 19246
rect 39396 18964 39448 18970
rect 39396 18906 39448 18912
rect 39684 18834 39712 19246
rect 39868 19242 39896 19790
rect 40040 19780 40092 19786
rect 40040 19722 40092 19728
rect 40052 19514 40080 19722
rect 40040 19508 40092 19514
rect 40040 19450 40092 19456
rect 39856 19236 39908 19242
rect 39856 19178 39908 19184
rect 38568 18828 38620 18834
rect 38568 18770 38620 18776
rect 39672 18828 39724 18834
rect 39672 18770 39724 18776
rect 38476 18624 38528 18630
rect 38476 18566 38528 18572
rect 38304 18414 38424 18442
rect 38016 18352 38068 18358
rect 38016 18294 38068 18300
rect 37740 18216 37792 18222
rect 37740 18158 37792 18164
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 37648 17876 37700 17882
rect 37648 17818 37700 17824
rect 37648 17740 37700 17746
rect 37648 17682 37700 17688
rect 37556 17672 37608 17678
rect 37556 17614 37608 17620
rect 37464 16992 37516 16998
rect 37464 16934 37516 16940
rect 37568 16726 37596 17614
rect 37556 16720 37608 16726
rect 37556 16662 37608 16668
rect 37384 16238 37596 16266
rect 37372 16108 37424 16114
rect 37372 16050 37424 16056
rect 37384 15570 37412 16050
rect 37464 16040 37516 16046
rect 37464 15982 37516 15988
rect 37372 15564 37424 15570
rect 37372 15506 37424 15512
rect 37384 15026 37412 15506
rect 37476 15162 37504 15982
rect 37464 15156 37516 15162
rect 37464 15098 37516 15104
rect 37372 15020 37424 15026
rect 37372 14962 37424 14968
rect 37384 14482 37412 14962
rect 37372 14476 37424 14482
rect 37372 14418 37424 14424
rect 37568 14278 37596 16238
rect 37660 15978 37688 17682
rect 37648 15972 37700 15978
rect 37648 15914 37700 15920
rect 37660 15706 37688 15914
rect 37752 15706 37780 18158
rect 37844 17134 37872 18158
rect 38028 18154 38056 18294
rect 38016 18148 38068 18154
rect 38016 18090 38068 18096
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 38304 16561 38332 18414
rect 38384 18284 38436 18290
rect 38384 18226 38436 18232
rect 38396 17626 38424 18226
rect 38488 17882 38516 18566
rect 38476 17876 38528 17882
rect 38476 17818 38528 17824
rect 38396 17598 38516 17626
rect 38384 17536 38436 17542
rect 38384 17478 38436 17484
rect 38290 16552 38346 16561
rect 38290 16487 38346 16496
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37648 15700 37700 15706
rect 37648 15642 37700 15648
rect 37740 15700 37792 15706
rect 37740 15642 37792 15648
rect 37752 15094 37780 15642
rect 37832 15360 37884 15366
rect 37832 15302 37884 15308
rect 37740 15088 37792 15094
rect 37740 15030 37792 15036
rect 37556 14272 37608 14278
rect 37556 14214 37608 14220
rect 37280 14000 37332 14006
rect 37280 13942 37332 13948
rect 37188 13932 37240 13938
rect 37188 13874 37240 13880
rect 37844 13530 37872 15302
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 38396 14618 38424 17478
rect 38488 17338 38516 17598
rect 38476 17332 38528 17338
rect 38476 17274 38528 17280
rect 38580 16454 38608 18770
rect 39684 18698 39712 18770
rect 39672 18692 39724 18698
rect 39672 18634 39724 18640
rect 39684 18442 39712 18634
rect 40144 18630 40172 20334
rect 40328 19922 40356 21111
rect 40420 21026 40448 22578
rect 40512 22234 40540 22918
rect 40696 22574 40724 23151
rect 40684 22568 40736 22574
rect 40684 22510 40736 22516
rect 40500 22228 40552 22234
rect 40500 22170 40552 22176
rect 40684 22092 40736 22098
rect 40684 22034 40736 22040
rect 40696 21962 40724 22034
rect 40684 21956 40736 21962
rect 40684 21898 40736 21904
rect 40592 21888 40644 21894
rect 40590 21856 40592 21865
rect 40644 21856 40646 21865
rect 40590 21791 40646 21800
rect 40972 21690 41000 24006
rect 41696 23860 41748 23866
rect 41696 23802 41748 23808
rect 41052 23656 41104 23662
rect 41052 23598 41104 23604
rect 41064 23186 41092 23598
rect 41512 23588 41564 23594
rect 41512 23530 41564 23536
rect 41052 23180 41104 23186
rect 41052 23122 41104 23128
rect 41064 22982 41092 23122
rect 41524 23118 41552 23530
rect 41604 23316 41656 23322
rect 41604 23258 41656 23264
rect 41512 23112 41564 23118
rect 41512 23054 41564 23060
rect 41236 23044 41288 23050
rect 41236 22986 41288 22992
rect 41052 22976 41104 22982
rect 41052 22918 41104 22924
rect 41144 22636 41196 22642
rect 41144 22578 41196 22584
rect 40960 21684 41012 21690
rect 40960 21626 41012 21632
rect 41052 21480 41104 21486
rect 41052 21422 41104 21428
rect 40868 21344 40920 21350
rect 41064 21332 41092 21422
rect 40920 21304 41092 21332
rect 40868 21286 40920 21292
rect 40868 21072 40920 21078
rect 40420 21020 40868 21026
rect 40420 21014 40920 21020
rect 40420 20998 40908 21014
rect 40316 19916 40368 19922
rect 40316 19858 40368 19864
rect 40132 18624 40184 18630
rect 40132 18566 40184 18572
rect 39684 18414 39804 18442
rect 39776 18290 39804 18414
rect 39764 18284 39816 18290
rect 39764 18226 39816 18232
rect 40040 18080 40092 18086
rect 40040 18022 40092 18028
rect 40052 17542 40080 18022
rect 38936 17536 38988 17542
rect 38936 17478 38988 17484
rect 39120 17536 39172 17542
rect 39120 17478 39172 17484
rect 40040 17536 40092 17542
rect 40040 17478 40092 17484
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 38672 16522 38700 17274
rect 38948 17202 38976 17478
rect 39132 17270 39160 17478
rect 40052 17338 40080 17478
rect 40040 17332 40092 17338
rect 40040 17274 40092 17280
rect 40144 17270 40172 18566
rect 40420 18057 40448 20998
rect 41050 20768 41106 20777
rect 41050 20703 41106 20712
rect 40684 20256 40736 20262
rect 40684 20198 40736 20204
rect 40590 19408 40646 19417
rect 40590 19343 40592 19352
rect 40644 19343 40646 19352
rect 40592 19314 40644 19320
rect 40500 19168 40552 19174
rect 40500 19110 40552 19116
rect 40512 18698 40540 19110
rect 40500 18692 40552 18698
rect 40500 18634 40552 18640
rect 40512 18086 40540 18634
rect 40500 18080 40552 18086
rect 40406 18048 40462 18057
rect 40500 18022 40552 18028
rect 40406 17983 40462 17992
rect 40696 17746 40724 20198
rect 41064 20058 41092 20703
rect 41156 20262 41184 22578
rect 41248 21894 41276 22986
rect 41418 22808 41474 22817
rect 41418 22743 41474 22752
rect 41236 21888 41288 21894
rect 41236 21830 41288 21836
rect 41328 21684 41380 21690
rect 41328 21626 41380 21632
rect 41340 20806 41368 21626
rect 41432 20913 41460 22743
rect 41616 22642 41644 23258
rect 41604 22636 41656 22642
rect 41604 22578 41656 22584
rect 41708 21894 41736 23802
rect 42168 23118 42196 24074
rect 42616 24064 42668 24070
rect 42616 24006 42668 24012
rect 42800 24064 42852 24070
rect 42800 24006 42852 24012
rect 42522 23896 42578 23905
rect 42522 23831 42524 23840
rect 42576 23831 42578 23840
rect 42524 23802 42576 23808
rect 42432 23520 42484 23526
rect 42432 23462 42484 23468
rect 42248 23248 42300 23254
rect 42444 23202 42472 23462
rect 42300 23196 42472 23202
rect 42248 23190 42472 23196
rect 42260 23174 42472 23190
rect 42156 23112 42208 23118
rect 42444 23089 42472 23174
rect 42156 23054 42208 23060
rect 42430 23080 42486 23089
rect 42430 23015 42486 23024
rect 42628 22642 42656 24006
rect 42812 23497 42840 24006
rect 42904 23526 42932 24278
rect 43364 24262 43484 24290
rect 43536 24278 43588 24284
rect 43352 24200 43404 24206
rect 43352 24142 43404 24148
rect 42982 23896 43038 23905
rect 42982 23831 43038 23840
rect 42996 23798 43024 23831
rect 42984 23792 43036 23798
rect 42984 23734 43036 23740
rect 42892 23520 42944 23526
rect 42798 23488 42854 23497
rect 42892 23462 42944 23468
rect 42798 23423 42854 23432
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 43364 23225 43392 24142
rect 43350 23216 43406 23225
rect 43350 23151 43406 23160
rect 43364 22982 43392 23151
rect 43352 22976 43404 22982
rect 43352 22918 43404 22924
rect 42798 22672 42854 22681
rect 42616 22636 42668 22642
rect 42798 22607 42854 22616
rect 42616 22578 42668 22584
rect 42812 22098 42840 22607
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 41972 22094 42024 22098
rect 42156 22094 42208 22098
rect 41972 22092 42208 22094
rect 42024 22066 42156 22092
rect 41972 22034 42024 22040
rect 42156 22034 42208 22040
rect 42800 22092 42852 22098
rect 43456 22094 43484 24262
rect 43548 24206 43576 24278
rect 43536 24200 43588 24206
rect 43536 24142 43588 24148
rect 43536 23588 43588 23594
rect 43536 23530 43588 23536
rect 43548 23322 43576 23530
rect 43628 23520 43680 23526
rect 43628 23462 43680 23468
rect 43640 23322 43668 23462
rect 43536 23316 43588 23322
rect 43536 23258 43588 23264
rect 43628 23316 43680 23322
rect 43628 23258 43680 23264
rect 42800 22034 42852 22040
rect 43364 22066 43484 22094
rect 42616 21956 42668 21962
rect 42800 21956 42852 21962
rect 42668 21916 42800 21944
rect 42616 21898 42668 21904
rect 42800 21898 42852 21904
rect 41696 21888 41748 21894
rect 41696 21830 41748 21836
rect 41512 21480 41564 21486
rect 41512 21422 41564 21428
rect 41418 20904 41474 20913
rect 41418 20839 41474 20848
rect 41328 20800 41380 20806
rect 41328 20742 41380 20748
rect 41144 20256 41196 20262
rect 41144 20198 41196 20204
rect 41052 20052 41104 20058
rect 41052 19994 41104 20000
rect 41064 19854 41092 19994
rect 41052 19848 41104 19854
rect 41052 19790 41104 19796
rect 40868 19712 40920 19718
rect 40868 19654 40920 19660
rect 40880 18426 40908 19654
rect 41340 19009 41368 20742
rect 41326 19000 41382 19009
rect 41524 18970 41552 21422
rect 41708 21146 41736 21830
rect 42616 21684 42668 21690
rect 42616 21626 42668 21632
rect 42628 21593 42656 21626
rect 42614 21584 42670 21593
rect 42432 21548 42484 21554
rect 43364 21554 43392 22066
rect 43444 22024 43496 22030
rect 43444 21966 43496 21972
rect 42614 21519 42670 21528
rect 43352 21548 43404 21554
rect 42432 21490 42484 21496
rect 43352 21490 43404 21496
rect 41696 21140 41748 21146
rect 41696 21082 41748 21088
rect 41326 18935 41382 18944
rect 41512 18964 41564 18970
rect 41512 18906 41564 18912
rect 40868 18420 40920 18426
rect 40868 18362 40920 18368
rect 41234 18184 41290 18193
rect 41234 18119 41290 18128
rect 40684 17740 40736 17746
rect 40684 17682 40736 17688
rect 40776 17672 40828 17678
rect 40776 17614 40828 17620
rect 40592 17604 40644 17610
rect 40592 17546 40644 17552
rect 39120 17264 39172 17270
rect 39120 17206 39172 17212
rect 40132 17264 40184 17270
rect 40132 17206 40184 17212
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 38844 16992 38896 16998
rect 38844 16934 38896 16940
rect 38856 16658 38884 16934
rect 38844 16652 38896 16658
rect 38844 16594 38896 16600
rect 38660 16516 38712 16522
rect 38660 16458 38712 16464
rect 38568 16448 38620 16454
rect 38568 16390 38620 16396
rect 38580 16182 38608 16390
rect 38672 16266 38700 16458
rect 38672 16238 38792 16266
rect 38764 16182 38792 16238
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38752 16176 38804 16182
rect 38752 16118 38804 16124
rect 38568 16040 38620 16046
rect 38568 15982 38620 15988
rect 38580 15366 38608 15982
rect 38764 15434 38792 16118
rect 38752 15428 38804 15434
rect 38752 15370 38804 15376
rect 38568 15360 38620 15366
rect 38568 15302 38620 15308
rect 38764 15094 38792 15370
rect 38752 15088 38804 15094
rect 38752 15030 38804 15036
rect 38476 14952 38528 14958
rect 38476 14894 38528 14900
rect 38764 14906 38792 15030
rect 38488 14618 38516 14894
rect 38764 14878 38884 14906
rect 38752 14816 38804 14822
rect 38752 14758 38804 14764
rect 38384 14612 38436 14618
rect 38384 14554 38436 14560
rect 38476 14612 38528 14618
rect 38476 14554 38528 14560
rect 38488 14278 38516 14554
rect 38476 14272 38528 14278
rect 38476 14214 38528 14220
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 38200 13796 38252 13802
rect 38200 13738 38252 13744
rect 38212 13530 38240 13738
rect 37832 13524 37884 13530
rect 37832 13466 37884 13472
rect 38200 13524 38252 13530
rect 38200 13466 38252 13472
rect 38212 13308 38240 13466
rect 38212 13280 38332 13308
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37648 13184 37700 13190
rect 37648 13126 37700 13132
rect 37188 12980 37240 12986
rect 37188 12922 37240 12928
rect 37200 12782 37228 12922
rect 37476 12850 37504 13126
rect 37660 12918 37688 13126
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37648 12912 37700 12918
rect 37648 12854 37700 12860
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 37188 12776 37240 12782
rect 37188 12718 37240 12724
rect 37096 12232 37148 12238
rect 37096 12174 37148 12180
rect 37280 12096 37332 12102
rect 37280 12038 37332 12044
rect 37292 10742 37320 12038
rect 37476 11218 37504 12786
rect 38304 12782 38332 13280
rect 38292 12776 38344 12782
rect 38292 12718 38344 12724
rect 38764 12306 38792 14758
rect 38856 14618 38884 14878
rect 38844 14612 38896 14618
rect 38844 14554 38896 14560
rect 38856 14346 38884 14554
rect 38844 14340 38896 14346
rect 38844 14282 38896 14288
rect 38856 14006 38884 14282
rect 38844 14000 38896 14006
rect 38844 13942 38896 13948
rect 38856 13530 38884 13942
rect 38844 13524 38896 13530
rect 38844 13466 38896 13472
rect 38856 13258 38884 13466
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 38856 12850 38884 13194
rect 38844 12844 38896 12850
rect 38844 12786 38896 12792
rect 38384 12300 38436 12306
rect 38384 12242 38436 12248
rect 38752 12300 38804 12306
rect 38752 12242 38804 12248
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 38396 11626 38424 12242
rect 38660 12096 38712 12102
rect 38660 12038 38712 12044
rect 38672 11898 38700 12038
rect 38660 11892 38712 11898
rect 38660 11834 38712 11840
rect 38384 11620 38436 11626
rect 38384 11562 38436 11568
rect 37464 11212 37516 11218
rect 37464 11154 37516 11160
rect 38396 11082 38424 11562
rect 38660 11348 38712 11354
rect 38660 11290 38712 11296
rect 38384 11076 38436 11082
rect 38384 11018 38436 11024
rect 38672 10996 38700 11290
rect 38580 10968 38700 10996
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 37280 10736 37332 10742
rect 37280 10678 37332 10684
rect 38580 10470 38608 10968
rect 38948 10538 38976 17138
rect 40224 16788 40276 16794
rect 40224 16730 40276 16736
rect 40236 16697 40264 16730
rect 40222 16688 40278 16697
rect 40222 16623 40278 16632
rect 40316 16652 40368 16658
rect 39488 16584 39540 16590
rect 39488 16526 39540 16532
rect 39946 16552 40002 16561
rect 39500 15570 39528 16526
rect 40236 16522 40264 16623
rect 40316 16594 40368 16600
rect 39946 16487 40002 16496
rect 40224 16516 40276 16522
rect 39488 15564 39540 15570
rect 39488 15506 39540 15512
rect 39960 15162 39988 16487
rect 40224 16458 40276 16464
rect 40328 15910 40356 16594
rect 40316 15904 40368 15910
rect 40316 15846 40368 15852
rect 40328 15570 40356 15846
rect 40316 15564 40368 15570
rect 40316 15506 40368 15512
rect 39948 15156 40000 15162
rect 39948 15098 40000 15104
rect 40604 15094 40632 17546
rect 40684 17128 40736 17134
rect 40684 17070 40736 17076
rect 40696 16590 40724 17070
rect 40788 16998 40816 17614
rect 41052 17332 41104 17338
rect 41052 17274 41104 17280
rect 40776 16992 40828 16998
rect 40776 16934 40828 16940
rect 41064 16794 41092 17274
rect 41248 16794 41276 18119
rect 41708 16998 41736 21082
rect 42444 21010 42472 21490
rect 42800 21344 42852 21350
rect 42800 21286 42852 21292
rect 42432 21004 42484 21010
rect 42432 20946 42484 20952
rect 42812 20330 42840 21286
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 43364 21078 43392 21490
rect 43352 21072 43404 21078
rect 43352 21014 43404 21020
rect 43352 20800 43404 20806
rect 43352 20742 43404 20748
rect 42800 20324 42852 20330
rect 42800 20266 42852 20272
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 43364 19990 43392 20742
rect 43352 19984 43404 19990
rect 43352 19926 43404 19932
rect 42064 19168 42116 19174
rect 42064 19110 42116 19116
rect 42076 18970 42104 19110
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42064 18964 42116 18970
rect 42064 18906 42116 18912
rect 41880 18896 41932 18902
rect 41880 18838 41932 18844
rect 41892 17241 41920 18838
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 43456 17542 43484 21966
rect 43536 21344 43588 21350
rect 43536 21286 43588 21292
rect 43548 21146 43576 21286
rect 43536 21140 43588 21146
rect 43536 21082 43588 21088
rect 43640 20602 43668 23258
rect 43810 22536 43866 22545
rect 43810 22471 43866 22480
rect 43824 21554 43852 22471
rect 43812 21548 43864 21554
rect 43812 21490 43864 21496
rect 43824 21146 43852 21490
rect 43812 21140 43864 21146
rect 43812 21082 43864 21088
rect 43916 20602 43944 24686
rect 43994 24304 44050 24313
rect 43994 24239 44050 24248
rect 44008 23594 44036 24239
rect 43996 23588 44048 23594
rect 43996 23530 44048 23536
rect 44100 22710 44128 26200
rect 44364 24676 44416 24682
rect 44364 24618 44416 24624
rect 44272 24404 44324 24410
rect 44272 24346 44324 24352
rect 44180 24064 44232 24070
rect 44180 24006 44232 24012
rect 44192 23118 44220 24006
rect 44284 23254 44312 24346
rect 44272 23248 44324 23254
rect 44272 23190 44324 23196
rect 44180 23112 44232 23118
rect 44180 23054 44232 23060
rect 44088 22704 44140 22710
rect 44088 22646 44140 22652
rect 44180 22636 44232 22642
rect 44180 22578 44232 22584
rect 43996 22568 44048 22574
rect 43996 22510 44048 22516
rect 43628 20596 43680 20602
rect 43628 20538 43680 20544
rect 43904 20596 43956 20602
rect 43904 20538 43956 20544
rect 44008 19961 44036 22510
rect 44192 22030 44220 22578
rect 44180 22024 44232 22030
rect 44180 21966 44232 21972
rect 44272 21480 44324 21486
rect 44272 21422 44324 21428
rect 44180 20868 44232 20874
rect 44180 20810 44232 20816
rect 44192 19990 44220 20810
rect 44180 19984 44232 19990
rect 43994 19952 44050 19961
rect 44180 19926 44232 19932
rect 43994 19887 44050 19896
rect 44284 19281 44312 21422
rect 44376 21078 44404 24618
rect 44456 24200 44508 24206
rect 44456 24142 44508 24148
rect 44468 22778 44496 24142
rect 44744 24138 44772 26200
rect 45388 24698 45416 26200
rect 46202 25120 46258 25129
rect 46202 25055 46258 25064
rect 45388 24682 45600 24698
rect 45388 24676 45612 24682
rect 45388 24670 45560 24676
rect 45560 24618 45612 24624
rect 44732 24132 44784 24138
rect 44732 24074 44784 24080
rect 44640 24064 44692 24070
rect 44640 24006 44692 24012
rect 45376 24064 45428 24070
rect 45376 24006 45428 24012
rect 44548 23316 44600 23322
rect 44548 23258 44600 23264
rect 44560 23118 44588 23258
rect 44548 23112 44600 23118
rect 44548 23054 44600 23060
rect 44456 22772 44508 22778
rect 44456 22714 44508 22720
rect 44548 22500 44600 22506
rect 44548 22442 44600 22448
rect 44560 22098 44588 22442
rect 44548 22092 44600 22098
rect 44548 22034 44600 22040
rect 44456 21684 44508 21690
rect 44456 21626 44508 21632
rect 44468 21146 44496 21626
rect 44652 21622 44680 24006
rect 44824 23724 44876 23730
rect 44824 23666 44876 23672
rect 44732 23520 44784 23526
rect 44732 23462 44784 23468
rect 44744 23050 44772 23462
rect 44836 23322 44864 23666
rect 44824 23316 44876 23322
rect 44824 23258 44876 23264
rect 45388 23118 45416 24006
rect 46020 23588 46072 23594
rect 46020 23530 46072 23536
rect 45376 23112 45428 23118
rect 45376 23054 45428 23060
rect 44732 23044 44784 23050
rect 44732 22986 44784 22992
rect 45742 22808 45798 22817
rect 45742 22743 45798 22752
rect 45756 22710 45784 22743
rect 44732 22704 44784 22710
rect 44732 22646 44784 22652
rect 45744 22704 45796 22710
rect 45744 22646 45796 22652
rect 44744 22234 44772 22646
rect 45008 22500 45060 22506
rect 45008 22442 45060 22448
rect 44732 22228 44784 22234
rect 44732 22170 44784 22176
rect 45020 21894 45048 22442
rect 45284 22432 45336 22438
rect 45284 22374 45336 22380
rect 45296 22166 45324 22374
rect 45284 22160 45336 22166
rect 45190 22128 45246 22137
rect 45284 22102 45336 22108
rect 45190 22063 45192 22072
rect 45244 22063 45246 22072
rect 45192 22034 45244 22040
rect 45008 21888 45060 21894
rect 45008 21830 45060 21836
rect 44640 21616 44692 21622
rect 44640 21558 44692 21564
rect 45204 21554 45232 22034
rect 45468 22024 45520 22030
rect 45468 21966 45520 21972
rect 45192 21548 45244 21554
rect 45192 21490 45244 21496
rect 45190 21448 45246 21457
rect 45190 21383 45246 21392
rect 45204 21146 45232 21383
rect 44456 21140 44508 21146
rect 44456 21082 44508 21088
rect 45192 21140 45244 21146
rect 45192 21082 45244 21088
rect 44364 21072 44416 21078
rect 44364 21014 44416 21020
rect 45376 21072 45428 21078
rect 45480 21049 45508 21966
rect 45836 21956 45888 21962
rect 45836 21898 45888 21904
rect 45848 21146 45876 21898
rect 45836 21140 45888 21146
rect 45836 21082 45888 21088
rect 45376 21014 45428 21020
rect 45466 21040 45522 21049
rect 45388 20942 45416 21014
rect 45466 20975 45522 20984
rect 45376 20936 45428 20942
rect 45376 20878 45428 20884
rect 46032 19854 46060 23530
rect 46216 20602 46244 25055
rect 46308 24410 46336 26302
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 49238 26330 49294 27000
rect 49160 26302 49294 26330
rect 46570 24712 46626 24721
rect 46570 24647 46626 24656
rect 46296 24404 46348 24410
rect 46296 24346 46348 24352
rect 46478 23760 46534 23769
rect 46388 23724 46440 23730
rect 46478 23695 46534 23704
rect 46388 23666 46440 23672
rect 46296 21412 46348 21418
rect 46296 21354 46348 21360
rect 46204 20596 46256 20602
rect 46204 20538 46256 20544
rect 46216 20398 46244 20538
rect 46308 20505 46336 21354
rect 46294 20496 46350 20505
rect 46294 20431 46350 20440
rect 46204 20392 46256 20398
rect 46204 20334 46256 20340
rect 46400 20058 46428 23666
rect 46492 20602 46520 23695
rect 46584 21978 46612 24647
rect 46676 22574 46704 26200
rect 46846 25528 46902 25537
rect 46846 25463 46902 25472
rect 46756 24676 46808 24682
rect 46756 24618 46808 24624
rect 46768 24342 46796 24618
rect 46756 24336 46808 24342
rect 46756 24278 46808 24284
rect 46860 23730 46888 25463
rect 47124 24608 47176 24614
rect 47124 24550 47176 24556
rect 46848 23724 46900 23730
rect 46848 23666 46900 23672
rect 46846 23488 46902 23497
rect 46846 23423 46902 23432
rect 46756 22976 46808 22982
rect 46756 22918 46808 22924
rect 46664 22568 46716 22574
rect 46664 22510 46716 22516
rect 46768 22030 46796 22918
rect 46860 22098 46888 23423
rect 47032 23248 47084 23254
rect 47032 23190 47084 23196
rect 47044 22234 47072 23190
rect 47032 22228 47084 22234
rect 47032 22170 47084 22176
rect 46848 22092 46900 22098
rect 46848 22034 46900 22040
rect 46756 22024 46808 22030
rect 46584 21950 46704 21978
rect 46756 21966 46808 21972
rect 46572 21888 46624 21894
rect 46572 21830 46624 21836
rect 46480 20596 46532 20602
rect 46480 20538 46532 20544
rect 46492 20466 46520 20538
rect 46480 20460 46532 20466
rect 46480 20402 46532 20408
rect 46584 20369 46612 21830
rect 46570 20360 46626 20369
rect 46570 20295 46626 20304
rect 46388 20052 46440 20058
rect 46388 19994 46440 20000
rect 46020 19848 46072 19854
rect 46020 19790 46072 19796
rect 46676 19718 46704 21950
rect 46860 21078 46888 22034
rect 47044 21622 47072 22170
rect 47032 21616 47084 21622
rect 47032 21558 47084 21564
rect 46848 21072 46900 21078
rect 46848 21014 46900 21020
rect 46848 20596 46900 20602
rect 46848 20538 46900 20544
rect 46860 19854 46888 20538
rect 47032 20256 47084 20262
rect 47032 20198 47084 20204
rect 46848 19848 46900 19854
rect 46848 19790 46900 19796
rect 46664 19712 46716 19718
rect 46664 19654 46716 19660
rect 44270 19272 44326 19281
rect 44270 19207 44326 19216
rect 46676 19174 46704 19654
rect 47044 19378 47072 20198
rect 47136 20058 47164 24550
rect 47320 23866 47348 26200
rect 47964 24562 47992 26200
rect 47412 24534 47992 24562
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 47320 22710 47348 23802
rect 47308 22704 47360 22710
rect 47308 22646 47360 22652
rect 47412 21554 47440 24534
rect 47860 24404 47912 24410
rect 47860 24346 47912 24352
rect 47676 24200 47728 24206
rect 47676 24142 47728 24148
rect 47584 23112 47636 23118
rect 47584 23054 47636 23060
rect 47596 22778 47624 23054
rect 47584 22772 47636 22778
rect 47584 22714 47636 22720
rect 47584 22568 47636 22574
rect 47584 22510 47636 22516
rect 47492 21956 47544 21962
rect 47492 21898 47544 21904
rect 47400 21548 47452 21554
rect 47400 21490 47452 21496
rect 47216 21412 47268 21418
rect 47216 21354 47268 21360
rect 47228 20466 47256 21354
rect 47412 21350 47440 21490
rect 47400 21344 47452 21350
rect 47400 21286 47452 21292
rect 47308 20800 47360 20806
rect 47400 20800 47452 20806
rect 47308 20742 47360 20748
rect 47398 20768 47400 20777
rect 47452 20768 47454 20777
rect 47216 20460 47268 20466
rect 47216 20402 47268 20408
rect 47124 20052 47176 20058
rect 47124 19994 47176 20000
rect 47032 19372 47084 19378
rect 47032 19314 47084 19320
rect 46664 19168 46716 19174
rect 46664 19110 46716 19116
rect 47320 18873 47348 20742
rect 47398 20703 47454 20712
rect 47504 18970 47532 21898
rect 47596 21554 47624 22510
rect 47688 22098 47716 24142
rect 47766 23080 47822 23089
rect 47766 23015 47822 23024
rect 47676 22092 47728 22098
rect 47676 22034 47728 22040
rect 47674 21584 47730 21593
rect 47584 21548 47636 21554
rect 47674 21519 47730 21528
rect 47584 21490 47636 21496
rect 47688 20602 47716 21519
rect 47780 21486 47808 23015
rect 47872 22710 47900 24346
rect 48042 24168 48098 24177
rect 48042 24103 48098 24112
rect 48056 24070 48084 24103
rect 48044 24064 48096 24070
rect 48044 24006 48096 24012
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 48228 23724 48280 23730
rect 48228 23666 48280 23672
rect 48044 23520 48096 23526
rect 48044 23462 48096 23468
rect 48056 23186 48084 23462
rect 48240 23322 48268 23666
rect 48228 23316 48280 23322
rect 48228 23258 48280 23264
rect 48608 23254 48636 26200
rect 48780 24064 48832 24070
rect 48780 24006 48832 24012
rect 48596 23248 48648 23254
rect 48596 23190 48648 23196
rect 48044 23180 48096 23186
rect 48044 23122 48096 23128
rect 48056 23089 48084 23122
rect 48042 23080 48098 23089
rect 48042 23015 48098 23024
rect 48320 22976 48372 22982
rect 48320 22918 48372 22924
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47860 22704 47912 22710
rect 47860 22646 47912 22652
rect 47860 22568 47912 22574
rect 47860 22510 47912 22516
rect 47768 21480 47820 21486
rect 47768 21422 47820 21428
rect 47872 20942 47900 22510
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 48332 21010 48360 22918
rect 48688 21888 48740 21894
rect 48688 21830 48740 21836
rect 48700 21622 48728 21830
rect 48688 21616 48740 21622
rect 48688 21558 48740 21564
rect 48320 21004 48372 21010
rect 48320 20946 48372 20952
rect 47860 20936 47912 20942
rect 47860 20878 47912 20884
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47676 20596 47728 20602
rect 47676 20538 47728 20544
rect 48410 20224 48466 20233
rect 48410 20159 48466 20168
rect 47584 19848 47636 19854
rect 47584 19790 47636 19796
rect 47596 19446 47624 19790
rect 47676 19780 47728 19786
rect 47676 19722 47728 19728
rect 47584 19440 47636 19446
rect 47584 19382 47636 19388
rect 47492 18964 47544 18970
rect 47492 18906 47544 18912
rect 47306 18864 47362 18873
rect 47306 18799 47362 18808
rect 47308 18624 47360 18630
rect 47308 18566 47360 18572
rect 47320 18358 47348 18566
rect 47308 18352 47360 18358
rect 47308 18294 47360 18300
rect 47688 18193 47716 19722
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 48424 19514 48452 20159
rect 48412 19508 48464 19514
rect 48412 19450 48464 19456
rect 48412 18828 48464 18834
rect 48412 18770 48464 18776
rect 48424 18601 48452 18770
rect 48410 18592 48466 18601
rect 47950 18524 48258 18533
rect 48410 18527 48466 18536
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 48424 18426 48452 18527
rect 48412 18420 48464 18426
rect 48412 18362 48464 18368
rect 47674 18184 47730 18193
rect 47674 18119 47730 18128
rect 48044 18080 48096 18086
rect 48044 18022 48096 18028
rect 46940 17808 46992 17814
rect 46938 17776 46940 17785
rect 46992 17776 46994 17785
rect 46938 17711 46994 17720
rect 48056 17649 48084 18022
rect 48042 17640 48098 17649
rect 47032 17604 47084 17610
rect 48042 17575 48098 17584
rect 47032 17546 47084 17552
rect 43444 17536 43496 17542
rect 43444 17478 43496 17484
rect 47044 17338 47072 17546
rect 47676 17536 47728 17542
rect 47676 17478 47728 17484
rect 47032 17332 47084 17338
rect 47032 17274 47084 17280
rect 47688 17270 47716 17478
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 47676 17264 47728 17270
rect 41878 17232 41934 17241
rect 47676 17206 47728 17212
rect 48228 17264 48280 17270
rect 48228 17206 48280 17212
rect 41878 17167 41934 17176
rect 47952 17128 48004 17134
rect 47950 17096 47952 17105
rect 48004 17096 48006 17105
rect 47950 17031 48006 17040
rect 41696 16992 41748 16998
rect 41696 16934 41748 16940
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 41052 16788 41104 16794
rect 41052 16730 41104 16736
rect 41236 16788 41288 16794
rect 41236 16730 41288 16736
rect 41064 16658 41092 16730
rect 41052 16652 41104 16658
rect 41052 16594 41104 16600
rect 40684 16584 40736 16590
rect 40684 16526 40736 16532
rect 40960 16448 41012 16454
rect 40960 16390 41012 16396
rect 40972 16250 41000 16390
rect 40960 16244 41012 16250
rect 40960 16186 41012 16192
rect 41064 15434 41092 16594
rect 41248 16522 41276 16730
rect 48240 16561 48268 17206
rect 48320 16992 48372 16998
rect 48318 16960 48320 16969
rect 48372 16960 48374 16969
rect 48318 16895 48374 16904
rect 48792 16726 48820 24006
rect 49160 23866 49188 26302
rect 49238 26200 49294 26302
rect 49514 24304 49570 24313
rect 49514 24239 49570 24248
rect 49528 23866 49556 24239
rect 49148 23860 49200 23866
rect 49148 23802 49200 23808
rect 49516 23860 49568 23866
rect 49516 23802 49568 23808
rect 49160 22642 49188 23802
rect 49332 23520 49384 23526
rect 49332 23462 49384 23468
rect 49344 23118 49372 23462
rect 49332 23112 49384 23118
rect 49332 23054 49384 23060
rect 49344 22681 49372 23054
rect 49330 22672 49386 22681
rect 49148 22636 49200 22642
rect 49148 22578 49200 22584
rect 49240 22636 49292 22642
rect 49330 22607 49386 22616
rect 49240 22578 49292 22584
rect 49252 22273 49280 22578
rect 49238 22264 49294 22273
rect 49238 22199 49294 22208
rect 49252 21690 49280 22199
rect 49528 22098 49556 23802
rect 49516 22092 49568 22098
rect 49516 22034 49568 22040
rect 49332 22024 49384 22030
rect 49332 21966 49384 21972
rect 49240 21684 49292 21690
rect 49240 21626 49292 21632
rect 49240 21548 49292 21554
rect 49240 21490 49292 21496
rect 49252 21049 49280 21490
rect 49344 21457 49372 21966
rect 49330 21448 49386 21457
rect 49330 21383 49386 21392
rect 49238 21040 49294 21049
rect 49238 20975 49294 20984
rect 49252 19922 49280 20975
rect 49332 20936 49384 20942
rect 49332 20878 49384 20884
rect 49344 20641 49372 20878
rect 49330 20632 49386 20641
rect 49330 20567 49386 20576
rect 49332 20460 49384 20466
rect 49332 20402 49384 20408
rect 49344 20330 49372 20402
rect 49332 20324 49384 20330
rect 49332 20266 49384 20272
rect 49240 19916 49292 19922
rect 49240 19858 49292 19864
rect 49344 19825 49372 20266
rect 49424 19848 49476 19854
rect 49330 19816 49386 19825
rect 49424 19790 49476 19796
rect 49330 19751 49386 19760
rect 49436 19417 49464 19790
rect 49422 19408 49478 19417
rect 49332 19372 49384 19378
rect 49422 19343 49478 19352
rect 49332 19314 49384 19320
rect 49344 19009 49372 19314
rect 49330 19000 49386 19009
rect 49330 18935 49386 18944
rect 49424 18760 49476 18766
rect 49424 18702 49476 18708
rect 49332 18284 49384 18290
rect 49332 18226 49384 18232
rect 49344 17785 49372 18226
rect 49436 18193 49464 18702
rect 49422 18184 49478 18193
rect 49422 18119 49478 18128
rect 49330 17776 49386 17785
rect 49330 17711 49386 17720
rect 49332 17672 49384 17678
rect 49332 17614 49384 17620
rect 49344 17377 49372 17614
rect 49330 17368 49386 17377
rect 49330 17303 49386 17312
rect 48780 16720 48832 16726
rect 48780 16662 48832 16668
rect 49332 16584 49384 16590
rect 48226 16552 48282 16561
rect 41236 16516 41288 16522
rect 49332 16526 49384 16532
rect 48226 16487 48282 16496
rect 41236 16458 41288 16464
rect 41604 16448 41656 16454
rect 41604 16390 41656 16396
rect 47860 16448 47912 16454
rect 47860 16390 47912 16396
rect 41616 15910 41644 16390
rect 41788 16040 41840 16046
rect 41788 15982 41840 15988
rect 41604 15904 41656 15910
rect 41604 15846 41656 15852
rect 41616 15706 41644 15846
rect 41604 15700 41656 15706
rect 41604 15642 41656 15648
rect 41800 15638 41828 15982
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 41788 15632 41840 15638
rect 41788 15574 41840 15580
rect 47872 15473 47900 16390
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 49344 16153 49372 16526
rect 49330 16144 49386 16153
rect 48320 16108 48372 16114
rect 48320 16050 48372 16056
rect 48688 16108 48740 16114
rect 49330 16079 49386 16088
rect 48688 16050 48740 16056
rect 48332 15706 48360 16050
rect 48700 15745 48728 16050
rect 49146 16008 49202 16017
rect 49146 15943 49202 15952
rect 48686 15736 48742 15745
rect 48320 15700 48372 15706
rect 49160 15706 49188 15943
rect 49332 15904 49384 15910
rect 49332 15846 49384 15852
rect 48686 15671 48742 15680
rect 49148 15700 49200 15706
rect 48320 15642 48372 15648
rect 49148 15642 49200 15648
rect 49344 15502 49372 15846
rect 48596 15496 48648 15502
rect 47858 15464 47914 15473
rect 41052 15428 41104 15434
rect 48596 15438 48648 15444
rect 49332 15496 49384 15502
rect 49332 15438 49384 15444
rect 47858 15399 47914 15408
rect 41052 15370 41104 15376
rect 48608 15337 48636 15438
rect 48594 15328 48650 15337
rect 47950 15260 48258 15269
rect 48594 15263 48650 15272
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 40592 15088 40644 15094
rect 40592 15030 40644 15036
rect 47858 15056 47914 15065
rect 47858 14991 47914 15000
rect 49332 15020 49384 15026
rect 40224 14952 40276 14958
rect 40224 14894 40276 14900
rect 46940 14952 46992 14958
rect 46940 14894 46992 14900
rect 39302 14512 39358 14521
rect 39302 14447 39358 14456
rect 39316 14414 39344 14447
rect 39304 14408 39356 14414
rect 39304 14350 39356 14356
rect 39488 14272 39540 14278
rect 39488 14214 39540 14220
rect 39500 14006 39528 14214
rect 39488 14000 39540 14006
rect 39488 13942 39540 13948
rect 40236 13938 40264 14894
rect 45652 14816 45704 14822
rect 45652 14758 45704 14764
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 41328 14068 41380 14074
rect 41328 14010 41380 14016
rect 40224 13932 40276 13938
rect 40224 13874 40276 13880
rect 39488 13524 39540 13530
rect 39488 13466 39540 13472
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39316 12782 39344 13126
rect 39304 12776 39356 12782
rect 39304 12718 39356 12724
rect 39120 12640 39172 12646
rect 39120 12582 39172 12588
rect 39132 11898 39160 12582
rect 39316 12442 39344 12718
rect 39500 12442 39528 13466
rect 39580 13388 39632 13394
rect 39580 13330 39632 13336
rect 39304 12436 39356 12442
rect 39304 12378 39356 12384
rect 39488 12436 39540 12442
rect 39488 12378 39540 12384
rect 39120 11892 39172 11898
rect 39120 11834 39172 11840
rect 39028 11756 39080 11762
rect 39028 11698 39080 11704
rect 38936 10532 38988 10538
rect 38936 10474 38988 10480
rect 38568 10464 38620 10470
rect 38568 10406 38620 10412
rect 38948 10062 38976 10474
rect 38936 10056 38988 10062
rect 38936 9998 38988 10004
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37832 8832 37884 8838
rect 37832 8774 37884 8780
rect 37844 8566 37872 8774
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 37832 8560 37884 8566
rect 37832 8502 37884 8508
rect 38752 8356 38804 8362
rect 38752 8298 38804 8304
rect 38764 7818 38792 8298
rect 39040 7886 39068 11698
rect 39500 11354 39528 12378
rect 39592 11354 39620 13330
rect 41340 13326 41368 14010
rect 45664 13938 45692 14758
rect 45652 13932 45704 13938
rect 45652 13874 45704 13880
rect 46952 13870 46980 14894
rect 47216 14068 47268 14074
rect 47216 14010 47268 14016
rect 46756 13864 46808 13870
rect 46756 13806 46808 13812
rect 46940 13864 46992 13870
rect 46940 13806 46992 13812
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 46768 13326 46796 13806
rect 41328 13320 41380 13326
rect 41328 13262 41380 13268
rect 46756 13320 46808 13326
rect 46756 13262 46808 13268
rect 45928 13184 45980 13190
rect 45928 13126 45980 13132
rect 40316 12980 40368 12986
rect 40316 12922 40368 12928
rect 40040 12844 40092 12850
rect 40040 12786 40092 12792
rect 40052 12753 40080 12786
rect 40038 12744 40094 12753
rect 40038 12679 40094 12688
rect 39948 12368 40000 12374
rect 39948 12310 40000 12316
rect 39960 11830 39988 12310
rect 39948 11824 40000 11830
rect 39948 11766 40000 11772
rect 40224 11552 40276 11558
rect 40224 11494 40276 11500
rect 39488 11348 39540 11354
rect 39488 11290 39540 11296
rect 39580 11348 39632 11354
rect 39580 11290 39632 11296
rect 39592 11150 39620 11290
rect 40236 11150 40264 11494
rect 39580 11144 39632 11150
rect 39580 11086 39632 11092
rect 40224 11144 40276 11150
rect 40224 11086 40276 11092
rect 39396 8968 39448 8974
rect 39396 8910 39448 8916
rect 39408 8430 39436 8910
rect 40040 8628 40092 8634
rect 40040 8570 40092 8576
rect 39396 8424 39448 8430
rect 39396 8366 39448 8372
rect 39028 7880 39080 7886
rect 39028 7822 39080 7828
rect 38752 7812 38804 7818
rect 38752 7754 38804 7760
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 38672 7478 38700 7686
rect 38660 7472 38712 7478
rect 38660 7414 38712 7420
rect 37280 7200 37332 7206
rect 37280 7142 37332 7148
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 36820 6316 36872 6322
rect 36820 6258 36872 6264
rect 37004 6316 37056 6322
rect 37004 6258 37056 6264
rect 36832 4826 36860 6258
rect 37292 5302 37320 7142
rect 37936 6934 37964 7142
rect 38476 6996 38528 7002
rect 38476 6938 38528 6944
rect 37924 6928 37976 6934
rect 37924 6870 37976 6876
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37740 6248 37792 6254
rect 37740 6190 37792 6196
rect 37648 6112 37700 6118
rect 37648 6054 37700 6060
rect 37660 5914 37688 6054
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37280 5296 37332 5302
rect 37280 5238 37332 5244
rect 36452 4820 36504 4826
rect 36452 4762 36504 4768
rect 36820 4820 36872 4826
rect 36820 4762 36872 4768
rect 35072 4072 35124 4078
rect 35072 4014 35124 4020
rect 35084 2854 35112 4014
rect 36464 3534 36492 4762
rect 36832 4622 36860 4762
rect 37752 4622 37780 6190
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 38488 5302 38516 6938
rect 40052 6390 40080 8570
rect 40328 8498 40356 12922
rect 45940 12850 45968 13126
rect 47228 12850 47256 14010
rect 47872 14006 47900 14991
rect 49332 14962 49384 14968
rect 49344 14929 49372 14962
rect 48042 14920 48098 14929
rect 48042 14855 48044 14864
rect 48096 14855 48098 14864
rect 49330 14920 49386 14929
rect 49330 14855 49386 14864
rect 48044 14826 48096 14832
rect 49330 14512 49386 14521
rect 49330 14447 49386 14456
rect 49344 14414 49372 14447
rect 47952 14408 48004 14414
rect 47950 14376 47952 14385
rect 49332 14408 49384 14414
rect 48004 14376 48006 14385
rect 49332 14350 49384 14356
rect 47950 14311 48006 14320
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 49330 14104 49386 14113
rect 49330 14039 49386 14048
rect 47860 14000 47912 14006
rect 47860 13942 47912 13948
rect 49344 13938 49372 14039
rect 49332 13932 49384 13938
rect 49332 13874 49384 13880
rect 47676 13864 47728 13870
rect 47676 13806 47728 13812
rect 47768 13864 47820 13870
rect 47768 13806 47820 13812
rect 47688 13705 47716 13806
rect 47674 13696 47730 13705
rect 47674 13631 47730 13640
rect 47780 13530 47808 13806
rect 47768 13524 47820 13530
rect 47768 13466 47820 13472
rect 49148 13320 49200 13326
rect 49146 13288 49148 13297
rect 49200 13288 49202 13297
rect 49146 13223 49202 13232
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 49146 12880 49202 12889
rect 45928 12844 45980 12850
rect 45928 12786 45980 12792
rect 47216 12844 47268 12850
rect 49146 12815 49148 12824
rect 47216 12786 47268 12792
rect 49200 12815 49202 12824
rect 49148 12786 49200 12792
rect 46940 12708 46992 12714
rect 46940 12650 46992 12656
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 40408 12164 40460 12170
rect 40408 12106 40460 12112
rect 40420 11830 40448 12106
rect 40960 12096 41012 12102
rect 40960 12038 41012 12044
rect 46112 12096 46164 12102
rect 46112 12038 46164 12044
rect 40972 11830 41000 12038
rect 40408 11824 40460 11830
rect 40406 11792 40408 11801
rect 40960 11824 41012 11830
rect 40460 11792 40462 11801
rect 40960 11766 41012 11772
rect 46124 11762 46152 12038
rect 40406 11727 40462 11736
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 46664 11620 46716 11626
rect 46664 11562 46716 11568
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 44364 11348 44416 11354
rect 44364 11290 44416 11296
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 44376 9994 44404 11290
rect 46112 11008 46164 11014
rect 46112 10950 46164 10956
rect 46124 10062 46152 10950
rect 46676 10062 46704 11562
rect 46952 11150 46980 12650
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 47400 12368 47452 12374
rect 47400 12310 47452 12316
rect 47032 11552 47084 11558
rect 47032 11494 47084 11500
rect 46940 11144 46992 11150
rect 46940 11086 46992 11092
rect 46940 10532 46992 10538
rect 46940 10474 46992 10480
rect 45836 10056 45888 10062
rect 45836 9998 45888 10004
rect 46112 10056 46164 10062
rect 46112 9998 46164 10004
rect 46664 10056 46716 10062
rect 46664 9998 46716 10004
rect 44364 9988 44416 9994
rect 44364 9930 44416 9936
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 43720 9172 43772 9178
rect 43720 9114 43772 9120
rect 40316 8492 40368 8498
rect 40316 8434 40368 8440
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 40592 7812 40644 7818
rect 40592 7754 40644 7760
rect 40604 6798 40632 7754
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 40592 6792 40644 6798
rect 40592 6734 40644 6740
rect 40040 6384 40092 6390
rect 40040 6326 40092 6332
rect 39212 6180 39264 6186
rect 39212 6122 39264 6128
rect 38476 5296 38528 5302
rect 38476 5238 38528 5244
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 37844 4826 37872 4966
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 36820 4616 36872 4622
rect 36820 4558 36872 4564
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 37372 4480 37424 4486
rect 37372 4422 37424 4428
rect 37384 4282 37412 4422
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 36556 3738 36584 4082
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 36452 3528 36504 3534
rect 36452 3470 36504 3476
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 35256 3052 35308 3058
rect 35256 2994 35308 3000
rect 35072 2848 35124 2854
rect 35072 2790 35124 2796
rect 35268 2650 35296 2994
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 38304 2650 38332 2926
rect 35256 2644 35308 2650
rect 35256 2586 35308 2592
rect 38292 2644 38344 2650
rect 38292 2586 38344 2592
rect 34152 2576 34204 2582
rect 34152 2518 34204 2524
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 29552 2508 29604 2514
rect 29552 2450 29604 2456
rect 27160 2440 27212 2446
rect 29012 2394 29040 2450
rect 27160 2382 27212 2388
rect 28920 2366 29040 2394
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28644 870 28764 898
rect 28644 800 28672 870
rect 18156 734 18368 762
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 28736 762 28764 870
rect 28920 762 28948 2366
rect 30760 800 30788 2382
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 32876 800 32904 2246
rect 34992 800 35020 2246
rect 37108 800 37136 2246
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 39224 800 39252 6122
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43732 5710 43760 9114
rect 45848 8498 45876 9998
rect 46756 9988 46808 9994
rect 46756 9930 46808 9936
rect 46480 8968 46532 8974
rect 46480 8910 46532 8916
rect 45836 8492 45888 8498
rect 45836 8434 45888 8440
rect 44916 8356 44968 8362
rect 44916 8298 44968 8304
rect 44928 7410 44956 8298
rect 44916 7404 44968 7410
rect 44916 7346 44968 7352
rect 45744 7200 45796 7206
rect 45744 7142 45796 7148
rect 43720 5704 43772 5710
rect 43720 5646 43772 5652
rect 45652 5636 45704 5642
rect 45652 5578 45704 5584
rect 40040 5092 40092 5098
rect 40040 5034 40092 5040
rect 39764 4548 39816 4554
rect 39764 4490 39816 4496
rect 39776 3058 39804 4490
rect 40052 3534 40080 5034
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 45560 3460 45612 3466
rect 45560 3402 45612 3408
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 40684 2916 40736 2922
rect 40684 2858 40736 2864
rect 40696 2446 40724 2858
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 40684 2440 40736 2446
rect 40684 2382 40736 2388
rect 41340 800 41368 2450
rect 43444 2304 43496 2310
rect 43444 2246 43496 2252
rect 43456 800 43484 2246
rect 45572 800 45600 3402
rect 45664 3058 45692 5578
rect 45756 5234 45784 7142
rect 45744 5228 45796 5234
rect 45744 5170 45796 5176
rect 46492 4758 46520 8910
rect 46768 8498 46796 9930
rect 46756 8492 46808 8498
rect 46756 8434 46808 8440
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46860 7993 46888 8366
rect 46846 7984 46902 7993
rect 46846 7919 46902 7928
rect 46952 7886 46980 10474
rect 47044 8974 47072 11494
rect 47216 11076 47268 11082
rect 47216 11018 47268 11024
rect 47228 10674 47256 11018
rect 47216 10668 47268 10674
rect 47216 10610 47268 10616
rect 47124 10124 47176 10130
rect 47124 10066 47176 10072
rect 47032 8968 47084 8974
rect 47032 8910 47084 8916
rect 46940 7880 46992 7886
rect 46940 7822 46992 7828
rect 46940 7472 46992 7478
rect 46940 7414 46992 7420
rect 46480 4752 46532 4758
rect 46480 4694 46532 4700
rect 46952 4622 46980 7414
rect 47136 7410 47164 10066
rect 47308 9988 47360 9994
rect 47308 9930 47360 9936
rect 47320 9625 47348 9930
rect 47306 9616 47362 9625
rect 47412 9586 47440 12310
rect 47964 12238 47992 12582
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49160 12306 49188 12407
rect 49148 12300 49200 12306
rect 49148 12242 49200 12248
rect 47952 12232 48004 12238
rect 47952 12174 48004 12180
rect 49146 12064 49202 12073
rect 47950 11996 48258 12005
rect 49146 11999 49202 12008
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 49160 11830 49188 11999
rect 49148 11824 49200 11830
rect 49148 11766 49200 11772
rect 49146 11656 49202 11665
rect 49146 11591 49202 11600
rect 49160 11218 49188 11591
rect 49238 11248 49294 11257
rect 49148 11212 49200 11218
rect 49238 11183 49294 11192
rect 49148 11154 49200 11160
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 49146 10840 49202 10849
rect 49146 10775 49202 10784
rect 49160 10130 49188 10775
rect 49252 10742 49280 11183
rect 49240 10736 49292 10742
rect 49240 10678 49292 10684
rect 49330 10432 49386 10441
rect 49330 10367 49386 10376
rect 49148 10124 49200 10130
rect 49148 10066 49200 10072
rect 49238 10024 49294 10033
rect 49238 9959 49294 9968
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47306 9551 47362 9560
rect 47400 9580 47452 9586
rect 47400 9522 47452 9528
rect 49146 9208 49202 9217
rect 49146 9143 49202 9152
rect 47584 8900 47636 8906
rect 47584 8842 47636 8848
rect 47124 7404 47176 7410
rect 47124 7346 47176 7352
rect 47032 6928 47084 6934
rect 47032 6870 47084 6876
rect 46940 4616 46992 4622
rect 46940 4558 46992 4564
rect 45836 4276 45888 4282
rect 45836 4218 45888 4224
rect 45652 3052 45704 3058
rect 45652 2994 45704 3000
rect 45848 2446 45876 4218
rect 47044 4146 47072 6870
rect 47596 6322 47624 8842
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 49160 8566 49188 9143
rect 49252 9042 49280 9959
rect 49344 9654 49372 10367
rect 49332 9648 49384 9654
rect 49332 9590 49384 9596
rect 49240 9036 49292 9042
rect 49240 8978 49292 8984
rect 49330 8800 49386 8809
rect 49330 8735 49386 8744
rect 47768 8560 47820 8566
rect 47768 8502 47820 8508
rect 49148 8560 49200 8566
rect 49148 8502 49200 8508
rect 47676 8356 47728 8362
rect 47676 8298 47728 8304
rect 47216 6316 47268 6322
rect 47216 6258 47268 6264
rect 47584 6316 47636 6322
rect 47584 6258 47636 6264
rect 47124 6180 47176 6186
rect 47124 6122 47176 6128
rect 47032 4140 47084 4146
rect 47032 4082 47084 4088
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 46676 1465 46704 4014
rect 47136 3534 47164 6122
rect 47228 4758 47256 6258
rect 47400 5908 47452 5914
rect 47400 5850 47452 5856
rect 47308 4820 47360 4826
rect 47308 4762 47360 4768
rect 47216 4752 47268 4758
rect 47216 4694 47268 4700
rect 47124 3528 47176 3534
rect 47124 3470 47176 3476
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46768 1873 46796 2926
rect 46860 2689 46888 2926
rect 46846 2680 46902 2689
rect 46846 2615 46902 2624
rect 47320 2446 47348 4762
rect 47412 3058 47440 5850
rect 47688 5710 47716 8298
rect 47780 6798 47808 8502
rect 49238 8392 49294 8401
rect 49238 8327 49294 8336
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49146 7576 49202 7585
rect 49146 7511 49202 7520
rect 47860 7268 47912 7274
rect 47860 7210 47912 7216
rect 47768 6792 47820 6798
rect 47768 6734 47820 6740
rect 47676 5704 47728 5710
rect 47676 5646 47728 5652
rect 47872 5234 47900 7210
rect 49160 6866 49188 7511
rect 49252 7478 49280 8327
rect 49344 7954 49372 8735
rect 49332 7948 49384 7954
rect 49332 7890 49384 7896
rect 49240 7472 49292 7478
rect 49240 7414 49292 7420
rect 49330 7168 49386 7177
rect 49330 7103 49386 7112
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 49238 6760 49294 6769
rect 48688 6724 48740 6730
rect 49238 6695 49294 6704
rect 48688 6666 48740 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48700 6361 48728 6666
rect 48686 6352 48742 6361
rect 48686 6287 48742 6296
rect 49146 5944 49202 5953
rect 49146 5879 49202 5888
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49160 5302 49188 5879
rect 49252 5778 49280 6695
rect 49344 6390 49372 7103
rect 49332 6384 49384 6390
rect 49332 6326 49384 6332
rect 49240 5772 49292 5778
rect 49240 5714 49292 5720
rect 49422 5536 49478 5545
rect 49422 5471 49478 5480
rect 49148 5296 49200 5302
rect 49148 5238 49200 5244
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 49330 5128 49386 5137
rect 48332 4729 48360 5102
rect 49330 5063 49386 5072
rect 48318 4720 48374 4729
rect 48318 4655 48374 4664
rect 47676 4548 47728 4554
rect 47676 4490 47728 4496
rect 47688 3942 47716 4490
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 47676 3936 47728 3942
rect 47676 3878 47728 3884
rect 47400 3052 47452 3058
rect 47400 2994 47452 3000
rect 47308 2440 47360 2446
rect 47308 2382 47360 2388
rect 46754 1864 46810 1873
rect 46754 1799 46810 1808
rect 46662 1456 46718 1465
rect 46662 1391 46718 1400
rect 47688 800 47716 3878
rect 49160 3602 49188 4247
rect 49344 4146 49372 5063
rect 49436 4690 49464 5471
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49792 4480 49844 4486
rect 49792 4422 49844 4428
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49238 3904 49294 3913
rect 49238 3839 49294 3848
rect 49148 3596 49200 3602
rect 49148 3538 49200 3544
rect 49146 3496 49202 3505
rect 48688 3460 48740 3466
rect 49146 3431 49202 3440
rect 48688 3402 48740 3408
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48700 3097 48728 3402
rect 48686 3088 48742 3097
rect 48686 3023 48742 3032
rect 49160 2514 49188 3431
rect 49252 3126 49280 3839
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 2281 48544 2314
rect 48502 2272 48558 2281
rect 47950 2204 48258 2213
rect 48502 2207 48558 2216
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49804 800 49832 4422
rect 28736 734 28948 762
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< via2 >>
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2778 24384 2834 24440
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 1766 21528 1822 21584
rect 1030 20712 1086 20768
rect 1306 20304 1362 20360
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 4066 25608 4122 25664
rect 3698 25200 3754 25256
rect 3606 24792 3662 24848
rect 3514 23976 3570 24032
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2778 21120 2834 21176
rect 1766 19896 1822 19952
rect 1490 18672 1546 18728
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2870 19488 2926 19544
rect 3514 21956 3570 21992
rect 3514 21936 3516 21956
rect 3516 21936 3568 21956
rect 3568 21936 3570 21956
rect 2778 19080 2834 19136
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3790 23160 3846 23216
rect 3974 23588 4030 23624
rect 3974 23568 3976 23588
rect 3976 23568 4028 23588
rect 4028 23568 4030 23588
rect 3974 22752 4030 22808
rect 1766 18264 1822 18320
rect 4158 22480 4214 22536
rect 1398 17856 1454 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 1766 17448 1822 17504
rect 1030 17040 1086 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 938 16632 994 16688
rect 1030 16224 1086 16280
rect 7470 24248 7526 24304
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 5262 19080 5318 19136
rect 1030 15816 1086 15872
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 938 15428 994 15464
rect 938 15408 940 15428
rect 940 15408 992 15428
rect 992 15408 994 15428
rect 938 15020 994 15056
rect 938 15000 940 15020
rect 940 15000 992 15020
rect 992 15000 994 15020
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 938 14592 994 14648
rect 1030 14184 1086 14240
rect 1766 13776 1822 13832
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3514 13368 3570 13424
rect 1306 12960 1362 13016
rect 1306 12552 1362 12608
rect 1214 12144 1270 12200
rect 1306 11756 1362 11792
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 1306 11736 1308 11756
rect 1308 11736 1360 11756
rect 1360 11736 1362 11756
rect 1306 11328 1362 11384
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 1306 10920 1362 10976
rect 1582 10512 1638 10568
rect 1214 10104 1270 10160
rect 1306 9696 1362 9752
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8390 20884 8392 20904
rect 8392 20884 8444 20904
rect 8444 20884 8446 20904
rect 8390 20848 8446 20884
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 11978 23160 12034 23216
rect 11334 23024 11390 23080
rect 11058 20340 11060 20360
rect 11060 20340 11112 20360
rect 11112 20340 11114 20360
rect 11058 20304 11114 20340
rect 10782 19796 10784 19816
rect 10784 19796 10836 19816
rect 10836 19796 10838 19816
rect 10782 19760 10838 19796
rect 10598 17720 10654 17776
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 11058 19216 11114 19272
rect 11610 21392 11666 21448
rect 11426 19896 11482 19952
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13542 22616 13598 22672
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 11794 20712 11850 20768
rect 11886 20304 11942 20360
rect 10506 15272 10562 15328
rect 11058 15952 11114 16008
rect 9954 14184 10010 14240
rect 10506 13812 10508 13832
rect 10508 13812 10560 13832
rect 10560 13812 10562 13832
rect 10506 13776 10562 13812
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 1306 9288 1362 9344
rect 3698 9460 3700 9480
rect 3700 9460 3752 9480
rect 3752 9460 3754 9480
rect 3698 9424 3754 9460
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 1582 8880 1638 8936
rect 1214 8472 1270 8528
rect 2410 8064 2466 8120
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 1306 7656 1362 7712
rect 1582 7248 1638 7304
rect 1306 6432 1362 6488
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3330 6840 3386 6896
rect 2870 6704 2926 6760
rect 1306 6024 1362 6080
rect 1306 5636 1362 5672
rect 1306 5616 1308 5636
rect 1308 5616 1360 5636
rect 1360 5616 1362 5636
rect 1398 5208 1454 5264
rect 1306 4800 1362 4856
rect 1306 4392 1362 4448
rect 1306 4020 1308 4040
rect 1308 4020 1360 4040
rect 1360 4020 1362 4040
rect 1306 3984 1362 4020
rect 1214 3576 1270 3632
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1306 3168 1362 3224
rect 1306 2760 1362 2816
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 1306 2372 1362 2408
rect 1306 2352 1308 2372
rect 1308 2352 1360 2372
rect 1360 2352 1362 2372
rect 1214 1944 1270 2000
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 11978 19080 12034 19136
rect 11610 16224 11666 16280
rect 11518 15408 11574 15464
rect 11242 14456 11298 14512
rect 11334 13096 11390 13152
rect 12438 20460 12494 20496
rect 12438 20440 12440 20460
rect 12440 20440 12492 20460
rect 12492 20440 12494 20460
rect 12346 18400 12402 18456
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12898 20984 12954 21040
rect 12714 20304 12770 20360
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 4066 1536 4122 1592
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12346 15544 12402 15600
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13818 20460 13874 20496
rect 13818 20440 13820 20460
rect 13820 20440 13872 20460
rect 13872 20440 13874 20460
rect 13634 20168 13690 20224
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12438 15272 12494 15328
rect 12346 15020 12402 15056
rect 12346 15000 12348 15020
rect 12348 15000 12400 15020
rect 12400 15000 12402 15020
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13266 15544 13322 15600
rect 13818 18264 13874 18320
rect 14278 17584 14334 17640
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12254 12688 12310 12744
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12898 12980 12954 13016
rect 12898 12960 12900 12980
rect 12900 12960 12952 12980
rect 12952 12960 12954 12980
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13358 12008 13414 12064
rect 14186 17196 14242 17232
rect 14186 17176 14188 17196
rect 14188 17176 14240 17196
rect 14240 17176 14242 17196
rect 15198 21528 15254 21584
rect 15658 19760 15714 19816
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 15198 19236 15254 19272
rect 15198 19216 15200 19236
rect 15200 19216 15252 19236
rect 15252 19216 15254 19236
rect 15658 18708 15660 18728
rect 15660 18708 15712 18728
rect 15712 18708 15714 18728
rect 15658 18672 15714 18708
rect 15934 19372 15990 19408
rect 15934 19352 15936 19372
rect 15936 19352 15988 19372
rect 15988 19352 15990 19372
rect 14002 14728 14058 14784
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13082 10104 13138 10160
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13450 10784 13506 10840
rect 13634 10668 13690 10704
rect 13634 10648 13636 10668
rect 13636 10648 13688 10668
rect 13688 10648 13690 10668
rect 14186 16088 14242 16144
rect 14646 15408 14702 15464
rect 14094 13368 14150 13424
rect 14002 13232 14058 13288
rect 14002 12552 14058 12608
rect 15106 16632 15162 16688
rect 14738 14900 14740 14920
rect 14740 14900 14792 14920
rect 14792 14900 14794 14920
rect 14738 14864 14794 14900
rect 14462 13368 14518 13424
rect 14370 13232 14426 13288
rect 14462 13096 14518 13152
rect 15014 13252 15070 13288
rect 15014 13232 15016 13252
rect 15016 13232 15068 13252
rect 15068 13232 15070 13252
rect 14922 12552 14978 12608
rect 14278 10512 14334 10568
rect 14370 8880 14426 8936
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 15198 12980 15254 13016
rect 15198 12960 15200 12980
rect 15200 12960 15252 12980
rect 15252 12960 15254 12980
rect 15842 16108 15898 16144
rect 15842 16088 15844 16108
rect 15844 16088 15896 16108
rect 15896 16088 15898 16108
rect 15750 15408 15806 15464
rect 16670 19760 16726 19816
rect 17222 19760 17278 19816
rect 16946 18672 17002 18728
rect 16302 13912 16358 13968
rect 16486 13640 16542 13696
rect 15934 10532 15990 10568
rect 15934 10512 15936 10532
rect 15936 10512 15988 10532
rect 15988 10512 15990 10532
rect 16670 15952 16726 16008
rect 17038 18284 17094 18320
rect 17038 18264 17040 18284
rect 17040 18264 17092 18284
rect 17092 18264 17094 18284
rect 17498 19352 17554 19408
rect 17406 18128 17462 18184
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17866 21936 17922 21992
rect 17590 17992 17646 18048
rect 17406 16244 17462 16280
rect 17406 16224 17408 16244
rect 17408 16224 17460 16244
rect 17460 16224 17462 16244
rect 16854 14220 16856 14240
rect 16856 14220 16908 14240
rect 16908 14220 16910 14240
rect 16854 14184 16910 14220
rect 16670 12688 16726 12744
rect 17130 13504 17186 13560
rect 17130 13252 17186 13288
rect 17130 13232 17132 13252
rect 17132 13232 17184 13252
rect 17184 13232 17186 13252
rect 17774 18400 17830 18456
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 19338 20712 19394 20768
rect 18694 19896 18750 19952
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17682 13232 17738 13288
rect 17222 12044 17224 12064
rect 17224 12044 17276 12064
rect 17276 12044 17278 12064
rect 17222 12008 17278 12044
rect 16486 9580 16542 9616
rect 16486 9560 16488 9580
rect 16488 9560 16540 9580
rect 16540 9560 16542 9580
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 15750 3984 15806 4040
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17498 10804 17554 10840
rect 17498 10784 17500 10804
rect 17500 10784 17552 10804
rect 17552 10784 17554 10804
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18602 16360 18658 16416
rect 18510 15544 18566 15600
rect 19338 19624 19394 19680
rect 19430 19252 19432 19272
rect 19432 19252 19484 19272
rect 19484 19252 19486 19272
rect 19430 19216 19486 19252
rect 18786 16360 18842 16416
rect 18786 15544 18842 15600
rect 18786 14592 18842 14648
rect 18050 13912 18106 13968
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17774 9560 17830 9616
rect 18602 14220 18604 14240
rect 18604 14220 18656 14240
rect 18656 14220 18658 14240
rect 18602 14184 18658 14220
rect 19154 15852 19156 15872
rect 19156 15852 19208 15872
rect 19208 15852 19210 15872
rect 19154 15816 19210 15852
rect 19430 17992 19486 18048
rect 22190 23160 22246 23216
rect 20350 20712 20406 20768
rect 19246 15156 19302 15192
rect 19246 15136 19248 15156
rect 19248 15136 19300 15156
rect 19300 15136 19302 15156
rect 18970 14884 19026 14920
rect 18970 14864 18972 14884
rect 18972 14864 19024 14884
rect 19024 14864 19026 14884
rect 19154 14728 19210 14784
rect 18510 12960 18566 13016
rect 18418 12824 18474 12880
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 20534 19216 20590 19272
rect 20626 18808 20682 18864
rect 22558 22072 22614 22128
rect 21822 20984 21878 21040
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 20626 14320 20682 14376
rect 20994 14456 21050 14512
rect 20994 13776 21050 13832
rect 20902 13232 20958 13288
rect 20994 12552 21050 12608
rect 22374 21664 22430 21720
rect 22374 21392 22430 21448
rect 22466 20984 22522 21040
rect 22190 20440 22246 20496
rect 21822 14320 21878 14376
rect 22466 20712 22522 20768
rect 22374 17176 22430 17232
rect 22374 17040 22430 17096
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23294 23024 23350 23080
rect 22834 22616 22890 22672
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23386 21392 23442 21448
rect 22742 20168 22798 20224
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23754 21800 23810 21856
rect 23938 22480 23994 22536
rect 23662 20848 23718 20904
rect 23386 19896 23442 19952
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 24122 21800 24178 21856
rect 25778 24284 25780 24304
rect 25780 24284 25832 24304
rect 25832 24284 25834 24304
rect 25778 24248 25834 24284
rect 24766 22616 24822 22672
rect 25318 22924 25320 22944
rect 25320 22924 25372 22944
rect 25372 22924 25374 22944
rect 25318 22888 25374 22924
rect 24766 22480 24822 22536
rect 24674 22208 24730 22264
rect 24582 21664 24638 21720
rect 23754 19488 23810 19544
rect 22742 15680 22798 15736
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 21546 9596 21548 9616
rect 21548 9596 21600 9616
rect 21600 9596 21602 9616
rect 21546 9560 21602 9596
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22374 12300 22430 12336
rect 22374 12280 22376 12300
rect 22376 12280 22428 12300
rect 22428 12280 22430 12300
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22834 12960 22890 13016
rect 22926 12724 22928 12744
rect 22928 12724 22980 12744
rect 22980 12724 22982 12744
rect 22926 12688 22982 12724
rect 22742 12552 22798 12608
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23570 12552 23626 12608
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 24582 18944 24638 19000
rect 24674 17584 24730 17640
rect 25226 21120 25282 21176
rect 25134 20712 25190 20768
rect 25226 20440 25282 20496
rect 25134 18284 25190 18320
rect 25134 18264 25136 18284
rect 25136 18264 25188 18284
rect 25188 18264 25190 18284
rect 25594 20712 25650 20768
rect 25870 21292 25872 21312
rect 25872 21292 25924 21312
rect 25924 21292 25926 21312
rect 25870 21256 25926 21292
rect 26606 24268 26662 24304
rect 26606 24248 26608 24268
rect 26608 24248 26660 24268
rect 26660 24248 26662 24268
rect 26422 22072 26478 22128
rect 26054 21428 26056 21448
rect 26056 21428 26108 21448
rect 26108 21428 26110 21448
rect 26054 21392 26110 21428
rect 26146 21120 26202 21176
rect 25962 20848 26018 20904
rect 23754 10104 23810 10160
rect 24582 13368 24638 13424
rect 24490 12552 24546 12608
rect 24858 14864 24914 14920
rect 26514 20884 26516 20904
rect 26516 20884 26568 20904
rect 26568 20884 26570 20904
rect 26514 20848 26570 20884
rect 26238 20712 26294 20768
rect 26054 19916 26110 19952
rect 26054 19896 26056 19916
rect 26056 19896 26108 19916
rect 26108 19896 26110 19916
rect 26146 19388 26148 19408
rect 26148 19388 26200 19408
rect 26200 19388 26202 19408
rect 26146 19352 26202 19388
rect 26146 18944 26202 19000
rect 25962 18264 26018 18320
rect 26330 17856 26386 17912
rect 26238 17620 26240 17640
rect 26240 17620 26292 17640
rect 26292 17620 26294 17640
rect 26238 17584 26294 17620
rect 26238 16904 26294 16960
rect 25686 15428 25742 15464
rect 25686 15408 25688 15428
rect 25688 15408 25740 15428
rect 25740 15408 25742 15428
rect 25226 12724 25228 12744
rect 25228 12724 25280 12744
rect 25280 12724 25282 12744
rect 25226 12688 25282 12724
rect 26330 15000 26386 15056
rect 26606 17720 26662 17776
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27066 21120 27122 21176
rect 27342 20868 27398 20904
rect 27342 20848 27344 20868
rect 27344 20848 27396 20868
rect 27396 20848 27398 20868
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27158 19660 27160 19680
rect 27160 19660 27212 19680
rect 27212 19660 27214 19680
rect 27158 19624 27214 19660
rect 26974 17076 26976 17096
rect 26976 17076 27028 17096
rect 27028 17076 27030 17096
rect 26974 17040 27030 17076
rect 27066 16088 27122 16144
rect 26790 12960 26846 13016
rect 27066 15544 27122 15600
rect 27158 12960 27214 13016
rect 27434 18944 27490 19000
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 28354 19372 28410 19408
rect 28354 19352 28356 19372
rect 28356 19352 28408 19372
rect 28408 19352 28410 19372
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 28354 18128 28410 18184
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27618 17196 27674 17232
rect 27618 17176 27620 17196
rect 27620 17176 27672 17196
rect 27672 17176 27674 17196
rect 28170 17176 28226 17232
rect 27342 15020 27398 15056
rect 27342 15000 27344 15020
rect 27344 15000 27396 15020
rect 27396 15000 27398 15020
rect 27986 17040 28042 17096
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 28814 20984 28870 21040
rect 28630 19488 28686 19544
rect 29182 19216 29238 19272
rect 28998 18672 29054 18728
rect 29182 18808 29238 18864
rect 29090 18536 29146 18592
rect 29366 21800 29422 21856
rect 29734 22208 29790 22264
rect 29550 21936 29606 21992
rect 29918 22072 29974 22128
rect 29734 21140 29790 21176
rect 29734 21120 29736 21140
rect 29736 21120 29788 21140
rect 29788 21120 29790 21140
rect 29550 19896 29606 19952
rect 29550 19292 29606 19348
rect 29734 19292 29790 19348
rect 30102 19796 30104 19816
rect 30104 19796 30156 19816
rect 30156 19796 30158 19816
rect 30102 19760 30158 19796
rect 30654 22480 30710 22536
rect 30562 20848 30618 20904
rect 30378 19780 30434 19816
rect 30378 19760 30380 19780
rect 30380 19760 30432 19780
rect 30432 19760 30434 19780
rect 30010 19250 30066 19306
rect 28906 17856 28962 17912
rect 28814 16904 28870 16960
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 25962 8916 25964 8936
rect 25964 8916 26016 8936
rect 26016 8916 26018 8936
rect 25962 8880 26018 8916
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27710 10104 27766 10160
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 28538 13132 28540 13152
rect 28540 13132 28592 13152
rect 28592 13132 28594 13152
rect 28538 13096 28594 13132
rect 29550 19080 29606 19136
rect 29642 18944 29698 19000
rect 29642 18672 29698 18728
rect 29366 15952 29422 16008
rect 28630 12688 28686 12744
rect 28814 13096 28870 13152
rect 30194 19080 30250 19136
rect 30102 17448 30158 17504
rect 30194 16632 30250 16688
rect 32494 24656 32550 24712
rect 31482 22616 31538 22672
rect 31206 21956 31262 21992
rect 31206 21936 31208 21956
rect 31208 21936 31260 21956
rect 31260 21936 31262 21956
rect 31206 21684 31262 21720
rect 31206 21664 31208 21684
rect 31208 21664 31260 21684
rect 31260 21664 31262 21684
rect 31390 20848 31446 20904
rect 30746 18944 30802 19000
rect 30746 18808 30802 18864
rect 29734 11736 29790 11792
rect 28630 10104 28686 10160
rect 31022 20440 31078 20496
rect 30930 18400 30986 18456
rect 31850 21936 31906 21992
rect 31666 20476 31668 20496
rect 31668 20476 31720 20496
rect 31720 20476 31722 20496
rect 31666 20440 31722 20476
rect 31114 17584 31170 17640
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33598 23432 33654 23488
rect 33414 23296 33470 23352
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 31942 20340 31944 20360
rect 31944 20340 31996 20360
rect 31996 20340 31998 20360
rect 31942 20304 31998 20340
rect 32862 21800 32918 21856
rect 33230 21800 33286 21856
rect 33230 21528 33286 21584
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32862 20984 32918 21040
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 34058 23568 34114 23624
rect 33690 22344 33746 22400
rect 33598 21684 33654 21720
rect 33598 21664 33600 21684
rect 33600 21664 33652 21684
rect 33652 21664 33654 21684
rect 33506 21548 33562 21584
rect 33506 21528 33508 21548
rect 33508 21528 33560 21548
rect 33560 21528 33562 21548
rect 30102 12280 30158 12336
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27894 4020 27896 4040
rect 27896 4020 27948 4040
rect 27948 4020 27950 4040
rect 27894 3984 27950 4020
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 30562 12824 30618 12880
rect 30470 11600 30526 11656
rect 30746 10512 30802 10568
rect 30930 9016 30986 9072
rect 31758 9696 31814 9752
rect 32770 19216 32826 19272
rect 32586 18536 32642 18592
rect 32770 18672 32826 18728
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 33138 18536 33194 18592
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 34242 23160 34298 23216
rect 35254 23704 35310 23760
rect 34610 22924 34612 22944
rect 34612 22924 34664 22944
rect 34664 22924 34666 22944
rect 34610 22888 34666 22924
rect 34794 22480 34850 22536
rect 34426 21664 34482 21720
rect 33782 19488 33838 19544
rect 33598 18944 33654 19000
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32310 9716 32366 9752
rect 32310 9696 32312 9716
rect 32312 9696 32364 9716
rect 32364 9696 32366 9716
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 33874 18572 33876 18592
rect 33876 18572 33928 18592
rect 33928 18572 33930 18592
rect 33874 18536 33930 18572
rect 33874 17584 33930 17640
rect 33690 16224 33746 16280
rect 34150 18828 34206 18864
rect 34150 18808 34152 18828
rect 34152 18808 34204 18828
rect 34204 18808 34206 18828
rect 35346 22344 35402 22400
rect 35254 21836 35256 21856
rect 35256 21836 35308 21856
rect 35308 21836 35310 21856
rect 35254 21800 35310 21836
rect 34610 20440 34666 20496
rect 33506 9424 33562 9480
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 34794 19080 34850 19136
rect 34886 15544 34942 15600
rect 35254 20712 35310 20768
rect 36082 23432 36138 23488
rect 35898 23024 35954 23080
rect 35990 22888 36046 22944
rect 35806 22616 35862 22672
rect 36082 22072 36138 22128
rect 35530 17584 35586 17640
rect 35714 17584 35770 17640
rect 35438 17484 35440 17504
rect 35440 17484 35492 17504
rect 35492 17484 35494 17504
rect 35438 17448 35494 17484
rect 35162 12824 35218 12880
rect 35714 16088 35770 16144
rect 35714 15952 35770 16008
rect 36082 18944 36138 19000
rect 37002 22888 37058 22944
rect 37370 23432 37426 23488
rect 37278 22480 37334 22536
rect 37278 22072 37334 22128
rect 36910 19116 36912 19136
rect 36912 19116 36964 19136
rect 36964 19116 36966 19136
rect 35714 14456 35770 14512
rect 35622 11600 35678 11656
rect 36910 19080 36966 19116
rect 36358 16224 36414 16280
rect 36634 16632 36690 16688
rect 36450 12824 36506 12880
rect 37278 21800 37334 21856
rect 37370 21664 37426 21720
rect 37186 21428 37188 21448
rect 37188 21428 37240 21448
rect 37240 21428 37242 21448
rect 37186 21392 37242 21428
rect 37554 21120 37610 21176
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37830 23704 37886 23760
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37278 20748 37280 20768
rect 37280 20748 37332 20768
rect 37332 20748 37334 20768
rect 37278 20712 37334 20748
rect 37094 18944 37150 19000
rect 37094 18128 37150 18184
rect 37186 14456 37242 14512
rect 35990 9052 35992 9072
rect 35992 9052 36044 9072
rect 36044 9052 36046 9072
rect 35990 9016 36046 9052
rect 36542 10532 36598 10568
rect 36542 10512 36544 10532
rect 36544 10512 36596 10532
rect 36596 10512 36598 10532
rect 38566 21800 38622 21856
rect 38382 20848 38438 20904
rect 39302 23704 39358 23760
rect 39394 23024 39450 23080
rect 39946 23568 40002 23624
rect 39486 21936 39542 21992
rect 40038 21256 40094 21312
rect 38474 20712 38530 20768
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37646 19080 37702 19136
rect 38014 18672 38070 18728
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 43534 24656 43590 24712
rect 40682 23160 40738 23216
rect 40314 22380 40316 22400
rect 40316 22380 40368 22400
rect 40368 22380 40370 22400
rect 40314 22344 40370 22380
rect 40314 21120 40370 21176
rect 40038 20712 40094 20768
rect 39762 19760 39818 19816
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 38290 16496 38346 16552
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 40590 21836 40592 21856
rect 40592 21836 40644 21856
rect 40644 21836 40646 21856
rect 40590 21800 40646 21836
rect 41050 20712 41106 20768
rect 40590 19372 40646 19408
rect 40590 19352 40592 19372
rect 40592 19352 40644 19372
rect 40644 19352 40646 19372
rect 40406 17992 40462 18048
rect 41418 22752 41474 22808
rect 42522 23860 42578 23896
rect 42522 23840 42524 23860
rect 42524 23840 42576 23860
rect 42576 23840 42578 23860
rect 42430 23024 42486 23080
rect 42982 23840 43038 23896
rect 42798 23432 42854 23488
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 43350 23160 43406 23216
rect 42798 22616 42854 22672
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 41418 20848 41474 20904
rect 41326 18944 41382 19000
rect 42614 21528 42670 21584
rect 41234 18128 41290 18184
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 40222 16632 40278 16688
rect 39946 16496 40002 16552
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 43810 22480 43866 22536
rect 43994 24248 44050 24304
rect 43994 19896 44050 19952
rect 46202 25064 46258 25120
rect 45742 22752 45798 22808
rect 45190 22092 45246 22128
rect 45190 22072 45192 22092
rect 45192 22072 45244 22092
rect 45244 22072 45246 22092
rect 45190 21392 45246 21448
rect 45466 20984 45522 21040
rect 46570 24656 46626 24712
rect 46478 23704 46534 23760
rect 46294 20440 46350 20496
rect 46846 25472 46902 25528
rect 46846 23432 46902 23488
rect 46570 20304 46626 20360
rect 44270 19216 44326 19272
rect 47398 20748 47400 20768
rect 47400 20748 47452 20768
rect 47452 20748 47454 20768
rect 47398 20712 47454 20748
rect 47766 23024 47822 23080
rect 47674 21528 47730 21584
rect 48042 24112 48098 24168
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 48042 23024 48098 23080
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 48410 20168 48466 20224
rect 47306 18808 47362 18864
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 48410 18536 48466 18592
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47674 18128 47730 18184
rect 46938 17756 46940 17776
rect 46940 17756 46992 17776
rect 46992 17756 46994 17776
rect 46938 17720 46994 17756
rect 48042 17584 48098 17640
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 41878 17176 41934 17232
rect 47950 17076 47952 17096
rect 47952 17076 48004 17096
rect 48004 17076 48006 17096
rect 47950 17040 48006 17076
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 48318 16940 48320 16960
rect 48320 16940 48372 16960
rect 48372 16940 48374 16960
rect 48318 16904 48374 16940
rect 49514 24248 49570 24304
rect 49330 22616 49386 22672
rect 49238 22208 49294 22264
rect 49330 21392 49386 21448
rect 49238 20984 49294 21040
rect 49330 20576 49386 20632
rect 49330 19760 49386 19816
rect 49422 19352 49478 19408
rect 49330 18944 49386 19000
rect 49422 18128 49478 18184
rect 49330 17720 49386 17776
rect 49330 17312 49386 17368
rect 48226 16496 48282 16552
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 49330 16088 49386 16144
rect 49146 15952 49202 16008
rect 48686 15680 48742 15736
rect 47858 15408 47914 15464
rect 48594 15272 48650 15328
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47858 15000 47914 15056
rect 39302 14456 39358 14512
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 40038 12688 40094 12744
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 48042 14884 48098 14920
rect 48042 14864 48044 14884
rect 48044 14864 48096 14884
rect 48096 14864 48098 14884
rect 49330 14864 49386 14920
rect 49330 14456 49386 14512
rect 47950 14356 47952 14376
rect 47952 14356 48004 14376
rect 48004 14356 48006 14376
rect 47950 14320 48006 14356
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 49330 14048 49386 14104
rect 47674 13640 47730 13696
rect 49146 13268 49148 13288
rect 49148 13268 49200 13288
rect 49200 13268 49202 13288
rect 49146 13232 49202 13268
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 49146 12844 49202 12880
rect 49146 12824 49148 12844
rect 49148 12824 49200 12844
rect 49200 12824 49202 12844
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 40406 11772 40408 11792
rect 40408 11772 40460 11792
rect 40460 11772 40462 11792
rect 40406 11736 40462 11772
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 46846 7928 46902 7984
rect 47306 9560 47362 9616
rect 49146 12416 49202 12472
rect 49146 12008 49202 12064
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 49146 11600 49202 11656
rect 49238 11192 49294 11248
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49146 10784 49202 10840
rect 49330 10376 49386 10432
rect 49238 9968 49294 10024
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 49146 9152 49202 9208
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 49330 8744 49386 8800
rect 46846 2624 46902 2680
rect 49238 8336 49294 8392
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7520 49202 7576
rect 49330 7112 49386 7168
rect 49238 6704 49294 6760
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 48686 6296 48742 6352
rect 49146 5888 49202 5944
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 49422 5480 49478 5536
rect 49330 5072 49386 5128
rect 48318 4664 48374 4720
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 4256 49202 4312
rect 46754 1808 46810 1864
rect 46662 1400 46718 1456
rect 49238 3848 49294 3904
rect 49146 3440 49202 3496
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 48686 3032 48742 3088
rect 48502 2216 48558 2272
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 4061 25666 4127 25669
rect 0 25664 4127 25666
rect 0 25608 4066 25664
rect 4122 25608 4127 25664
rect 0 25606 4127 25608
rect 0 25576 800 25606
rect 4061 25603 4127 25606
rect 46841 25530 46907 25533
rect 50200 25530 51000 25560
rect 46841 25528 51000 25530
rect 46841 25472 46846 25528
rect 46902 25472 51000 25528
rect 46841 25470 51000 25472
rect 46841 25467 46907 25470
rect 50200 25440 51000 25470
rect 0 25258 800 25288
rect 3693 25258 3759 25261
rect 0 25256 3759 25258
rect 0 25200 3698 25256
rect 3754 25200 3759 25256
rect 0 25198 3759 25200
rect 0 25168 800 25198
rect 3693 25195 3759 25198
rect 46197 25122 46263 25125
rect 50200 25122 51000 25152
rect 46197 25120 51000 25122
rect 46197 25064 46202 25120
rect 46258 25064 51000 25120
rect 46197 25062 51000 25064
rect 46197 25059 46263 25062
rect 50200 25032 51000 25062
rect 0 24850 800 24880
rect 3601 24850 3667 24853
rect 0 24848 3667 24850
rect 0 24792 3606 24848
rect 3662 24792 3667 24848
rect 0 24790 3667 24792
rect 0 24760 800 24790
rect 3601 24787 3667 24790
rect 32489 24714 32555 24717
rect 43529 24714 43595 24717
rect 32489 24712 43595 24714
rect 32489 24656 32494 24712
rect 32550 24656 43534 24712
rect 43590 24656 43595 24712
rect 32489 24654 43595 24656
rect 32489 24651 32555 24654
rect 43529 24651 43595 24654
rect 46565 24714 46631 24717
rect 50200 24714 51000 24744
rect 46565 24712 51000 24714
rect 46565 24656 46570 24712
rect 46626 24656 51000 24712
rect 46565 24654 51000 24656
rect 46565 24651 46631 24654
rect 50200 24624 51000 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 7465 24306 7531 24309
rect 25773 24306 25839 24309
rect 7465 24304 25839 24306
rect 7465 24248 7470 24304
rect 7526 24248 25778 24304
rect 25834 24248 25839 24304
rect 7465 24246 25839 24248
rect 7465 24243 7531 24246
rect 25773 24243 25839 24246
rect 26601 24306 26667 24309
rect 43989 24306 44055 24309
rect 26601 24304 44055 24306
rect 26601 24248 26606 24304
rect 26662 24248 43994 24304
rect 44050 24248 44055 24304
rect 26601 24246 44055 24248
rect 26601 24243 26667 24246
rect 43989 24243 44055 24246
rect 49509 24306 49575 24309
rect 50200 24306 51000 24336
rect 49509 24304 51000 24306
rect 49509 24248 49514 24304
rect 49570 24248 51000 24304
rect 49509 24246 51000 24248
rect 49509 24243 49575 24246
rect 50200 24216 51000 24246
rect 28574 24108 28580 24172
rect 28644 24170 28650 24172
rect 48037 24170 48103 24173
rect 28644 24168 48103 24170
rect 28644 24112 48042 24168
rect 48098 24112 48103 24168
rect 28644 24110 48103 24112
rect 28644 24108 28650 24110
rect 48037 24107 48103 24110
rect 0 24034 800 24064
rect 3509 24034 3575 24037
rect 0 24032 3575 24034
rect 0 23976 3514 24032
rect 3570 23976 3575 24032
rect 0 23974 3575 23976
rect 0 23944 800 23974
rect 3509 23971 3575 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 42517 23898 42583 23901
rect 42977 23898 43043 23901
rect 50200 23898 51000 23928
rect 42517 23896 43043 23898
rect 42517 23840 42522 23896
rect 42578 23840 42982 23896
rect 43038 23840 43043 23896
rect 42517 23838 43043 23840
rect 42517 23835 42583 23838
rect 42977 23835 43043 23838
rect 48454 23838 51000 23898
rect 28942 23700 28948 23764
rect 29012 23762 29018 23764
rect 35249 23762 35315 23765
rect 37825 23762 37891 23765
rect 39297 23762 39363 23765
rect 29012 23760 39363 23762
rect 29012 23704 35254 23760
rect 35310 23704 37830 23760
rect 37886 23704 39302 23760
rect 39358 23704 39363 23760
rect 29012 23702 39363 23704
rect 29012 23700 29018 23702
rect 35249 23699 35315 23702
rect 37825 23699 37891 23702
rect 39297 23699 39363 23702
rect 46473 23762 46539 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 46473 23760 48514 23762
rect 46473 23704 46478 23760
rect 46534 23704 48514 23760
rect 46473 23702 48514 23704
rect 46473 23699 46539 23702
rect 0 23626 800 23656
rect 3969 23626 4035 23629
rect 0 23624 4035 23626
rect 0 23568 3974 23624
rect 4030 23568 4035 23624
rect 0 23566 4035 23568
rect 0 23536 800 23566
rect 3969 23563 4035 23566
rect 34053 23626 34119 23629
rect 39941 23626 40007 23629
rect 34053 23624 40007 23626
rect 34053 23568 34058 23624
rect 34114 23568 39946 23624
rect 40002 23568 40007 23624
rect 34053 23566 40007 23568
rect 34053 23563 34119 23566
rect 39941 23563 40007 23566
rect 33593 23490 33659 23493
rect 36077 23490 36143 23493
rect 33593 23488 36143 23490
rect 33593 23432 33598 23488
rect 33654 23432 36082 23488
rect 36138 23432 36143 23488
rect 33593 23430 36143 23432
rect 33593 23427 33659 23430
rect 36077 23427 36143 23430
rect 37365 23490 37431 23493
rect 42793 23490 42859 23493
rect 37365 23488 42859 23490
rect 37365 23432 37370 23488
rect 37426 23432 42798 23488
rect 42854 23432 42859 23488
rect 37365 23430 42859 23432
rect 37365 23427 37431 23430
rect 42793 23427 42859 23430
rect 46841 23490 46907 23493
rect 50200 23490 51000 23520
rect 46841 23488 51000 23490
rect 46841 23432 46846 23488
rect 46902 23432 51000 23488
rect 46841 23430 51000 23432
rect 46841 23427 46907 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 50200 23400 51000 23430
rect 42946 23359 43262 23360
rect 33409 23354 33475 23357
rect 33409 23352 41430 23354
rect 33409 23296 33414 23352
rect 33470 23296 41430 23352
rect 33409 23294 41430 23296
rect 33409 23291 33475 23294
rect 0 23218 800 23248
rect 3785 23218 3851 23221
rect 0 23216 3851 23218
rect 0 23160 3790 23216
rect 3846 23160 3851 23216
rect 0 23158 3851 23160
rect 0 23128 800 23158
rect 3785 23155 3851 23158
rect 11973 23218 12039 23221
rect 22185 23218 22251 23221
rect 11973 23216 22251 23218
rect 11973 23160 11978 23216
rect 12034 23160 22190 23216
rect 22246 23160 22251 23216
rect 11973 23158 22251 23160
rect 11973 23155 12039 23158
rect 22185 23155 22251 23158
rect 34237 23218 34303 23221
rect 40677 23218 40743 23221
rect 34237 23216 40743 23218
rect 34237 23160 34242 23216
rect 34298 23160 40682 23216
rect 40738 23160 40743 23216
rect 34237 23158 40743 23160
rect 41370 23218 41430 23294
rect 43345 23218 43411 23221
rect 41370 23216 43411 23218
rect 41370 23160 43350 23216
rect 43406 23160 43411 23216
rect 41370 23158 43411 23160
rect 34237 23155 34303 23158
rect 40677 23155 40743 23158
rect 43345 23155 43411 23158
rect 11329 23082 11395 23085
rect 23289 23082 23355 23085
rect 11329 23080 23355 23082
rect 11329 23024 11334 23080
rect 11390 23024 23294 23080
rect 23350 23024 23355 23080
rect 11329 23022 23355 23024
rect 11329 23019 11395 23022
rect 23289 23019 23355 23022
rect 35893 23082 35959 23085
rect 39389 23082 39455 23085
rect 35893 23080 39455 23082
rect 35893 23024 35898 23080
rect 35954 23024 39394 23080
rect 39450 23024 39455 23080
rect 35893 23022 39455 23024
rect 35893 23019 35959 23022
rect 39389 23019 39455 23022
rect 42425 23082 42491 23085
rect 47761 23082 47827 23085
rect 42425 23080 47827 23082
rect 42425 23024 42430 23080
rect 42486 23024 47766 23080
rect 47822 23024 47827 23080
rect 42425 23022 47827 23024
rect 42425 23019 42491 23022
rect 47761 23019 47827 23022
rect 48037 23082 48103 23085
rect 50200 23082 51000 23112
rect 48037 23080 51000 23082
rect 48037 23024 48042 23080
rect 48098 23024 51000 23080
rect 48037 23022 51000 23024
rect 48037 23019 48103 23022
rect 50200 22992 51000 23022
rect 25313 22948 25379 22949
rect 25262 22884 25268 22948
rect 25332 22946 25379 22948
rect 34605 22946 34671 22949
rect 35985 22946 36051 22949
rect 36997 22946 37063 22949
rect 25332 22944 25424 22946
rect 25374 22888 25424 22944
rect 25332 22886 25424 22888
rect 34605 22944 37063 22946
rect 34605 22888 34610 22944
rect 34666 22888 35990 22944
rect 36046 22888 37002 22944
rect 37058 22888 37063 22944
rect 34605 22886 37063 22888
rect 25332 22884 25379 22886
rect 25313 22883 25379 22884
rect 34605 22883 34671 22886
rect 35985 22883 36051 22886
rect 36997 22883 37063 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 3969 22810 4035 22813
rect 0 22808 4035 22810
rect 0 22752 3974 22808
rect 4030 22752 4035 22808
rect 0 22750 4035 22752
rect 0 22720 800 22750
rect 3969 22747 4035 22750
rect 41413 22810 41479 22813
rect 45737 22810 45803 22813
rect 41413 22808 45803 22810
rect 41413 22752 41418 22808
rect 41474 22752 45742 22808
rect 45798 22752 45803 22808
rect 41413 22750 45803 22752
rect 41413 22747 41479 22750
rect 45737 22747 45803 22750
rect 13537 22674 13603 22677
rect 22829 22674 22895 22677
rect 13537 22672 22895 22674
rect 13537 22616 13542 22672
rect 13598 22616 22834 22672
rect 22890 22616 22895 22672
rect 13537 22614 22895 22616
rect 13537 22611 13603 22614
rect 22829 22611 22895 22614
rect 24761 22674 24827 22677
rect 31477 22674 31543 22677
rect 24761 22672 31543 22674
rect 24761 22616 24766 22672
rect 24822 22616 31482 22672
rect 31538 22616 31543 22672
rect 24761 22614 31543 22616
rect 24761 22611 24827 22614
rect 31477 22611 31543 22614
rect 35801 22674 35867 22677
rect 42793 22674 42859 22677
rect 35801 22672 42859 22674
rect 35801 22616 35806 22672
rect 35862 22616 42798 22672
rect 42854 22616 42859 22672
rect 35801 22614 42859 22616
rect 35801 22611 35867 22614
rect 42793 22611 42859 22614
rect 49325 22674 49391 22677
rect 50200 22674 51000 22704
rect 49325 22672 51000 22674
rect 49325 22616 49330 22672
rect 49386 22616 51000 22672
rect 49325 22614 51000 22616
rect 49325 22611 49391 22614
rect 50200 22584 51000 22614
rect 4153 22538 4219 22541
rect 2086 22536 4219 22538
rect 2086 22480 4158 22536
rect 4214 22480 4219 22536
rect 2086 22478 4219 22480
rect 0 22402 800 22432
rect 2086 22402 2146 22478
rect 4153 22475 4219 22478
rect 23933 22538 23999 22541
rect 24761 22538 24827 22541
rect 23933 22536 24827 22538
rect 23933 22480 23938 22536
rect 23994 22480 24766 22536
rect 24822 22480 24827 22536
rect 23933 22478 24827 22480
rect 23933 22475 23999 22478
rect 24761 22475 24827 22478
rect 30649 22538 30715 22541
rect 34789 22538 34855 22541
rect 30649 22536 34855 22538
rect 30649 22480 30654 22536
rect 30710 22480 34794 22536
rect 34850 22480 34855 22536
rect 30649 22478 34855 22480
rect 30649 22475 30715 22478
rect 34789 22475 34855 22478
rect 37273 22538 37339 22541
rect 43805 22538 43871 22541
rect 37273 22536 43871 22538
rect 37273 22480 37278 22536
rect 37334 22480 43810 22536
rect 43866 22480 43871 22536
rect 37273 22478 43871 22480
rect 37273 22475 37339 22478
rect 43805 22475 43871 22478
rect 0 22342 2146 22402
rect 33685 22402 33751 22405
rect 35341 22402 35407 22405
rect 40309 22402 40375 22405
rect 33685 22400 40375 22402
rect 33685 22344 33690 22400
rect 33746 22344 35346 22400
rect 35402 22344 40314 22400
rect 40370 22344 40375 22400
rect 33685 22342 40375 22344
rect 0 22312 800 22342
rect 33685 22339 33751 22342
rect 35341 22339 35407 22342
rect 40309 22339 40375 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 24669 22266 24735 22269
rect 29729 22266 29795 22269
rect 24669 22264 29795 22266
rect 24669 22208 24674 22264
rect 24730 22208 29734 22264
rect 29790 22208 29795 22264
rect 24669 22206 29795 22208
rect 24669 22203 24735 22206
rect 29729 22203 29795 22206
rect 49233 22266 49299 22269
rect 50200 22266 51000 22296
rect 49233 22264 51000 22266
rect 49233 22208 49238 22264
rect 49294 22208 51000 22264
rect 49233 22206 51000 22208
rect 49233 22203 49299 22206
rect 50200 22176 51000 22206
rect 22553 22130 22619 22133
rect 26417 22130 26483 22133
rect 22553 22128 26483 22130
rect 22553 22072 22558 22128
rect 22614 22072 26422 22128
rect 26478 22072 26483 22128
rect 22553 22070 26483 22072
rect 22553 22067 22619 22070
rect 26417 22067 26483 22070
rect 29913 22130 29979 22133
rect 36077 22130 36143 22133
rect 29913 22128 36143 22130
rect 29913 22072 29918 22128
rect 29974 22072 36082 22128
rect 36138 22072 36143 22128
rect 29913 22070 36143 22072
rect 29913 22067 29979 22070
rect 36077 22067 36143 22070
rect 37273 22130 37339 22133
rect 45185 22130 45251 22133
rect 37273 22128 45251 22130
rect 37273 22072 37278 22128
rect 37334 22072 45190 22128
rect 45246 22072 45251 22128
rect 37273 22070 45251 22072
rect 37273 22067 37339 22070
rect 45185 22067 45251 22070
rect 0 21994 800 22024
rect 3509 21994 3575 21997
rect 0 21992 3575 21994
rect 0 21936 3514 21992
rect 3570 21936 3575 21992
rect 0 21934 3575 21936
rect 0 21904 800 21934
rect 3509 21931 3575 21934
rect 17861 21994 17927 21997
rect 29545 21994 29611 21997
rect 31201 21994 31267 21997
rect 17861 21992 26986 21994
rect 17861 21936 17866 21992
rect 17922 21936 26986 21992
rect 17861 21934 26986 21936
rect 17861 21931 17927 21934
rect 23749 21858 23815 21861
rect 24117 21858 24183 21861
rect 23749 21856 24183 21858
rect 23749 21800 23754 21856
rect 23810 21800 24122 21856
rect 24178 21800 24183 21856
rect 23749 21798 24183 21800
rect 23749 21795 23815 21798
rect 24117 21795 24183 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 22369 21722 22435 21725
rect 24577 21722 24643 21725
rect 22369 21720 24643 21722
rect 22369 21664 22374 21720
rect 22430 21664 24582 21720
rect 24638 21664 24643 21720
rect 22369 21662 24643 21664
rect 22369 21659 22435 21662
rect 24577 21659 24643 21662
rect 0 21586 800 21616
rect 1761 21586 1827 21589
rect 0 21584 1827 21586
rect 0 21528 1766 21584
rect 1822 21528 1827 21584
rect 0 21526 1827 21528
rect 0 21496 800 21526
rect 1761 21523 1827 21526
rect 15193 21586 15259 21589
rect 26926 21586 26986 21934
rect 29545 21992 31267 21994
rect 29545 21936 29550 21992
rect 29606 21936 31206 21992
rect 31262 21936 31267 21992
rect 29545 21934 31267 21936
rect 29545 21931 29611 21934
rect 31201 21931 31267 21934
rect 31845 21994 31911 21997
rect 39481 21994 39547 21997
rect 31845 21992 39547 21994
rect 31845 21936 31850 21992
rect 31906 21936 39486 21992
rect 39542 21936 39547 21992
rect 31845 21934 39547 21936
rect 31845 21931 31911 21934
rect 39481 21931 39547 21934
rect 29361 21858 29427 21861
rect 32857 21858 32923 21861
rect 29361 21856 32923 21858
rect 29361 21800 29366 21856
rect 29422 21800 32862 21856
rect 32918 21800 32923 21856
rect 29361 21798 32923 21800
rect 29361 21795 29427 21798
rect 32857 21795 32923 21798
rect 33225 21858 33291 21861
rect 35249 21858 35315 21861
rect 37273 21858 37339 21861
rect 33225 21856 37339 21858
rect 33225 21800 33230 21856
rect 33286 21800 35254 21856
rect 35310 21800 37278 21856
rect 37334 21800 37339 21856
rect 33225 21798 37339 21800
rect 33225 21795 33291 21798
rect 35249 21795 35315 21798
rect 37273 21795 37339 21798
rect 38561 21858 38627 21861
rect 40585 21858 40651 21861
rect 50200 21858 51000 21888
rect 38561 21856 40651 21858
rect 38561 21800 38566 21856
rect 38622 21800 40590 21856
rect 40646 21800 40651 21856
rect 38561 21798 40651 21800
rect 38561 21795 38627 21798
rect 40585 21795 40651 21798
rect 48454 21798 51000 21858
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 31201 21722 31267 21725
rect 33593 21722 33659 21725
rect 31201 21720 33659 21722
rect 31201 21664 31206 21720
rect 31262 21664 33598 21720
rect 33654 21664 33659 21720
rect 31201 21662 33659 21664
rect 31201 21659 31267 21662
rect 33593 21659 33659 21662
rect 34421 21722 34487 21725
rect 37365 21722 37431 21725
rect 34421 21720 37431 21722
rect 34421 21664 34426 21720
rect 34482 21664 37370 21720
rect 37426 21664 37431 21720
rect 34421 21662 37431 21664
rect 34421 21659 34487 21662
rect 37365 21659 37431 21662
rect 33225 21586 33291 21589
rect 15193 21584 22754 21586
rect 15193 21528 15198 21584
rect 15254 21528 22754 21584
rect 15193 21526 22754 21528
rect 26926 21584 33291 21586
rect 26926 21528 33230 21584
rect 33286 21528 33291 21584
rect 26926 21526 33291 21528
rect 15193 21523 15259 21526
rect 11605 21450 11671 21453
rect 22369 21450 22435 21453
rect 11605 21448 22435 21450
rect 11605 21392 11610 21448
rect 11666 21392 22374 21448
rect 22430 21392 22435 21448
rect 11605 21390 22435 21392
rect 11605 21387 11671 21390
rect 22369 21387 22435 21390
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 12893 21042 12959 21045
rect 21817 21042 21883 21045
rect 22461 21042 22527 21045
rect 12893 21040 22527 21042
rect 12893 20984 12898 21040
rect 12954 20984 21822 21040
rect 21878 20984 22466 21040
rect 22522 20984 22527 21040
rect 12893 20982 22527 20984
rect 22694 21042 22754 21526
rect 33225 21523 33291 21526
rect 33501 21586 33567 21589
rect 42609 21586 42675 21589
rect 33501 21584 42675 21586
rect 33501 21528 33506 21584
rect 33562 21528 42614 21584
rect 42670 21528 42675 21584
rect 33501 21526 42675 21528
rect 33501 21523 33567 21526
rect 42609 21523 42675 21526
rect 47669 21586 47735 21589
rect 48454 21586 48514 21798
rect 50200 21768 51000 21798
rect 47669 21584 48514 21586
rect 47669 21528 47674 21584
rect 47730 21528 48514 21584
rect 47669 21526 48514 21528
rect 47669 21523 47735 21526
rect 23381 21450 23447 21453
rect 26049 21450 26115 21453
rect 37181 21450 37247 21453
rect 45185 21450 45251 21453
rect 23381 21448 37106 21450
rect 23381 21392 23386 21448
rect 23442 21392 26054 21448
rect 26110 21392 37106 21448
rect 23381 21390 37106 21392
rect 23381 21387 23447 21390
rect 26049 21387 26115 21390
rect 25865 21314 25931 21317
rect 30414 21314 30420 21316
rect 25865 21312 30420 21314
rect 25865 21256 25870 21312
rect 25926 21256 30420 21312
rect 25865 21254 30420 21256
rect 25865 21251 25931 21254
rect 30414 21252 30420 21254
rect 30484 21252 30490 21316
rect 37046 21314 37106 21390
rect 37181 21448 45251 21450
rect 37181 21392 37186 21448
rect 37242 21392 45190 21448
rect 45246 21392 45251 21448
rect 37181 21390 45251 21392
rect 37181 21387 37247 21390
rect 45185 21387 45251 21390
rect 49325 21450 49391 21453
rect 50200 21450 51000 21480
rect 49325 21448 51000 21450
rect 49325 21392 49330 21448
rect 49386 21392 51000 21448
rect 49325 21390 51000 21392
rect 49325 21387 49391 21390
rect 50200 21360 51000 21390
rect 40033 21314 40099 21317
rect 37046 21312 40099 21314
rect 37046 21256 40038 21312
rect 40094 21256 40099 21312
rect 37046 21254 40099 21256
rect 40033 21251 40099 21254
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 25221 21178 25287 21181
rect 26141 21178 26207 21181
rect 25221 21176 26207 21178
rect 25221 21120 25226 21176
rect 25282 21120 26146 21176
rect 26202 21120 26207 21176
rect 25221 21118 26207 21120
rect 25221 21115 25287 21118
rect 26141 21115 26207 21118
rect 27061 21178 27127 21181
rect 29729 21178 29795 21181
rect 27061 21176 29795 21178
rect 27061 21120 27066 21176
rect 27122 21120 29734 21176
rect 29790 21120 29795 21176
rect 27061 21118 29795 21120
rect 27061 21115 27127 21118
rect 29729 21115 29795 21118
rect 37549 21178 37615 21181
rect 40309 21178 40375 21181
rect 37549 21176 40375 21178
rect 37549 21120 37554 21176
rect 37610 21120 40314 21176
rect 40370 21120 40375 21176
rect 37549 21118 40375 21120
rect 37549 21115 37615 21118
rect 40309 21115 40375 21118
rect 28809 21042 28875 21045
rect 22694 21040 28875 21042
rect 22694 20984 28814 21040
rect 28870 20984 28875 21040
rect 22694 20982 28875 20984
rect 12893 20979 12959 20982
rect 21817 20979 21883 20982
rect 22461 20979 22527 20982
rect 28809 20979 28875 20982
rect 32857 21042 32923 21045
rect 45461 21042 45527 21045
rect 32857 21040 45527 21042
rect 32857 20984 32862 21040
rect 32918 20984 45466 21040
rect 45522 20984 45527 21040
rect 32857 20982 45527 20984
rect 32857 20979 32923 20982
rect 45461 20979 45527 20982
rect 49233 21042 49299 21045
rect 50200 21042 51000 21072
rect 49233 21040 51000 21042
rect 49233 20984 49238 21040
rect 49294 20984 51000 21040
rect 49233 20982 51000 20984
rect 49233 20979 49299 20982
rect 50200 20952 51000 20982
rect 8385 20906 8451 20909
rect 23657 20906 23723 20909
rect 8385 20904 23723 20906
rect 8385 20848 8390 20904
rect 8446 20848 23662 20904
rect 23718 20848 23723 20904
rect 8385 20846 23723 20848
rect 8385 20843 8451 20846
rect 23657 20843 23723 20846
rect 25957 20906 26023 20909
rect 26509 20906 26575 20909
rect 25957 20904 26575 20906
rect 25957 20848 25962 20904
rect 26018 20848 26514 20904
rect 26570 20848 26575 20904
rect 25957 20846 26575 20848
rect 25957 20843 26023 20846
rect 26509 20843 26575 20846
rect 27337 20906 27403 20909
rect 29494 20906 29500 20908
rect 27337 20904 29500 20906
rect 27337 20848 27342 20904
rect 27398 20848 29500 20904
rect 27337 20846 29500 20848
rect 27337 20843 27403 20846
rect 29494 20844 29500 20846
rect 29564 20844 29570 20908
rect 30557 20906 30623 20909
rect 31385 20906 31451 20909
rect 38377 20906 38443 20909
rect 41413 20906 41479 20909
rect 30557 20904 38443 20906
rect 30557 20848 30562 20904
rect 30618 20848 31390 20904
rect 31446 20848 38382 20904
rect 38438 20848 38443 20904
rect 30557 20846 38443 20848
rect 30557 20843 30623 20846
rect 31385 20843 31451 20846
rect 38377 20843 38443 20846
rect 38518 20904 41479 20906
rect 38518 20848 41418 20904
rect 41474 20848 41479 20904
rect 38518 20846 41479 20848
rect 0 20770 800 20800
rect 38518 20773 38578 20846
rect 41413 20843 41479 20846
rect 1025 20770 1091 20773
rect 0 20768 1091 20770
rect 0 20712 1030 20768
rect 1086 20712 1091 20768
rect 0 20710 1091 20712
rect 0 20680 800 20710
rect 1025 20707 1091 20710
rect 11789 20770 11855 20773
rect 19333 20770 19399 20773
rect 20345 20770 20411 20773
rect 11789 20768 17280 20770
rect 11789 20712 11794 20768
rect 11850 20712 17280 20768
rect 11789 20710 17280 20712
rect 11789 20707 11855 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 12433 20498 12499 20501
rect 13813 20498 13879 20501
rect 12433 20496 13879 20498
rect 12433 20440 12438 20496
rect 12494 20440 13818 20496
rect 13874 20440 13879 20496
rect 12433 20438 13879 20440
rect 17220 20498 17280 20710
rect 19333 20768 20411 20770
rect 19333 20712 19338 20768
rect 19394 20712 20350 20768
rect 20406 20712 20411 20768
rect 19333 20710 20411 20712
rect 19333 20707 19399 20710
rect 20345 20707 20411 20710
rect 22461 20770 22527 20773
rect 25129 20770 25195 20773
rect 22461 20768 25195 20770
rect 22461 20712 22466 20768
rect 22522 20712 25134 20768
rect 25190 20712 25195 20768
rect 22461 20710 25195 20712
rect 22461 20707 22527 20710
rect 25129 20707 25195 20710
rect 25589 20770 25655 20773
rect 26233 20770 26299 20773
rect 25589 20768 26299 20770
rect 25589 20712 25594 20768
rect 25650 20712 26238 20768
rect 26294 20712 26299 20768
rect 25589 20710 26299 20712
rect 25589 20707 25655 20710
rect 26233 20707 26299 20710
rect 35249 20770 35315 20773
rect 37273 20770 37339 20773
rect 35249 20768 37339 20770
rect 35249 20712 35254 20768
rect 35310 20712 37278 20768
rect 37334 20712 37339 20768
rect 35249 20710 37339 20712
rect 35249 20707 35315 20710
rect 37273 20707 37339 20710
rect 38469 20768 38578 20773
rect 38469 20712 38474 20768
rect 38530 20712 38578 20768
rect 38469 20710 38578 20712
rect 40033 20770 40099 20773
rect 41045 20770 41111 20773
rect 47393 20770 47459 20773
rect 40033 20768 47459 20770
rect 40033 20712 40038 20768
rect 40094 20712 41050 20768
rect 41106 20712 47398 20768
rect 47454 20712 47459 20768
rect 40033 20710 47459 20712
rect 38469 20707 38535 20710
rect 40033 20707 40099 20710
rect 41045 20707 41111 20710
rect 47393 20707 47459 20710
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 49325 20634 49391 20637
rect 50200 20634 51000 20664
rect 49325 20632 51000 20634
rect 49325 20576 49330 20632
rect 49386 20576 51000 20632
rect 49325 20574 51000 20576
rect 49325 20571 49391 20574
rect 50200 20544 51000 20574
rect 22185 20498 22251 20501
rect 25221 20498 25287 20501
rect 31017 20498 31083 20501
rect 31661 20498 31727 20501
rect 17220 20496 31727 20498
rect 17220 20440 22190 20496
rect 22246 20440 25226 20496
rect 25282 20440 31022 20496
rect 31078 20440 31666 20496
rect 31722 20440 31727 20496
rect 17220 20438 31727 20440
rect 12433 20435 12499 20438
rect 13813 20435 13879 20438
rect 22185 20435 22251 20438
rect 25221 20435 25287 20438
rect 31017 20435 31083 20438
rect 31661 20435 31727 20438
rect 34605 20498 34671 20501
rect 46289 20498 46355 20501
rect 34605 20496 46355 20498
rect 34605 20440 34610 20496
rect 34666 20440 46294 20496
rect 46350 20440 46355 20496
rect 34605 20438 46355 20440
rect 34605 20435 34671 20438
rect 46289 20435 46355 20438
rect 0 20362 800 20392
rect 1301 20362 1367 20365
rect 0 20360 1367 20362
rect 0 20304 1306 20360
rect 1362 20304 1367 20360
rect 0 20302 1367 20304
rect 0 20272 800 20302
rect 1301 20299 1367 20302
rect 11053 20362 11119 20365
rect 11881 20362 11947 20365
rect 11053 20360 11947 20362
rect 11053 20304 11058 20360
rect 11114 20304 11886 20360
rect 11942 20304 11947 20360
rect 11053 20302 11947 20304
rect 11053 20299 11119 20302
rect 11881 20299 11947 20302
rect 12709 20362 12775 20365
rect 31937 20362 32003 20365
rect 46565 20362 46631 20365
rect 12709 20360 13508 20362
rect 12709 20304 12714 20360
rect 12770 20304 13508 20360
rect 12709 20302 13508 20304
rect 12709 20299 12775 20302
rect 13448 20226 13508 20302
rect 31937 20360 46631 20362
rect 31937 20304 31942 20360
rect 31998 20304 46570 20360
rect 46626 20304 46631 20360
rect 31937 20302 46631 20304
rect 31937 20299 32003 20302
rect 46565 20299 46631 20302
rect 13629 20226 13695 20229
rect 22737 20226 22803 20229
rect 13448 20224 22803 20226
rect 13448 20168 13634 20224
rect 13690 20168 22742 20224
rect 22798 20168 22803 20224
rect 13448 20166 22803 20168
rect 13629 20163 13695 20166
rect 22737 20163 22803 20166
rect 48405 20226 48471 20229
rect 50200 20226 51000 20256
rect 48405 20224 51000 20226
rect 48405 20168 48410 20224
rect 48466 20168 51000 20224
rect 48405 20166 51000 20168
rect 48405 20163 48471 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 50200 20136 51000 20166
rect 42946 20095 43262 20096
rect 0 19954 800 19984
rect 1761 19954 1827 19957
rect 0 19952 1827 19954
rect 0 19896 1766 19952
rect 1822 19896 1827 19952
rect 0 19894 1827 19896
rect 0 19864 800 19894
rect 1761 19891 1827 19894
rect 11421 19954 11487 19957
rect 18689 19954 18755 19957
rect 23381 19954 23447 19957
rect 11421 19952 23447 19954
rect 11421 19896 11426 19952
rect 11482 19896 18694 19952
rect 18750 19896 23386 19952
rect 23442 19896 23447 19952
rect 11421 19894 23447 19896
rect 11421 19891 11487 19894
rect 18689 19891 18755 19894
rect 23381 19891 23447 19894
rect 26049 19954 26115 19957
rect 29545 19954 29611 19957
rect 43989 19954 44055 19957
rect 26049 19952 44055 19954
rect 26049 19896 26054 19952
rect 26110 19896 29550 19952
rect 29606 19896 43994 19952
rect 44050 19896 44055 19952
rect 26049 19894 44055 19896
rect 26049 19891 26115 19894
rect 29545 19891 29611 19894
rect 43989 19891 44055 19894
rect 10777 19818 10843 19821
rect 15653 19818 15719 19821
rect 10777 19816 15719 19818
rect 10777 19760 10782 19816
rect 10838 19760 15658 19816
rect 15714 19760 15719 19816
rect 10777 19758 15719 19760
rect 10777 19755 10843 19758
rect 15653 19755 15719 19758
rect 16665 19818 16731 19821
rect 17217 19818 17283 19821
rect 30097 19818 30163 19821
rect 16665 19816 30163 19818
rect 16665 19760 16670 19816
rect 16726 19760 17222 19816
rect 17278 19760 30102 19816
rect 30158 19760 30163 19816
rect 16665 19758 30163 19760
rect 16665 19755 16731 19758
rect 17217 19755 17283 19758
rect 30097 19755 30163 19758
rect 30373 19818 30439 19821
rect 39757 19818 39823 19821
rect 30373 19816 39823 19818
rect 30373 19760 30378 19816
rect 30434 19760 39762 19816
rect 39818 19760 39823 19816
rect 30373 19758 39823 19760
rect 30373 19755 30439 19758
rect 39757 19755 39823 19758
rect 49325 19818 49391 19821
rect 50200 19818 51000 19848
rect 49325 19816 51000 19818
rect 49325 19760 49330 19816
rect 49386 19760 51000 19816
rect 49325 19758 51000 19760
rect 49325 19755 49391 19758
rect 50200 19728 51000 19758
rect 19333 19682 19399 19685
rect 27153 19682 27219 19685
rect 19333 19680 27219 19682
rect 19333 19624 19338 19680
rect 19394 19624 27158 19680
rect 27214 19624 27219 19680
rect 19333 19622 27219 19624
rect 19333 19619 19399 19622
rect 27153 19619 27219 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2865 19546 2931 19549
rect 0 19544 2931 19546
rect 0 19488 2870 19544
rect 2926 19488 2931 19544
rect 0 19486 2931 19488
rect 0 19456 800 19486
rect 2865 19483 2931 19486
rect 23749 19546 23815 19549
rect 28625 19546 28691 19549
rect 33777 19546 33843 19549
rect 23749 19544 26434 19546
rect 23749 19488 23754 19544
rect 23810 19488 26434 19544
rect 23749 19486 26434 19488
rect 23749 19483 23815 19486
rect 15929 19410 15995 19413
rect 17493 19410 17559 19413
rect 26141 19410 26207 19413
rect 15929 19408 26207 19410
rect 15929 19352 15934 19408
rect 15990 19352 17498 19408
rect 17554 19352 26146 19408
rect 26202 19352 26207 19408
rect 15929 19350 26207 19352
rect 26374 19410 26434 19486
rect 28625 19544 33843 19546
rect 28625 19488 28630 19544
rect 28686 19488 33782 19544
rect 33838 19488 33843 19544
rect 28625 19486 33843 19488
rect 28625 19483 28691 19486
rect 33777 19483 33843 19486
rect 28349 19410 28415 19413
rect 28574 19410 28580 19412
rect 26374 19408 28580 19410
rect 26374 19352 28354 19408
rect 28410 19352 28580 19408
rect 26374 19350 28580 19352
rect 15929 19347 15995 19350
rect 17493 19347 17559 19350
rect 26141 19347 26207 19350
rect 28349 19347 28415 19350
rect 28574 19348 28580 19350
rect 28644 19348 28650 19412
rect 29545 19350 29611 19353
rect 29502 19348 29611 19350
rect 29502 19292 29550 19348
rect 29606 19292 29611 19348
rect 29502 19287 29611 19292
rect 29729 19348 29795 19353
rect 30414 19348 30420 19412
rect 30484 19410 30490 19412
rect 40585 19410 40651 19413
rect 30484 19408 40651 19410
rect 30484 19352 40590 19408
rect 40646 19352 40651 19408
rect 30484 19350 40651 19352
rect 30484 19348 30490 19350
rect 29729 19292 29734 19348
rect 29790 19292 29795 19348
rect 40585 19347 40651 19350
rect 49417 19410 49483 19413
rect 50200 19410 51000 19440
rect 49417 19408 51000 19410
rect 49417 19352 49422 19408
rect 49478 19352 51000 19408
rect 49417 19350 51000 19352
rect 49417 19347 49483 19350
rect 50200 19320 51000 19350
rect 29729 19287 29795 19292
rect 30005 19308 30071 19311
rect 30005 19306 30114 19308
rect 11053 19274 11119 19277
rect 15193 19274 15259 19277
rect 11053 19272 15259 19274
rect 11053 19216 11058 19272
rect 11114 19216 15198 19272
rect 15254 19216 15259 19272
rect 11053 19214 15259 19216
rect 11053 19211 11119 19214
rect 15193 19211 15259 19214
rect 19425 19274 19491 19277
rect 20529 19274 20595 19277
rect 29177 19276 29243 19277
rect 19425 19272 20595 19274
rect 19425 19216 19430 19272
rect 19486 19216 20534 19272
rect 20590 19216 20595 19272
rect 19425 19214 20595 19216
rect 19425 19211 19491 19214
rect 20529 19211 20595 19214
rect 29126 19212 29132 19276
rect 29196 19274 29243 19276
rect 29196 19272 29288 19274
rect 29238 19216 29288 19272
rect 29196 19214 29288 19216
rect 29196 19212 29243 19214
rect 29177 19211 29243 19212
rect 0 19138 800 19168
rect 29502 19141 29562 19287
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 5257 19138 5323 19141
rect 11973 19138 12039 19141
rect 5257 19136 12039 19138
rect 5257 19080 5262 19136
rect 5318 19080 11978 19136
rect 12034 19080 12039 19136
rect 5257 19078 12039 19080
rect 29502 19136 29611 19141
rect 29502 19080 29550 19136
rect 29606 19080 29611 19136
rect 29502 19078 29611 19080
rect 29732 19138 29792 19287
rect 30005 19250 30010 19306
rect 30066 19274 30114 19306
rect 32765 19274 32831 19277
rect 44265 19274 44331 19277
rect 30066 19272 32831 19274
rect 30066 19250 32770 19272
rect 30005 19245 32770 19250
rect 30054 19216 32770 19245
rect 32826 19216 32831 19272
rect 30054 19214 32831 19216
rect 32765 19211 32831 19214
rect 33366 19272 44331 19274
rect 33366 19216 44270 19272
rect 44326 19216 44331 19272
rect 33366 19214 44331 19216
rect 30189 19138 30255 19141
rect 29732 19136 30255 19138
rect 29732 19080 30194 19136
rect 30250 19080 30255 19136
rect 29732 19078 30255 19080
rect 5257 19075 5323 19078
rect 11973 19075 12039 19078
rect 29545 19075 29611 19078
rect 30189 19075 30255 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 24577 19002 24643 19005
rect 26141 19002 26207 19005
rect 27429 19002 27495 19005
rect 24577 19000 27495 19002
rect 24577 18944 24582 19000
rect 24638 18944 26146 19000
rect 26202 18944 27434 19000
rect 27490 18944 27495 19000
rect 24577 18942 27495 18944
rect 24577 18939 24643 18942
rect 26141 18939 26207 18942
rect 27429 18939 27495 18942
rect 29637 19002 29703 19005
rect 30741 19002 30807 19005
rect 29637 19000 30807 19002
rect 29637 18944 29642 19000
rect 29698 18944 30746 19000
rect 30802 18944 30807 19000
rect 29637 18942 30807 18944
rect 29637 18939 29703 18942
rect 30741 18939 30807 18942
rect 20621 18866 20687 18869
rect 29177 18866 29243 18869
rect 20621 18864 29243 18866
rect 20621 18808 20626 18864
rect 20682 18808 29182 18864
rect 29238 18808 29243 18864
rect 20621 18806 29243 18808
rect 20621 18803 20687 18806
rect 29177 18803 29243 18806
rect 30741 18866 30807 18869
rect 33366 18866 33426 19214
rect 44265 19211 44331 19214
rect 34646 19076 34652 19140
rect 34716 19138 34722 19140
rect 34789 19138 34855 19141
rect 36905 19138 36971 19141
rect 37641 19138 37707 19141
rect 38510 19138 38516 19140
rect 34716 19136 38516 19138
rect 34716 19080 34794 19136
rect 34850 19080 36910 19136
rect 36966 19080 37646 19136
rect 37702 19080 38516 19136
rect 34716 19078 38516 19080
rect 34716 19076 34722 19078
rect 34789 19075 34855 19078
rect 36905 19075 36971 19078
rect 37641 19075 37707 19078
rect 38510 19076 38516 19078
rect 38580 19076 38586 19140
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 33593 19002 33659 19005
rect 36077 19002 36143 19005
rect 33593 19000 36143 19002
rect 33593 18944 33598 19000
rect 33654 18944 36082 19000
rect 36138 18944 36143 19000
rect 33593 18942 36143 18944
rect 33593 18939 33659 18942
rect 36077 18939 36143 18942
rect 37089 19002 37155 19005
rect 41321 19002 41387 19005
rect 37089 19000 41387 19002
rect 37089 18944 37094 19000
rect 37150 18944 41326 19000
rect 41382 18944 41387 19000
rect 37089 18942 41387 18944
rect 37089 18939 37155 18942
rect 41321 18939 41387 18942
rect 49325 19002 49391 19005
rect 50200 19002 51000 19032
rect 49325 19000 51000 19002
rect 49325 18944 49330 19000
rect 49386 18944 51000 19000
rect 49325 18942 51000 18944
rect 49325 18939 49391 18942
rect 50200 18912 51000 18942
rect 30741 18864 33426 18866
rect 30741 18808 30746 18864
rect 30802 18808 33426 18864
rect 30741 18806 33426 18808
rect 34145 18866 34211 18869
rect 47301 18866 47367 18869
rect 34145 18864 47367 18866
rect 34145 18808 34150 18864
rect 34206 18808 47306 18864
rect 47362 18808 47367 18864
rect 34145 18806 47367 18808
rect 30741 18803 30807 18806
rect 34145 18803 34211 18806
rect 47301 18803 47367 18806
rect 0 18730 800 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 800 18670
rect 1485 18667 1551 18670
rect 15653 18730 15719 18733
rect 16941 18730 17007 18733
rect 15653 18728 17007 18730
rect 15653 18672 15658 18728
rect 15714 18672 16946 18728
rect 17002 18672 17007 18728
rect 15653 18670 17007 18672
rect 15653 18667 15719 18670
rect 16941 18667 17007 18670
rect 28993 18730 29059 18733
rect 29126 18730 29132 18732
rect 28993 18728 29132 18730
rect 28993 18672 28998 18728
rect 29054 18672 29132 18728
rect 28993 18670 29132 18672
rect 28993 18667 29059 18670
rect 29126 18668 29132 18670
rect 29196 18668 29202 18732
rect 29494 18668 29500 18732
rect 29564 18730 29570 18732
rect 29637 18730 29703 18733
rect 29564 18728 29703 18730
rect 29564 18672 29642 18728
rect 29698 18672 29703 18728
rect 29564 18670 29703 18672
rect 29564 18668 29570 18670
rect 29637 18667 29703 18670
rect 32765 18730 32831 18733
rect 38009 18730 38075 18733
rect 32765 18728 38075 18730
rect 32765 18672 32770 18728
rect 32826 18672 38014 18728
rect 38070 18672 38075 18728
rect 32765 18670 38075 18672
rect 32765 18667 32831 18670
rect 38009 18667 38075 18670
rect 29085 18594 29151 18597
rect 32581 18594 32647 18597
rect 29085 18592 32647 18594
rect 29085 18536 29090 18592
rect 29146 18536 32586 18592
rect 32642 18536 32647 18592
rect 29085 18534 32647 18536
rect 29085 18531 29151 18534
rect 32581 18531 32647 18534
rect 33133 18594 33199 18597
rect 33869 18594 33935 18597
rect 33133 18592 33935 18594
rect 33133 18536 33138 18592
rect 33194 18536 33874 18592
rect 33930 18536 33935 18592
rect 33133 18534 33935 18536
rect 33133 18531 33199 18534
rect 33869 18531 33935 18534
rect 48405 18594 48471 18597
rect 50200 18594 51000 18624
rect 48405 18592 51000 18594
rect 48405 18536 48410 18592
rect 48466 18536 51000 18592
rect 48405 18534 51000 18536
rect 48405 18531 48471 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 12341 18458 12407 18461
rect 17769 18458 17835 18461
rect 12341 18456 17835 18458
rect 12341 18400 12346 18456
rect 12402 18400 17774 18456
rect 17830 18400 17835 18456
rect 12341 18398 17835 18400
rect 12341 18395 12407 18398
rect 17769 18395 17835 18398
rect 30925 18458 30991 18461
rect 30925 18456 37842 18458
rect 30925 18400 30930 18456
rect 30986 18400 37842 18456
rect 30925 18398 37842 18400
rect 30925 18395 30991 18398
rect 0 18322 800 18352
rect 1761 18322 1827 18325
rect 0 18320 1827 18322
rect 0 18264 1766 18320
rect 1822 18264 1827 18320
rect 0 18262 1827 18264
rect 0 18232 800 18262
rect 1761 18259 1827 18262
rect 13813 18322 13879 18325
rect 17033 18322 17099 18325
rect 13813 18320 17099 18322
rect 13813 18264 13818 18320
rect 13874 18264 17038 18320
rect 17094 18264 17099 18320
rect 13813 18262 17099 18264
rect 13813 18259 13879 18262
rect 17033 18259 17099 18262
rect 25129 18322 25195 18325
rect 25957 18322 26023 18325
rect 25129 18320 37658 18322
rect 25129 18264 25134 18320
rect 25190 18264 25962 18320
rect 26018 18264 37658 18320
rect 25129 18262 37658 18264
rect 25129 18259 25195 18262
rect 25957 18259 26023 18262
rect 17401 18186 17467 18189
rect 28349 18186 28415 18189
rect 37089 18186 37155 18189
rect 17401 18184 37155 18186
rect 17401 18128 17406 18184
rect 17462 18128 28354 18184
rect 28410 18128 37094 18184
rect 37150 18128 37155 18184
rect 17401 18126 37155 18128
rect 17401 18123 17467 18126
rect 28349 18123 28415 18126
rect 37089 18123 37155 18126
rect 17585 18050 17651 18053
rect 19425 18050 19491 18053
rect 25262 18050 25268 18052
rect 17585 18048 19491 18050
rect 17585 17992 17590 18048
rect 17646 17992 19430 18048
rect 19486 17992 19491 18048
rect 17585 17990 19491 17992
rect 17585 17987 17651 17990
rect 19425 17987 19491 17990
rect 23614 17990 25268 18050
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 10593 17778 10659 17781
rect 23614 17778 23674 17990
rect 25262 17988 25268 17990
rect 25332 17988 25338 18052
rect 37598 18050 37658 18262
rect 37782 18186 37842 18398
rect 41229 18186 41295 18189
rect 47669 18186 47735 18189
rect 37782 18184 47735 18186
rect 37782 18128 41234 18184
rect 41290 18128 47674 18184
rect 47730 18128 47735 18184
rect 37782 18126 47735 18128
rect 41229 18123 41295 18126
rect 47669 18123 47735 18126
rect 49417 18186 49483 18189
rect 50200 18186 51000 18216
rect 49417 18184 51000 18186
rect 49417 18128 49422 18184
rect 49478 18128 51000 18184
rect 49417 18126 51000 18128
rect 49417 18123 49483 18126
rect 50200 18096 51000 18126
rect 40401 18050 40467 18053
rect 37598 18048 40467 18050
rect 37598 17992 40406 18048
rect 40462 17992 40467 18048
rect 37598 17990 40467 17992
rect 40401 17987 40467 17990
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 26325 17914 26391 17917
rect 28901 17914 28967 17917
rect 26325 17912 28967 17914
rect 26325 17856 26330 17912
rect 26386 17856 28906 17912
rect 28962 17856 28967 17912
rect 26325 17854 28967 17856
rect 26325 17851 26391 17854
rect 28901 17851 28967 17854
rect 10593 17776 23674 17778
rect 10593 17720 10598 17776
rect 10654 17720 23674 17776
rect 10593 17718 23674 17720
rect 26601 17778 26667 17781
rect 46933 17778 46999 17781
rect 26601 17776 46999 17778
rect 26601 17720 26606 17776
rect 26662 17720 46938 17776
rect 46994 17720 46999 17776
rect 26601 17718 46999 17720
rect 10593 17715 10659 17718
rect 26601 17715 26667 17718
rect 46933 17715 46999 17718
rect 49325 17778 49391 17781
rect 50200 17778 51000 17808
rect 49325 17776 51000 17778
rect 49325 17720 49330 17776
rect 49386 17720 51000 17776
rect 49325 17718 51000 17720
rect 49325 17715 49391 17718
rect 50200 17688 51000 17718
rect 14273 17642 14339 17645
rect 24669 17642 24735 17645
rect 26233 17642 26299 17645
rect 14273 17640 26299 17642
rect 14273 17584 14278 17640
rect 14334 17584 24674 17640
rect 24730 17584 26238 17640
rect 26294 17584 26299 17640
rect 14273 17582 26299 17584
rect 14273 17579 14339 17582
rect 24669 17579 24735 17582
rect 26233 17579 26299 17582
rect 31109 17642 31175 17645
rect 33869 17642 33935 17645
rect 35525 17642 35591 17645
rect 31109 17640 35591 17642
rect 31109 17584 31114 17640
rect 31170 17584 33874 17640
rect 33930 17584 35530 17640
rect 35586 17584 35591 17640
rect 31109 17582 35591 17584
rect 31109 17579 31175 17582
rect 33869 17579 33935 17582
rect 35525 17579 35591 17582
rect 35709 17642 35775 17645
rect 48037 17642 48103 17645
rect 35709 17640 48103 17642
rect 35709 17584 35714 17640
rect 35770 17584 48042 17640
rect 48098 17584 48103 17640
rect 35709 17582 48103 17584
rect 35709 17579 35775 17582
rect 48037 17579 48103 17582
rect 0 17506 800 17536
rect 1761 17506 1827 17509
rect 0 17504 1827 17506
rect 0 17448 1766 17504
rect 1822 17448 1827 17504
rect 0 17446 1827 17448
rect 0 17416 800 17446
rect 1761 17443 1827 17446
rect 30097 17506 30163 17509
rect 35433 17506 35499 17509
rect 30097 17504 35499 17506
rect 30097 17448 30102 17504
rect 30158 17448 35438 17504
rect 35494 17448 35499 17504
rect 30097 17446 35499 17448
rect 30097 17443 30163 17446
rect 35433 17443 35499 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 49325 17370 49391 17373
rect 50200 17370 51000 17400
rect 49325 17368 51000 17370
rect 49325 17312 49330 17368
rect 49386 17312 51000 17368
rect 49325 17310 51000 17312
rect 49325 17307 49391 17310
rect 50200 17280 51000 17310
rect 14181 17234 14247 17237
rect 18454 17234 18460 17236
rect 14181 17232 18460 17234
rect 14181 17176 14186 17232
rect 14242 17176 18460 17232
rect 14181 17174 18460 17176
rect 14181 17171 14247 17174
rect 18454 17172 18460 17174
rect 18524 17234 18530 17236
rect 22369 17234 22435 17237
rect 27613 17234 27679 17237
rect 28165 17234 28231 17237
rect 41873 17234 41939 17237
rect 18524 17232 41939 17234
rect 18524 17176 22374 17232
rect 22430 17176 27618 17232
rect 27674 17176 28170 17232
rect 28226 17176 41878 17232
rect 41934 17176 41939 17232
rect 18524 17174 41939 17176
rect 18524 17172 18530 17174
rect 22369 17171 22435 17174
rect 27613 17171 27679 17174
rect 28165 17171 28231 17174
rect 41873 17171 41939 17174
rect 0 17098 800 17128
rect 1025 17098 1091 17101
rect 0 17096 1091 17098
rect 0 17040 1030 17096
rect 1086 17040 1091 17096
rect 0 17038 1091 17040
rect 0 17008 800 17038
rect 1025 17035 1091 17038
rect 22369 17098 22435 17101
rect 26969 17098 27035 17101
rect 22369 17096 27035 17098
rect 22369 17040 22374 17096
rect 22430 17040 26974 17096
rect 27030 17040 27035 17096
rect 22369 17038 27035 17040
rect 22369 17035 22435 17038
rect 26969 17035 27035 17038
rect 27981 17098 28047 17101
rect 28758 17098 28764 17100
rect 27981 17096 28764 17098
rect 27981 17040 27986 17096
rect 28042 17040 28764 17096
rect 27981 17038 28764 17040
rect 27981 17035 28047 17038
rect 28758 17036 28764 17038
rect 28828 17036 28834 17100
rect 47945 17098 48011 17101
rect 31710 17096 48011 17098
rect 31710 17040 47950 17096
rect 48006 17040 48011 17096
rect 31710 17038 48011 17040
rect 26233 16962 26299 16965
rect 28809 16962 28875 16965
rect 31710 16962 31770 17038
rect 47945 17035 48011 17038
rect 26233 16960 31770 16962
rect 26233 16904 26238 16960
rect 26294 16904 28814 16960
rect 28870 16904 31770 16960
rect 26233 16902 31770 16904
rect 48313 16962 48379 16965
rect 50200 16962 51000 16992
rect 48313 16960 51000 16962
rect 48313 16904 48318 16960
rect 48374 16904 51000 16960
rect 48313 16902 51000 16904
rect 26233 16899 26299 16902
rect 28809 16899 28875 16902
rect 48313 16899 48379 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 50200 16872 51000 16902
rect 42946 16831 43262 16832
rect 0 16690 800 16720
rect 933 16690 999 16693
rect 0 16688 999 16690
rect 0 16632 938 16688
rect 994 16632 999 16688
rect 0 16630 999 16632
rect 0 16600 800 16630
rect 933 16627 999 16630
rect 15101 16692 15167 16693
rect 15101 16688 15148 16692
rect 15212 16690 15218 16692
rect 30189 16690 30255 16693
rect 36629 16690 36695 16693
rect 15101 16632 15106 16688
rect 15101 16628 15148 16632
rect 15212 16630 15258 16690
rect 30189 16688 36695 16690
rect 30189 16632 30194 16688
rect 30250 16632 36634 16688
rect 36690 16632 36695 16688
rect 30189 16630 36695 16632
rect 15212 16628 15218 16630
rect 15101 16627 15167 16628
rect 30189 16627 30255 16630
rect 36629 16627 36695 16630
rect 38510 16628 38516 16692
rect 38580 16690 38586 16692
rect 40217 16690 40283 16693
rect 38580 16688 40283 16690
rect 38580 16632 40222 16688
rect 40278 16632 40283 16688
rect 38580 16630 40283 16632
rect 38580 16628 38586 16630
rect 40217 16627 40283 16630
rect 38285 16554 38351 16557
rect 39941 16554 40007 16557
rect 38285 16552 40007 16554
rect 38285 16496 38290 16552
rect 38346 16496 39946 16552
rect 40002 16496 40007 16552
rect 38285 16494 40007 16496
rect 38285 16491 38351 16494
rect 39941 16491 40007 16494
rect 48221 16554 48287 16557
rect 50200 16554 51000 16584
rect 48221 16552 51000 16554
rect 48221 16496 48226 16552
rect 48282 16496 51000 16552
rect 48221 16494 51000 16496
rect 48221 16491 48287 16494
rect 50200 16464 51000 16494
rect 18597 16418 18663 16421
rect 18781 16418 18847 16421
rect 18597 16416 18847 16418
rect 18597 16360 18602 16416
rect 18658 16360 18786 16416
rect 18842 16360 18847 16416
rect 18597 16358 18847 16360
rect 18597 16355 18663 16358
rect 18781 16355 18847 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1025 16282 1091 16285
rect 0 16280 1091 16282
rect 0 16224 1030 16280
rect 1086 16224 1091 16280
rect 0 16222 1091 16224
rect 0 16192 800 16222
rect 1025 16219 1091 16222
rect 11605 16282 11671 16285
rect 17401 16282 17467 16285
rect 11605 16280 17467 16282
rect 11605 16224 11610 16280
rect 11666 16224 17406 16280
rect 17462 16224 17467 16280
rect 11605 16222 17467 16224
rect 11605 16219 11671 16222
rect 17401 16219 17467 16222
rect 33685 16282 33751 16285
rect 36353 16282 36419 16285
rect 33685 16280 36419 16282
rect 33685 16224 33690 16280
rect 33746 16224 36358 16280
rect 36414 16224 36419 16280
rect 33685 16222 36419 16224
rect 33685 16219 33751 16222
rect 36353 16219 36419 16222
rect 14181 16146 14247 16149
rect 15837 16146 15903 16149
rect 27061 16146 27127 16149
rect 35709 16146 35775 16149
rect 14181 16144 22110 16146
rect 14181 16088 14186 16144
rect 14242 16088 15842 16144
rect 15898 16088 22110 16144
rect 14181 16086 22110 16088
rect 14181 16083 14247 16086
rect 15837 16083 15903 16086
rect 11053 16010 11119 16013
rect 16665 16010 16731 16013
rect 11053 16008 16731 16010
rect 11053 15952 11058 16008
rect 11114 15952 16670 16008
rect 16726 15952 16731 16008
rect 11053 15950 16731 15952
rect 22050 16010 22110 16086
rect 27061 16144 35775 16146
rect 27061 16088 27066 16144
rect 27122 16088 35714 16144
rect 35770 16088 35775 16144
rect 27061 16086 35775 16088
rect 27061 16083 27127 16086
rect 35709 16083 35775 16086
rect 49325 16146 49391 16149
rect 50200 16146 51000 16176
rect 49325 16144 51000 16146
rect 49325 16088 49330 16144
rect 49386 16088 51000 16144
rect 49325 16086 51000 16088
rect 49325 16083 49391 16086
rect 50200 16056 51000 16086
rect 29361 16010 29427 16013
rect 22050 16008 29427 16010
rect 22050 15952 29366 16008
rect 29422 15952 29427 16008
rect 22050 15950 29427 15952
rect 11053 15947 11119 15950
rect 16665 15947 16731 15950
rect 29361 15947 29427 15950
rect 35709 16010 35775 16013
rect 49141 16010 49207 16013
rect 35709 16008 49207 16010
rect 35709 15952 35714 16008
rect 35770 15952 49146 16008
rect 49202 15952 49207 16008
rect 35709 15950 49207 15952
rect 35709 15947 35775 15950
rect 49141 15947 49207 15950
rect 0 15874 800 15904
rect 1025 15874 1091 15877
rect 0 15872 1091 15874
rect 0 15816 1030 15872
rect 1086 15816 1091 15872
rect 0 15814 1091 15816
rect 0 15784 800 15814
rect 1025 15811 1091 15814
rect 19006 15812 19012 15876
rect 19076 15874 19082 15876
rect 19149 15874 19215 15877
rect 19076 15872 19215 15874
rect 19076 15816 19154 15872
rect 19210 15816 19215 15872
rect 19076 15814 19215 15816
rect 19076 15812 19082 15814
rect 19149 15811 19215 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 22737 15738 22803 15741
rect 17910 15736 22803 15738
rect 17910 15680 22742 15736
rect 22798 15680 22803 15736
rect 17910 15678 22803 15680
rect 12341 15602 12407 15605
rect 13261 15602 13327 15605
rect 12341 15600 13327 15602
rect 12341 15544 12346 15600
rect 12402 15544 13266 15600
rect 13322 15544 13327 15600
rect 12341 15542 13327 15544
rect 12341 15539 12407 15542
rect 13261 15539 13327 15542
rect 0 15466 800 15496
rect 933 15466 999 15469
rect 0 15464 999 15466
rect 0 15408 938 15464
rect 994 15408 999 15464
rect 0 15406 999 15408
rect 0 15376 800 15406
rect 933 15403 999 15406
rect 11513 15466 11579 15469
rect 14641 15466 14707 15469
rect 15745 15466 15811 15469
rect 17910 15466 17970 15678
rect 22737 15675 22803 15678
rect 48681 15738 48747 15741
rect 50200 15738 51000 15768
rect 48681 15736 51000 15738
rect 48681 15680 48686 15736
rect 48742 15680 51000 15736
rect 48681 15678 51000 15680
rect 48681 15675 48747 15678
rect 50200 15648 51000 15678
rect 18505 15602 18571 15605
rect 18781 15604 18847 15605
rect 18505 15600 18706 15602
rect 18505 15544 18510 15600
rect 18566 15544 18706 15600
rect 18505 15542 18706 15544
rect 18505 15539 18571 15542
rect 11513 15464 17970 15466
rect 11513 15408 11518 15464
rect 11574 15408 14646 15464
rect 14702 15408 15750 15464
rect 15806 15408 17970 15464
rect 11513 15406 17970 15408
rect 11513 15403 11579 15406
rect 14641 15403 14707 15406
rect 15745 15403 15811 15406
rect 10501 15330 10567 15333
rect 12433 15330 12499 15333
rect 10501 15328 12499 15330
rect 10501 15272 10506 15328
rect 10562 15272 12438 15328
rect 12494 15272 12499 15328
rect 10501 15270 12499 15272
rect 10501 15267 10567 15270
rect 12433 15267 12499 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 18646 15194 18706 15542
rect 18781 15600 18828 15604
rect 18892 15602 18898 15604
rect 27061 15602 27127 15605
rect 34881 15602 34947 15605
rect 18781 15544 18786 15600
rect 18781 15540 18828 15544
rect 18892 15542 18938 15602
rect 27061 15600 34947 15602
rect 27061 15544 27066 15600
rect 27122 15544 34886 15600
rect 34942 15544 34947 15600
rect 27061 15542 34947 15544
rect 18892 15540 18898 15542
rect 18781 15539 18847 15540
rect 27061 15539 27127 15542
rect 34881 15539 34947 15542
rect 25681 15466 25747 15469
rect 47853 15466 47919 15469
rect 25681 15464 47919 15466
rect 25681 15408 25686 15464
rect 25742 15408 47858 15464
rect 47914 15408 47919 15464
rect 25681 15406 47919 15408
rect 25681 15403 25747 15406
rect 47853 15403 47919 15406
rect 48589 15330 48655 15333
rect 50200 15330 51000 15360
rect 48589 15328 51000 15330
rect 48589 15272 48594 15328
rect 48650 15272 51000 15328
rect 48589 15270 51000 15272
rect 48589 15267 48655 15270
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 50200 15240 51000 15270
rect 47946 15199 48262 15200
rect 19241 15194 19307 15197
rect 18646 15192 19307 15194
rect 18646 15136 19246 15192
rect 19302 15136 19307 15192
rect 18646 15134 19307 15136
rect 19241 15131 19307 15134
rect 0 15058 800 15088
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14968 800 14998
rect 933 14995 999 14998
rect 12341 15058 12407 15061
rect 26325 15058 26391 15061
rect 12341 15056 19212 15058
rect 12341 15000 12346 15056
rect 12402 15024 19212 15056
rect 19290 15056 26391 15058
rect 19290 15024 26330 15056
rect 12402 15000 26330 15024
rect 26386 15000 26391 15056
rect 12341 14998 26391 15000
rect 12341 14995 12407 14998
rect 19152 14964 19350 14998
rect 26325 14995 26391 14998
rect 27337 15058 27403 15061
rect 47853 15058 47919 15061
rect 27337 15056 47919 15058
rect 27337 15000 27342 15056
rect 27398 15000 47858 15056
rect 47914 15000 47919 15056
rect 27337 14998 47919 15000
rect 27337 14995 27403 14998
rect 47853 14995 47919 14998
rect 14733 14922 14799 14925
rect 18965 14922 19031 14925
rect 14733 14920 19031 14922
rect 14733 14864 14738 14920
rect 14794 14864 18970 14920
rect 19026 14864 19031 14920
rect 14733 14862 19031 14864
rect 14733 14859 14799 14862
rect 18965 14859 19031 14862
rect 24853 14922 24919 14925
rect 48037 14922 48103 14925
rect 24853 14920 48103 14922
rect 24853 14864 24858 14920
rect 24914 14864 48042 14920
rect 48098 14864 48103 14920
rect 24853 14862 48103 14864
rect 24853 14859 24919 14862
rect 48037 14859 48103 14862
rect 49325 14922 49391 14925
rect 50200 14922 51000 14952
rect 49325 14920 51000 14922
rect 49325 14864 49330 14920
rect 49386 14864 51000 14920
rect 49325 14862 51000 14864
rect 49325 14859 49391 14862
rect 50200 14832 51000 14862
rect 13997 14786 14063 14789
rect 19149 14786 19215 14789
rect 13997 14784 19215 14786
rect 13997 14728 14002 14784
rect 14058 14728 19154 14784
rect 19210 14728 19215 14784
rect 13997 14726 19215 14728
rect 13997 14723 14063 14726
rect 19149 14723 19215 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 933 14650 999 14653
rect 18781 14652 18847 14653
rect 18781 14650 18828 14652
rect 0 14648 999 14650
rect 0 14592 938 14648
rect 994 14592 999 14648
rect 0 14590 999 14592
rect 18736 14648 18828 14650
rect 18736 14592 18786 14648
rect 18736 14590 18828 14592
rect 0 14560 800 14590
rect 933 14587 999 14590
rect 18781 14588 18828 14590
rect 18892 14588 18898 14652
rect 18781 14587 18847 14588
rect 11237 14514 11303 14517
rect 20989 14514 21055 14517
rect 35709 14514 35775 14517
rect 11237 14512 19810 14514
rect 11237 14456 11242 14512
rect 11298 14456 19810 14512
rect 11237 14454 19810 14456
rect 11237 14451 11303 14454
rect 19750 14378 19810 14454
rect 20989 14512 35775 14514
rect 20989 14456 20994 14512
rect 21050 14456 35714 14512
rect 35770 14456 35775 14512
rect 20989 14454 35775 14456
rect 20989 14451 21055 14454
rect 35709 14451 35775 14454
rect 37181 14514 37247 14517
rect 39297 14514 39363 14517
rect 37181 14512 39363 14514
rect 37181 14456 37186 14512
rect 37242 14456 39302 14512
rect 39358 14456 39363 14512
rect 37181 14454 39363 14456
rect 37181 14451 37247 14454
rect 39297 14451 39363 14454
rect 49325 14514 49391 14517
rect 50200 14514 51000 14544
rect 49325 14512 51000 14514
rect 49325 14456 49330 14512
rect 49386 14456 51000 14512
rect 49325 14454 51000 14456
rect 49325 14451 49391 14454
rect 50200 14424 51000 14454
rect 20621 14378 20687 14381
rect 21817 14378 21883 14381
rect 47945 14378 48011 14381
rect 19750 14376 48011 14378
rect 19750 14320 20626 14376
rect 20682 14320 21822 14376
rect 21878 14320 47950 14376
rect 48006 14320 48011 14376
rect 19750 14318 48011 14320
rect 20621 14315 20687 14318
rect 21817 14315 21883 14318
rect 47945 14315 48011 14318
rect 0 14242 800 14272
rect 1025 14242 1091 14245
rect 0 14240 1091 14242
rect 0 14184 1030 14240
rect 1086 14184 1091 14240
rect 0 14182 1091 14184
rect 0 14152 800 14182
rect 1025 14179 1091 14182
rect 9949 14242 10015 14245
rect 16849 14242 16915 14245
rect 9949 14240 16915 14242
rect 9949 14184 9954 14240
rect 10010 14184 16854 14240
rect 16910 14184 16915 14240
rect 9949 14182 16915 14184
rect 9949 14179 10015 14182
rect 16849 14179 16915 14182
rect 18597 14242 18663 14245
rect 19006 14242 19012 14244
rect 18597 14240 19012 14242
rect 18597 14184 18602 14240
rect 18658 14184 19012 14240
rect 18597 14182 19012 14184
rect 18597 14179 18663 14182
rect 19006 14180 19012 14182
rect 19076 14180 19082 14244
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 49325 14106 49391 14109
rect 50200 14106 51000 14136
rect 49325 14104 51000 14106
rect 49325 14048 49330 14104
rect 49386 14048 51000 14104
rect 49325 14046 51000 14048
rect 49325 14043 49391 14046
rect 50200 14016 51000 14046
rect 16297 13970 16363 13973
rect 18045 13970 18111 13973
rect 16297 13968 18111 13970
rect 16297 13912 16302 13968
rect 16358 13912 18050 13968
rect 18106 13912 18111 13968
rect 16297 13910 18111 13912
rect 16297 13907 16363 13910
rect 18045 13907 18111 13910
rect 0 13834 800 13864
rect 1761 13834 1827 13837
rect 0 13832 1827 13834
rect 0 13776 1766 13832
rect 1822 13776 1827 13832
rect 0 13774 1827 13776
rect 0 13744 800 13774
rect 1761 13771 1827 13774
rect 10501 13834 10567 13837
rect 20989 13834 21055 13837
rect 10501 13832 21055 13834
rect 10501 13776 10506 13832
rect 10562 13776 20994 13832
rect 21050 13776 21055 13832
rect 10501 13774 21055 13776
rect 10501 13771 10567 13774
rect 20989 13771 21055 13774
rect 15142 13636 15148 13700
rect 15212 13698 15218 13700
rect 16481 13698 16547 13701
rect 15212 13696 16547 13698
rect 15212 13640 16486 13696
rect 16542 13640 16547 13696
rect 15212 13638 16547 13640
rect 15212 13636 15218 13638
rect 16481 13635 16547 13638
rect 47669 13698 47735 13701
rect 50200 13698 51000 13728
rect 47669 13696 51000 13698
rect 47669 13640 47674 13696
rect 47730 13640 51000 13696
rect 47669 13638 51000 13640
rect 47669 13635 47735 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 50200 13608 51000 13638
rect 42946 13567 43262 13568
rect 13854 13500 13860 13564
rect 13924 13562 13930 13564
rect 17125 13562 17191 13565
rect 13924 13560 17191 13562
rect 13924 13504 17130 13560
rect 17186 13504 17191 13560
rect 13924 13502 17191 13504
rect 13924 13500 13930 13502
rect 17125 13499 17191 13502
rect 0 13426 800 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 800 13366
rect 3509 13363 3575 13366
rect 14089 13426 14155 13429
rect 14457 13426 14523 13429
rect 24577 13426 24643 13429
rect 14089 13424 14290 13426
rect 14089 13368 14094 13424
rect 14150 13368 14290 13424
rect 14089 13366 14290 13368
rect 14089 13363 14155 13366
rect 13997 13292 14063 13293
rect 13997 13288 14044 13292
rect 14108 13290 14114 13292
rect 14230 13290 14290 13366
rect 14457 13424 24643 13426
rect 14457 13368 14462 13424
rect 14518 13368 24582 13424
rect 24638 13368 24643 13424
rect 14457 13366 24643 13368
rect 14457 13363 14523 13366
rect 24577 13363 24643 13366
rect 14365 13290 14431 13293
rect 13997 13232 14002 13288
rect 13997 13228 14044 13232
rect 14108 13230 14154 13290
rect 14230 13288 14431 13290
rect 14230 13232 14370 13288
rect 14426 13232 14431 13288
rect 14230 13230 14431 13232
rect 14108 13228 14114 13230
rect 13997 13227 14063 13228
rect 14365 13227 14431 13230
rect 15009 13290 15075 13293
rect 17125 13290 17191 13293
rect 15009 13288 17191 13290
rect 15009 13232 15014 13288
rect 15070 13232 17130 13288
rect 17186 13232 17191 13288
rect 15009 13230 17191 13232
rect 15009 13227 15075 13230
rect 17125 13227 17191 13230
rect 17677 13290 17743 13293
rect 20897 13290 20963 13293
rect 17677 13288 20963 13290
rect 17677 13232 17682 13288
rect 17738 13232 20902 13288
rect 20958 13232 20963 13288
rect 17677 13230 20963 13232
rect 17677 13227 17743 13230
rect 20897 13227 20963 13230
rect 49141 13290 49207 13293
rect 50200 13290 51000 13320
rect 49141 13288 51000 13290
rect 49141 13232 49146 13288
rect 49202 13232 51000 13288
rect 49141 13230 51000 13232
rect 49141 13227 49207 13230
rect 50200 13200 51000 13230
rect 11329 13154 11395 13157
rect 14457 13154 14523 13157
rect 11329 13152 14523 13154
rect 11329 13096 11334 13152
rect 11390 13096 14462 13152
rect 14518 13096 14523 13152
rect 11329 13094 14523 13096
rect 11329 13091 11395 13094
rect 14457 13091 14523 13094
rect 28533 13154 28599 13157
rect 28809 13154 28875 13157
rect 28533 13152 28875 13154
rect 28533 13096 28538 13152
rect 28594 13096 28814 13152
rect 28870 13096 28875 13152
rect 28533 13094 28875 13096
rect 28533 13091 28599 13094
rect 28809 13091 28875 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 12893 13018 12959 13021
rect 15193 13018 15259 13021
rect 18505 13020 18571 13021
rect 12893 13016 15259 13018
rect 12893 12960 12898 13016
rect 12954 12960 15198 13016
rect 15254 12960 15259 13016
rect 12893 12958 15259 12960
rect 12893 12955 12959 12958
rect 15193 12955 15259 12958
rect 18454 12956 18460 13020
rect 18524 13018 18571 13020
rect 22829 13018 22895 13021
rect 26785 13018 26851 13021
rect 27153 13018 27219 13021
rect 18524 13016 18616 13018
rect 18566 12960 18616 13016
rect 18524 12958 18616 12960
rect 22829 13016 27219 13018
rect 22829 12960 22834 13016
rect 22890 12960 26790 13016
rect 26846 12960 27158 13016
rect 27214 12960 27219 13016
rect 22829 12958 27219 12960
rect 18524 12956 18571 12958
rect 18505 12955 18571 12956
rect 22829 12955 22895 12958
rect 26785 12955 26851 12958
rect 27153 12955 27219 12958
rect 18413 12884 18479 12885
rect 18413 12882 18460 12884
rect 18332 12880 18460 12882
rect 18524 12882 18530 12884
rect 30557 12882 30623 12885
rect 35157 12882 35223 12885
rect 36445 12882 36511 12885
rect 18524 12880 36511 12882
rect 18332 12824 18418 12880
rect 18524 12824 30562 12880
rect 30618 12824 35162 12880
rect 35218 12824 36450 12880
rect 36506 12824 36511 12880
rect 18332 12822 18460 12824
rect 18413 12820 18460 12822
rect 18524 12822 36511 12824
rect 18524 12820 18530 12822
rect 18413 12819 18479 12820
rect 30557 12819 30623 12822
rect 35157 12819 35223 12822
rect 36445 12819 36511 12822
rect 49141 12882 49207 12885
rect 50200 12882 51000 12912
rect 49141 12880 51000 12882
rect 49141 12824 49146 12880
rect 49202 12824 51000 12880
rect 49141 12822 51000 12824
rect 49141 12819 49207 12822
rect 50200 12792 51000 12822
rect 12249 12746 12315 12749
rect 16665 12746 16731 12749
rect 12249 12744 16731 12746
rect 12249 12688 12254 12744
rect 12310 12688 16670 12744
rect 16726 12688 16731 12744
rect 12249 12686 16731 12688
rect 12249 12683 12315 12686
rect 16665 12683 16731 12686
rect 22921 12746 22987 12749
rect 25221 12746 25287 12749
rect 22921 12744 25287 12746
rect 22921 12688 22926 12744
rect 22982 12688 25226 12744
rect 25282 12688 25287 12744
rect 22921 12686 25287 12688
rect 22921 12683 22987 12686
rect 25221 12683 25287 12686
rect 28625 12746 28691 12749
rect 40033 12746 40099 12749
rect 28625 12744 40099 12746
rect 28625 12688 28630 12744
rect 28686 12688 40038 12744
rect 40094 12688 40099 12744
rect 28625 12686 40099 12688
rect 28625 12683 28691 12686
rect 40033 12683 40099 12686
rect 0 12610 800 12640
rect 1301 12610 1367 12613
rect 0 12608 1367 12610
rect 0 12552 1306 12608
rect 1362 12552 1367 12608
rect 0 12550 1367 12552
rect 0 12520 800 12550
rect 1301 12547 1367 12550
rect 13997 12610 14063 12613
rect 14917 12610 14983 12613
rect 13997 12608 14983 12610
rect 13997 12552 14002 12608
rect 14058 12552 14922 12608
rect 14978 12552 14983 12608
rect 13997 12550 14983 12552
rect 13997 12547 14063 12550
rect 14917 12547 14983 12550
rect 20989 12610 21055 12613
rect 22737 12610 22803 12613
rect 20989 12608 22803 12610
rect 20989 12552 20994 12608
rect 21050 12552 22742 12608
rect 22798 12552 22803 12608
rect 20989 12550 22803 12552
rect 20989 12547 21055 12550
rect 22737 12547 22803 12550
rect 23565 12610 23631 12613
rect 24485 12610 24551 12613
rect 23565 12608 24551 12610
rect 23565 12552 23570 12608
rect 23626 12552 24490 12608
rect 24546 12552 24551 12608
rect 23565 12550 24551 12552
rect 23565 12547 23631 12550
rect 24485 12547 24551 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 22369 12338 22435 12341
rect 30097 12338 30163 12341
rect 22369 12336 30163 12338
rect 22369 12280 22374 12336
rect 22430 12280 30102 12336
rect 30158 12280 30163 12336
rect 22369 12278 30163 12280
rect 22369 12275 22435 12278
rect 30097 12275 30163 12278
rect 0 12202 800 12232
rect 1209 12202 1275 12205
rect 0 12200 1275 12202
rect 0 12144 1214 12200
rect 1270 12144 1275 12200
rect 0 12142 1275 12144
rect 0 12112 800 12142
rect 1209 12139 1275 12142
rect 13353 12066 13419 12069
rect 17217 12066 17283 12069
rect 13353 12064 17283 12066
rect 13353 12008 13358 12064
rect 13414 12008 17222 12064
rect 17278 12008 17283 12064
rect 13353 12006 17283 12008
rect 13353 12003 13419 12006
rect 17217 12003 17283 12006
rect 49141 12066 49207 12069
rect 50200 12066 51000 12096
rect 49141 12064 51000 12066
rect 49141 12008 49146 12064
rect 49202 12008 51000 12064
rect 49141 12006 51000 12008
rect 49141 12003 49207 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 50200 11976 51000 12006
rect 47946 11935 48262 11936
rect 0 11794 800 11824
rect 1301 11794 1367 11797
rect 0 11792 1367 11794
rect 0 11736 1306 11792
rect 1362 11736 1367 11792
rect 0 11734 1367 11736
rect 0 11704 800 11734
rect 1301 11731 1367 11734
rect 29729 11794 29795 11797
rect 40401 11794 40467 11797
rect 29729 11792 40467 11794
rect 29729 11736 29734 11792
rect 29790 11736 40406 11792
rect 40462 11736 40467 11792
rect 29729 11734 40467 11736
rect 29729 11731 29795 11734
rect 40401 11731 40467 11734
rect 30465 11658 30531 11661
rect 35617 11658 35683 11661
rect 30465 11656 35683 11658
rect 30465 11600 30470 11656
rect 30526 11600 35622 11656
rect 35678 11600 35683 11656
rect 30465 11598 35683 11600
rect 30465 11595 30531 11598
rect 35617 11595 35683 11598
rect 49141 11658 49207 11661
rect 50200 11658 51000 11688
rect 49141 11656 51000 11658
rect 49141 11600 49146 11656
rect 49202 11600 51000 11656
rect 49141 11598 51000 11600
rect 49141 11595 49207 11598
rect 50200 11568 51000 11598
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 1301 11386 1367 11389
rect 0 11384 1367 11386
rect 0 11328 1306 11384
rect 1362 11328 1367 11384
rect 0 11326 1367 11328
rect 0 11296 800 11326
rect 1301 11323 1367 11326
rect 49233 11250 49299 11253
rect 50200 11250 51000 11280
rect 49233 11248 51000 11250
rect 49233 11192 49238 11248
rect 49294 11192 51000 11248
rect 49233 11190 51000 11192
rect 49233 11187 49299 11190
rect 50200 11160 51000 11190
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 13445 10842 13511 10845
rect 17493 10842 17559 10845
rect 13445 10840 17559 10842
rect 13445 10784 13450 10840
rect 13506 10784 17498 10840
rect 17554 10784 17559 10840
rect 13445 10782 17559 10784
rect 13445 10779 13511 10782
rect 17493 10779 17559 10782
rect 49141 10842 49207 10845
rect 50200 10842 51000 10872
rect 49141 10840 51000 10842
rect 49141 10784 49146 10840
rect 49202 10784 51000 10840
rect 49141 10782 51000 10784
rect 49141 10779 49207 10782
rect 50200 10752 51000 10782
rect 13629 10706 13695 10709
rect 34646 10706 34652 10708
rect 13629 10704 34652 10706
rect 13629 10648 13634 10704
rect 13690 10648 34652 10704
rect 13629 10646 34652 10648
rect 13629 10643 13695 10646
rect 34646 10644 34652 10646
rect 34716 10644 34722 10708
rect 0 10570 800 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 800 10510
rect 1577 10507 1643 10510
rect 14273 10570 14339 10573
rect 15929 10570 15995 10573
rect 14273 10568 15995 10570
rect 14273 10512 14278 10568
rect 14334 10512 15934 10568
rect 15990 10512 15995 10568
rect 14273 10510 15995 10512
rect 14273 10507 14339 10510
rect 15929 10507 15995 10510
rect 30741 10570 30807 10573
rect 36537 10570 36603 10573
rect 30741 10568 36603 10570
rect 30741 10512 30746 10568
rect 30802 10512 36542 10568
rect 36598 10512 36603 10568
rect 30741 10510 36603 10512
rect 30741 10507 30807 10510
rect 36537 10507 36603 10510
rect 49325 10434 49391 10437
rect 50200 10434 51000 10464
rect 49325 10432 51000 10434
rect 49325 10376 49330 10432
rect 49386 10376 51000 10432
rect 49325 10374 51000 10376
rect 49325 10371 49391 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 1209 10162 1275 10165
rect 0 10160 1275 10162
rect 0 10104 1214 10160
rect 1270 10104 1275 10160
rect 0 10102 1275 10104
rect 0 10072 800 10102
rect 1209 10099 1275 10102
rect 13077 10162 13143 10165
rect 13854 10162 13860 10164
rect 13077 10160 13860 10162
rect 13077 10104 13082 10160
rect 13138 10104 13860 10160
rect 13077 10102 13860 10104
rect 13077 10099 13143 10102
rect 13854 10100 13860 10102
rect 13924 10100 13930 10164
rect 23749 10162 23815 10165
rect 27705 10162 27771 10165
rect 28625 10162 28691 10165
rect 23749 10160 28691 10162
rect 23749 10104 23754 10160
rect 23810 10104 27710 10160
rect 27766 10104 28630 10160
rect 28686 10104 28691 10160
rect 23749 10102 28691 10104
rect 23749 10099 23815 10102
rect 27705 10099 27771 10102
rect 28625 10099 28691 10102
rect 49233 10026 49299 10029
rect 50200 10026 51000 10056
rect 49233 10024 51000 10026
rect 49233 9968 49238 10024
rect 49294 9968 51000 10024
rect 49233 9966 51000 9968
rect 49233 9963 49299 9966
rect 50200 9936 51000 9966
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1301 9754 1367 9757
rect 0 9752 1367 9754
rect 0 9696 1306 9752
rect 1362 9696 1367 9752
rect 0 9694 1367 9696
rect 0 9664 800 9694
rect 1301 9691 1367 9694
rect 31753 9754 31819 9757
rect 32305 9754 32371 9757
rect 31753 9752 32371 9754
rect 31753 9696 31758 9752
rect 31814 9696 32310 9752
rect 32366 9696 32371 9752
rect 31753 9694 32371 9696
rect 31753 9691 31819 9694
rect 32305 9691 32371 9694
rect 16481 9618 16547 9621
rect 17769 9618 17835 9621
rect 21541 9618 21607 9621
rect 16481 9616 21607 9618
rect 16481 9560 16486 9616
rect 16542 9560 17774 9616
rect 17830 9560 21546 9616
rect 21602 9560 21607 9616
rect 16481 9558 21607 9560
rect 16481 9555 16547 9558
rect 17769 9555 17835 9558
rect 21541 9555 21607 9558
rect 47301 9618 47367 9621
rect 50200 9618 51000 9648
rect 47301 9616 51000 9618
rect 47301 9560 47306 9616
rect 47362 9560 51000 9616
rect 47301 9558 51000 9560
rect 47301 9555 47367 9558
rect 50200 9528 51000 9558
rect 3693 9482 3759 9485
rect 33501 9482 33567 9485
rect 3693 9480 33567 9482
rect 3693 9424 3698 9480
rect 3754 9424 33506 9480
rect 33562 9424 33567 9480
rect 3693 9422 33567 9424
rect 3693 9419 3759 9422
rect 33501 9419 33567 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9210 49207 9213
rect 50200 9210 51000 9240
rect 49141 9208 51000 9210
rect 49141 9152 49146 9208
rect 49202 9152 51000 9208
rect 49141 9150 51000 9152
rect 49141 9147 49207 9150
rect 50200 9120 51000 9150
rect 30925 9074 30991 9077
rect 35985 9074 36051 9077
rect 30925 9072 36051 9074
rect 30925 9016 30930 9072
rect 30986 9016 35990 9072
rect 36046 9016 36051 9072
rect 30925 9014 36051 9016
rect 30925 9011 30991 9014
rect 35985 9011 36051 9014
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 14038 8876 14044 8940
rect 14108 8938 14114 8940
rect 14365 8938 14431 8941
rect 25957 8938 26023 8941
rect 14108 8936 26023 8938
rect 14108 8880 14370 8936
rect 14426 8880 25962 8936
rect 26018 8880 26023 8936
rect 14108 8878 26023 8880
rect 14108 8876 14114 8878
rect 14365 8875 14431 8878
rect 25957 8875 26023 8878
rect 49325 8802 49391 8805
rect 50200 8802 51000 8832
rect 49325 8800 51000 8802
rect 49325 8744 49330 8800
rect 49386 8744 51000 8800
rect 49325 8742 51000 8744
rect 49325 8739 49391 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 50200 8712 51000 8742
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 49233 8394 49299 8397
rect 50200 8394 51000 8424
rect 49233 8392 51000 8394
rect 49233 8336 49238 8392
rect 49294 8336 51000 8392
rect 49233 8334 51000 8336
rect 49233 8331 49299 8334
rect 50200 8304 51000 8334
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 2405 8122 2471 8125
rect 0 8120 2471 8122
rect 0 8064 2410 8120
rect 2466 8064 2471 8120
rect 0 8062 2471 8064
rect 0 8032 800 8062
rect 2405 8059 2471 8062
rect 46841 7986 46907 7989
rect 50200 7986 51000 8016
rect 46841 7984 51000 7986
rect 46841 7928 46846 7984
rect 46902 7928 51000 7984
rect 46841 7926 51000 7928
rect 46841 7923 46907 7926
rect 50200 7896 51000 7926
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 49141 7578 49207 7581
rect 50200 7578 51000 7608
rect 49141 7576 51000 7578
rect 49141 7520 49146 7576
rect 49202 7520 51000 7576
rect 49141 7518 51000 7520
rect 49141 7515 49207 7518
rect 50200 7488 51000 7518
rect 0 7306 800 7336
rect 1577 7306 1643 7309
rect 0 7304 1643 7306
rect 0 7248 1582 7304
rect 1638 7248 1643 7304
rect 0 7246 1643 7248
rect 0 7216 800 7246
rect 1577 7243 1643 7246
rect 49325 7170 49391 7173
rect 50200 7170 51000 7200
rect 49325 7168 51000 7170
rect 49325 7112 49330 7168
rect 49386 7112 51000 7168
rect 49325 7110 51000 7112
rect 49325 7107 49391 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 50200 7080 51000 7110
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 3325 6898 3391 6901
rect 0 6896 3391 6898
rect 0 6840 3330 6896
rect 3386 6840 3391 6896
rect 0 6838 3391 6840
rect 0 6808 800 6838
rect 3325 6835 3391 6838
rect 2865 6762 2931 6765
rect 18454 6762 18460 6764
rect 2865 6760 18460 6762
rect 2865 6704 2870 6760
rect 2926 6704 18460 6760
rect 2865 6702 18460 6704
rect 2865 6699 2931 6702
rect 18454 6700 18460 6702
rect 18524 6700 18530 6764
rect 49233 6762 49299 6765
rect 50200 6762 51000 6792
rect 49233 6760 51000 6762
rect 49233 6704 49238 6760
rect 49294 6704 51000 6760
rect 49233 6702 51000 6704
rect 49233 6699 49299 6702
rect 50200 6672 51000 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 48681 6354 48747 6357
rect 50200 6354 51000 6384
rect 48681 6352 51000 6354
rect 48681 6296 48686 6352
rect 48742 6296 51000 6352
rect 48681 6294 51000 6296
rect 48681 6291 48747 6294
rect 50200 6264 51000 6294
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5946 49207 5949
rect 50200 5946 51000 5976
rect 49141 5944 51000 5946
rect 49141 5888 49146 5944
rect 49202 5888 51000 5944
rect 49141 5886 51000 5888
rect 49141 5883 49207 5886
rect 50200 5856 51000 5886
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 49417 5538 49483 5541
rect 50200 5538 51000 5568
rect 49417 5536 51000 5538
rect 49417 5480 49422 5536
rect 49478 5480 51000 5536
rect 49417 5478 51000 5480
rect 49417 5475 49483 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 50200 5448 51000 5478
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 1393 5266 1459 5269
rect 0 5264 1459 5266
rect 0 5208 1398 5264
rect 1454 5208 1459 5264
rect 0 5206 1459 5208
rect 0 5176 800 5206
rect 1393 5203 1459 5206
rect 49325 5130 49391 5133
rect 50200 5130 51000 5160
rect 49325 5128 51000 5130
rect 49325 5072 49330 5128
rect 49386 5072 51000 5128
rect 49325 5070 51000 5072
rect 49325 5067 49391 5070
rect 50200 5040 51000 5070
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 48313 4722 48379 4725
rect 50200 4722 51000 4752
rect 48313 4720 51000 4722
rect 48313 4664 48318 4720
rect 48374 4664 51000 4720
rect 48313 4662 51000 4664
rect 48313 4659 48379 4662
rect 50200 4632 51000 4662
rect 0 4450 800 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 800 4390
rect 1301 4387 1367 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4042 800 4072
rect 1301 4042 1367 4045
rect 0 4040 1367 4042
rect 0 3984 1306 4040
rect 1362 3984 1367 4040
rect 0 3982 1367 3984
rect 0 3952 800 3982
rect 1301 3979 1367 3982
rect 15745 4042 15811 4045
rect 27889 4042 27955 4045
rect 15745 4040 27955 4042
rect 15745 3984 15750 4040
rect 15806 3984 27894 4040
rect 27950 3984 27955 4040
rect 15745 3982 27955 3984
rect 15745 3979 15811 3982
rect 27889 3979 27955 3982
rect 49233 3906 49299 3909
rect 50200 3906 51000 3936
rect 49233 3904 51000 3906
rect 49233 3848 49238 3904
rect 49294 3848 51000 3904
rect 49233 3846 51000 3848
rect 49233 3843 49299 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 50200 3816 51000 3846
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1209 3634 1275 3637
rect 0 3632 1275 3634
rect 0 3576 1214 3632
rect 1270 3576 1275 3632
rect 0 3574 1275 3576
rect 0 3544 800 3574
rect 1209 3571 1275 3574
rect 49141 3498 49207 3501
rect 50200 3498 51000 3528
rect 49141 3496 51000 3498
rect 49141 3440 49146 3496
rect 49202 3440 51000 3496
rect 49141 3438 51000 3440
rect 49141 3435 49207 3438
rect 50200 3408 51000 3438
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 48681 3090 48747 3093
rect 50200 3090 51000 3120
rect 48681 3088 51000 3090
rect 48681 3032 48686 3088
rect 48742 3032 51000 3088
rect 48681 3030 51000 3032
rect 48681 3027 48747 3030
rect 50200 3000 51000 3030
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 46841 2682 46907 2685
rect 50200 2682 51000 2712
rect 46841 2680 51000 2682
rect 46841 2624 46846 2680
rect 46902 2624 51000 2680
rect 46841 2622 51000 2624
rect 46841 2619 46907 2622
rect 50200 2592 51000 2622
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 48497 2274 48563 2277
rect 50200 2274 51000 2304
rect 48497 2272 51000 2274
rect 48497 2216 48502 2272
rect 48558 2216 51000 2272
rect 48497 2214 51000 2216
rect 48497 2211 48563 2214
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 50200 2184 51000 2214
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 46749 1866 46815 1869
rect 50200 1866 51000 1896
rect 46749 1864 51000 1866
rect 46749 1808 46754 1864
rect 46810 1808 51000 1864
rect 46749 1806 51000 1808
rect 46749 1803 46815 1806
rect 50200 1776 51000 1806
rect 0 1594 800 1624
rect 4061 1594 4127 1597
rect 0 1592 4127 1594
rect 0 1536 4066 1592
rect 4122 1536 4127 1592
rect 0 1534 4127 1536
rect 0 1504 800 1534
rect 4061 1531 4127 1534
rect 46657 1458 46723 1461
rect 50200 1458 51000 1488
rect 46657 1456 51000 1458
rect 46657 1400 46662 1456
rect 46718 1400 51000 1456
rect 46657 1398 51000 1400
rect 46657 1395 46723 1398
rect 50200 1368 51000 1398
<< via3 >>
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 28580 24108 28644 24172
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 28948 23700 29012 23764
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 25268 22944 25332 22948
rect 25268 22888 25318 22944
rect 25318 22888 25332 22944
rect 25268 22884 25332 22888
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 30420 21252 30484 21316
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 29500 20844 29564 20908
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 28580 19348 28644 19412
rect 30420 19348 30484 19412
rect 29132 19272 29196 19276
rect 29132 19216 29182 19272
rect 29182 19216 29196 19272
rect 29132 19212 29196 19216
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 34652 19076 34716 19140
rect 38516 19076 38580 19140
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 29132 18668 29196 18732
rect 29500 18668 29564 18732
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 25268 17988 25332 18052
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 18460 17172 18524 17236
rect 28764 17036 28828 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 15148 16688 15212 16692
rect 15148 16632 15162 16688
rect 15162 16632 15212 16688
rect 15148 16628 15212 16632
rect 38516 16628 38580 16692
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 19012 15812 19076 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18828 15600 18892 15604
rect 18828 15544 18842 15600
rect 18842 15544 18892 15600
rect 18828 15540 18892 15544
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 18828 14648 18892 14652
rect 18828 14592 18842 14648
rect 18842 14592 18892 14648
rect 18828 14588 18892 14592
rect 19012 14180 19076 14244
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 15148 13636 15212 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 13860 13500 13924 13564
rect 14044 13288 14108 13292
rect 14044 13232 14058 13288
rect 14058 13232 14108 13288
rect 14044 13228 14108 13232
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 18460 13016 18524 13020
rect 18460 12960 18510 13016
rect 18510 12960 18524 13016
rect 18460 12956 18524 12960
rect 18460 12880 18524 12884
rect 18460 12824 18474 12880
rect 18474 12824 18524 12880
rect 18460 12820 18524 12824
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 34652 10644 34716 10708
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 13860 10100 13924 10164
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 14044 8876 14108 8940
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 18460 6700 18524 6764
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 15147 16692 15213 16693
rect 15147 16628 15148 16692
rect 15212 16628 15213 16692
rect 15147 16627 15213 16628
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 15150 13701 15210 16627
rect 17944 16352 18264 17376
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 27944 23968 28264 24528
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 28579 24172 28645 24173
rect 28579 24108 28580 24172
rect 28644 24108 28645 24172
rect 28579 24107 28645 24108
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 25267 22948 25333 22949
rect 25267 22884 25268 22948
rect 25332 22884 25333 22948
rect 25267 22883 25333 22884
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 25270 18053 25330 22883
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 28582 19413 28642 24107
rect 28947 23764 29013 23765
rect 28947 23700 28948 23764
rect 29012 23700 29013 23764
rect 28947 23699 29013 23700
rect 28579 19412 28645 19413
rect 28579 19348 28580 19412
rect 28644 19348 28645 19412
rect 28950 19350 29010 23699
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 30419 21316 30485 21317
rect 30419 21252 30420 21316
rect 30484 21252 30485 21316
rect 30419 21251 30485 21252
rect 29499 20908 29565 20909
rect 29499 20844 29500 20908
rect 29564 20844 29565 20908
rect 29499 20843 29565 20844
rect 28579 19347 28645 19348
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 25267 18052 25333 18053
rect 25267 17988 25268 18052
rect 25332 17988 25333 18052
rect 25267 17987 25333 17988
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 18459 17236 18525 17237
rect 18459 17172 18460 17236
rect 18524 17172 18525 17236
rect 18459 17171 18525 17172
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 15147 13700 15213 13701
rect 15147 13636 15148 13700
rect 15212 13636 15213 13700
rect 15147 13635 15213 13636
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 13859 13564 13925 13565
rect 13859 13500 13860 13564
rect 13924 13500 13925 13564
rect 13859 13499 13925 13500
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 13862 10165 13922 13499
rect 14043 13292 14109 13293
rect 14043 13228 14044 13292
rect 14108 13228 14109 13292
rect 14043 13227 14109 13228
rect 13859 10164 13925 10165
rect 13859 10100 13860 10164
rect 13924 10100 13925 10164
rect 13859 10099 13925 10100
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 14046 8941 14106 13227
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 18462 13021 18522 17171
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 19011 15876 19077 15877
rect 19011 15812 19012 15876
rect 19076 15812 19077 15876
rect 19011 15811 19077 15812
rect 18827 15604 18893 15605
rect 18827 15540 18828 15604
rect 18892 15540 18893 15604
rect 18827 15539 18893 15540
rect 18830 14653 18890 15539
rect 18827 14652 18893 14653
rect 18827 14588 18828 14652
rect 18892 14588 18893 14652
rect 18827 14587 18893 14588
rect 19014 14245 19074 15811
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 19011 14244 19077 14245
rect 19011 14180 19012 14244
rect 19076 14180 19077 14244
rect 19011 14179 19077 14180
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 18459 13020 18525 13021
rect 18459 12956 18460 13020
rect 18524 12956 18525 13020
rect 18459 12955 18525 12956
rect 18459 12884 18525 12885
rect 18459 12820 18460 12884
rect 18524 12820 18525 12884
rect 18459 12819 18525 12820
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 14043 8940 14109 8941
rect 14043 8876 14044 8940
rect 14108 8876 14109 8940
rect 14043 8875 14109 8876
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 18462 6765 18522 12819
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 18459 6764 18525 6765
rect 18459 6700 18460 6764
rect 18524 6700 18525 6764
rect 18459 6699 18525 6700
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 28766 19290 29010 19350
rect 28766 17101 28826 19290
rect 29131 19276 29197 19277
rect 29131 19212 29132 19276
rect 29196 19212 29197 19276
rect 29131 19211 29197 19212
rect 29134 18733 29194 19211
rect 29502 18733 29562 20843
rect 30422 19413 30482 21251
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 30419 19412 30485 19413
rect 30419 19348 30420 19412
rect 30484 19348 30485 19412
rect 30419 19347 30485 19348
rect 32944 19072 33264 20096
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 34651 19140 34717 19141
rect 34651 19076 34652 19140
rect 34716 19076 34717 19140
rect 34651 19075 34717 19076
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 29131 18732 29197 18733
rect 29131 18668 29132 18732
rect 29196 18668 29197 18732
rect 29131 18667 29197 18668
rect 29499 18732 29565 18733
rect 29499 18668 29500 18732
rect 29564 18668 29565 18732
rect 29499 18667 29565 18668
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 28763 17100 28829 17101
rect 28763 17036 28764 17100
rect 28828 17036 28829 17100
rect 28763 17035 28829 17036
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 34654 10709 34714 19075
rect 37944 18528 38264 19552
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 38515 19140 38581 19141
rect 38515 19076 38516 19140
rect 38580 19076 38581 19140
rect 38515 19075 38581 19076
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 38518 16693 38578 19075
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 38515 16692 38581 16693
rect 38515 16628 38516 16692
rect 38580 16628 38581 16692
rect 38515 16627 38581 16628
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 34651 10708 34717 10709
rect 34651 10644 34652 10708
rect 34716 10644 34717 10708
rect 34651 10643 34717 10644
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform -1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1679235063
transform -1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform -1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1679235063
transform -1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1679235063
transform -1 0 11224 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform -1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform -1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform -1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform -1 0 11224 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1679235063
transform -1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform -1 0 9476 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform -1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1679235063
transform -1 0 16376 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform -1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform -1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform -1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform -1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform -1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform -1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform -1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform -1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1679235063
transform -1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1679235063
transform -1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform -1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1679235063
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1679235063
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1679235063
transform -1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 37904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 37168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 37628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 44804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 39192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 44068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 39836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 40020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 45540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 39928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1679235063
transform -1 0 46184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1679235063
transform -1 0 46184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1679235063
transform -1 0 45908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1679235063
transform -1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1679235063
transform -1 0 5612 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4140 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1679235063
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1679235063
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1679235063
transform -1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1679235063
transform -1 0 2392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1679235063
transform -1 0 6808 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1679235063
transform -1 0 4232 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1679235063
transform -1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1679235063
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1679235063
transform -1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1679235063
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1679235063
transform -1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1679235063
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1679235063
transform 1 0 13892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1679235063
transform -1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1679235063
transform -1 0 7544 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1679235063
transform -1 0 23736 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1679235063
transform -1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1679235063
transform -1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1679235063
transform -1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1679235063
transform -1 0 21528 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1679235063
transform -1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1679235063
transform -1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1679235063
transform -1 0 21528 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1679235063
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1679235063
transform -1 0 17204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _195_
timestamp 1679235063
transform -1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1679235063
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1679235063
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1679235063
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1679235063
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1679235063
transform -1 0 21528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1679235063
transform -1 0 26680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 11408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform -1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1679235063
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1679235063
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1679235063
transform -1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1679235063
transform -1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform -1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1679235063
transform -1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1679235063
transform -1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1679235063
transform -1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1679235063
transform -1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1679235063
transform -1 0 9752 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1679235063
transform -1 0 11776 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1679235063
transform -1 0 11408 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1679235063
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1679235063
transform -1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1679235063
transform -1 0 10304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1679235063
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1679235063
transform -1 0 37076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1679235063
transform -1 0 38640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1679235063
transform 1 0 36800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1679235063
transform -1 0 39100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1679235063
transform -1 0 38180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform -1 0 39192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 37352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 37536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform -1 0 39376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform -1 0 40940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform -1 0 40020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform -1 0 40756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform -1 0 38916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform -1 0 40388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1679235063
transform -1 0 40756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform -1 0 40572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform -1 0 40664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1679235063
transform 1 0 5796 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1679235063
transform -1 0 26496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1679235063
transform -1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 19320 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 12880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform -1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 20516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform -1 0 16560 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S
timestamp 1679235063
transform -1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S
timestamp 1679235063
transform -1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform -1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S
timestamp 1679235063
transform -1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 16744 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform -1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 11960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform -1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 28060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform -1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform -1 0 22724 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 24656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 30360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform -1 0 37168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 35328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1679235063
transform -1 0 46092 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold11_A
timestamp 1679235063
transform -1 0 29716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold13_A
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold14_A
timestamp 1679235063
transform -1 0 32016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold16_A
timestamp 1679235063
transform -1 0 34960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold18_A
timestamp 1679235063
transform -1 0 32844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold20_A
timestamp 1679235063
transform -1 0 3404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold21_A
timestamp 1679235063
transform -1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold22_A
timestamp 1679235063
transform -1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold23_A
timestamp 1679235063
transform -1 0 46644 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold24_A
timestamp 1679235063
transform -1 0 47748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold25_A
timestamp 1679235063
transform -1 0 47748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold26_A
timestamp 1679235063
transform -1 0 46460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold27_A
timestamp 1679235063
transform -1 0 46920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold28_A
timestamp 1679235063
transform -1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold29_A
timestamp 1679235063
transform -1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold30_A
timestamp 1679235063
transform -1 0 47748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold31_A
timestamp 1679235063
transform -1 0 47932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold32_A
timestamp 1679235063
transform -1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold33_A
timestamp 1679235063
transform -1 0 47564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold34_A
timestamp 1679235063
transform -1 0 47748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold35_A
timestamp 1679235063
transform -1 0 44988 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold36_A
timestamp 1679235063
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold37_A
timestamp 1679235063
transform -1 0 3588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold38_A
timestamp 1679235063
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold39_A
timestamp 1679235063
transform -1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold40_A
timestamp 1679235063
transform -1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold41_A
timestamp 1679235063
transform -1 0 44528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold42_A
timestamp 1679235063
transform -1 0 3404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold43_A
timestamp 1679235063
transform -1 0 47472 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold44_A
timestamp 1679235063
transform -1 0 4140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold45_A
timestamp 1679235063
transform -1 0 47748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold46_A
timestamp 1679235063
transform -1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold47_A
timestamp 1679235063
transform -1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold48_A
timestamp 1679235063
transform -1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold49_A
timestamp 1679235063
transform -1 0 47104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold50_A
timestamp 1679235063
transform -1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold51_A
timestamp 1679235063
transform -1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold52_A
timestamp 1679235063
transform -1 0 45816 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold53_A
timestamp 1679235063
transform -1 0 48484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold54_A
timestamp 1679235063
transform -1 0 4140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold55_A
timestamp 1679235063
transform -1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold56_A
timestamp 1679235063
transform -1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold57_A
timestamp 1679235063
transform -1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold58_A
timestamp 1679235063
transform -1 0 4140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold59_A
timestamp 1679235063
transform -1 0 3588 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold60_A
timestamp 1679235063
transform -1 0 3404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold61_A
timestamp 1679235063
transform -1 0 37168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold62_A
timestamp 1679235063
transform 1 0 49036 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold65_A
timestamp 1679235063
transform -1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform -1 0 5336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform -1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform -1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform -1 0 4140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform -1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform -1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform -1 0 3588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform -1 0 3956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform -1 0 47748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform -1 0 47748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 47564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 47012 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform -1 0 46644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform -1 0 46828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform -1 0 46460 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform -1 0 47472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform -1 0 48208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 47564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform -1 0 27048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform -1 0 29716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform -1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform -1 0 34500 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform -1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform -1 0 42596 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform -1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform -1 0 43332 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform -1 0 47380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform -1 0 46276 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform -1 0 44068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform -1 0 9384 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform -1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform -1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1679235063
transform -1 0 44528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1679235063
transform -1 0 44252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform -1 0 46000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform -1 0 43700 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1679235063
transform -1 0 43884 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1679235063
transform -1 0 44344 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1679235063
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1679235063
transform -1 0 42596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1679235063
transform -1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1679235063
transform -1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1679235063
transform -1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1679235063
transform -1 0 31648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1679235063
transform -1 0 25300 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1679235063
transform -1 0 29164 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1679235063
transform -1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1679235063
transform -1 0 29348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1679235063
transform -1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1679235063
transform -1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1679235063
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1679235063
transform -1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1679235063
transform -1 0 49588 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1679235063
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1679235063
transform -1 0 48484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1679235063
transform -1 0 47748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1679235063
transform -1 0 48484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1679235063
transform 1 0 47196 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1679235063
transform -1 0 44896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1679235063
transform -1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 27048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 24472 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22080 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 17020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20516 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform -1 0 22172 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23184 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 27784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 30176 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 30728 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 27600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 28152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 34316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 34224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 36708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform -1 0 37076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 38456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 38456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform -1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 37444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 38640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 35880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 36064 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 36892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 33488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 34684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 33672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 34132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 28980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 30636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 32752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 32936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 30176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform -1 0 45908 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 43700 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 33304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 36892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 37628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 38456 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 39836 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 39468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 37076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 37260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 35512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 39468 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 41032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 40572 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 39376 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 40020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 40388 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 37076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 40204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 37260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 39192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 37444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 37444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 41124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 40020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 42044 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 40940 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 41032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 41492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 42044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 40020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 38916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 35880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 27416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21160 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 12328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform -1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 19596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform -1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__S
timestamp 1679235063
transform -1 0 31924 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 28336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 28152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 26036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 23460 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__S
timestamp 1679235063
transform -1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 30360 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 25852 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 27968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 30176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 27508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 25760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 22172 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 29440 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 25944 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26680 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 24288 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 30912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1
timestamp 1679235063
transform -1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1
timestamp 1679235063
transform -1 0 30544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 31188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 25576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1
timestamp 1679235063
transform -1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 30360 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 36064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 34316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__S
timestamp 1679235063
transform -1 0 34500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 27600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__S
timestamp 1679235063
transform -1 0 27968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform -1 0 34040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 29532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__S
timestamp 1679235063
transform -1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform -1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 37444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__S
timestamp 1679235063
transform -1 0 37076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1
timestamp 1679235063
transform -1 0 29440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__S
timestamp 1679235063
transform -1 0 31924 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__S
timestamp 1679235063
transform -1 0 35880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform -1 0 34592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 33948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 36616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 36800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 32752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__S
timestamp 1679235063
transform -1 0 33488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 34224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 34316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 34500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 34316 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 30452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__S
timestamp 1679235063
transform -1 0 32016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 26036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 31832 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 32292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 29440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 26036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0
timestamp 1679235063
transform -1 0 29072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 32016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 25668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 33764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 33304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 30268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 27784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 35696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 43332 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform -1 0 43148 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__S
timestamp 1679235063
transform -1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 28520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 39284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 41216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 44804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 31096 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 42596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 29716 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42412 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 42596 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 42780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform -1 0 33856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 34040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42596 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 42780 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 42228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 34224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1
timestamp 1679235063
transform -1 0 34592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 36892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 41308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 31740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 41032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 41216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1
timestamp 1679235063
transform -1 0 39192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 41584 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 41952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 36892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 41216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 41400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 36432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 38824 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 39008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1
timestamp 1679235063
transform -1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 28336 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 28612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 21712 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15640 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 19136 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12052 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 10488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0
timestamp 1679235063
transform -1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A1
timestamp 1679235063
transform -1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 20148 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16376 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 18216 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 18952 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 16192 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 16100 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 13616 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 15456 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10764 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9476 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform -1 0 12788 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 15180 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 12604 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform -1 0 11040 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 15272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform -1 0 16376 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform -1 0 16376 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform -1 0 16008 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17112 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform -1 0 16376 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform -1 0 17480 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform -1 0 18676 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform -1 0 11224 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform -1 0 13524 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 17940 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform -1 0 13800 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform -1 0 13524 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255
timestamp 1679235063
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 17112 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform -1 0 14720 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform -1 0 16008 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform -1 0 8556 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform -1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 14444 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 16744 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform -1 0 10212 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256
timestamp 1679235063
transform -1 0 11224 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform -1 0 12512 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform -1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform -1 0 12972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform -1 0 13800 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 15640 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 18308 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13156 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 14352 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257
timestamp 1679235063
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform -1 0 11868 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 29072 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23552 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 22724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform -1 0 27048 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform -1 0 23828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20976 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform -1 0 26128 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 23000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform -1 0 24104 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24196 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform -1 0 26496 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform -1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 18032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28888 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 28980 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 18952 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 17848 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 22448 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 22540 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform -1 0 18768 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform -1 0 23000 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 23276 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 28796 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform -1 0 29256 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 33304 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 34040 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 29900 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 30728 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform -1 0 35604 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform -1 0 35880 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1679235063
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42
timestamp 1679235063
transform 1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1679235063
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1679235063
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1679235063
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1679235063
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1679235063
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1679235063
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1679235063
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1679235063
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1679235063
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1679235063
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1679235063
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1679235063
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1679235063
transform 1 0 26036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1679235063
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1679235063
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1679235063
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1679235063
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1679235063
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1679235063
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_319
timestamp 1679235063
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_323
timestamp 1679235063
transform 1 0 30820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_332
timestamp 1679235063
transform 1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1679235063
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_345
timestamp 1679235063
transform 1 0 32844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1679235063
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1679235063
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_365
timestamp 1679235063
transform 1 0 34684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_368
timestamp 1679235063
transform 1 0 34960 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_378
timestamp 1679235063
transform 1 0 35880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1679235063
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_403
timestamp 1679235063
transform 1 0 38180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1679235063
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1679235063
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1679235063
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1679235063
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1679235063
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1679235063
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_459
timestamp 1679235063
transform 1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1679235063
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1679235063
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1679235063
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1679235063
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1679235063
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1679235063
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1679235063
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1679235063
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1679235063
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1679235063
transform 1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_35
timestamp 1679235063
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1679235063
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1679235063
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81
timestamp 1679235063
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1679235063
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1679235063
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1679235063
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_132
timestamp 1679235063
transform 1 0 13248 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1679235063
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1679235063
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_171
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1679235063
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1679235063
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1679235063
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1679235063
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1679235063
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1679235063
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_235
timestamp 1679235063
transform 1 0 22724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1679235063
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1679235063
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1679235063
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1679235063
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1679235063
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_301
timestamp 1679235063
transform 1 0 28796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_323
timestamp 1679235063
transform 1 0 30820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_330
timestamp 1679235063
transform 1 0 31464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1679235063
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1679235063
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1679235063
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1679235063
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_361
timestamp 1679235063
transform 1 0 34316 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_372
timestamp 1679235063
transform 1 0 35328 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1679235063
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1679235063
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1679235063
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1679235063
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1679235063
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1679235063
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1679235063
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1679235063
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1679235063
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1679235063
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1679235063
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1679235063
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1679235063
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1679235063
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1679235063
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_31
timestamp 1679235063
transform 1 0 3956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_43
timestamp 1679235063
transform 1 0 5060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_55
timestamp 1679235063
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_67
timestamp 1679235063
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1679235063
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1679235063
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_101
timestamp 1679235063
transform 1 0 10396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1679235063
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1679235063
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1679235063
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_180
timestamp 1679235063
transform 1 0 17664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1679235063
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_209
timestamp 1679235063
transform 1 0 20332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_236
timestamp 1679235063
transform 1 0 22816 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1679235063
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_261
timestamp 1679235063
transform 1 0 25116 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1679235063
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1679235063
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1679235063
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_311
timestamp 1679235063
transform 1 0 29716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_323
timestamp 1679235063
transform 1 0 30820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_335
timestamp 1679235063
transform 1 0 31924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_347
timestamp 1679235063
transform 1 0 33028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1679235063
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1679235063
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1679235063
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1679235063
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_387
timestamp 1679235063
transform 1 0 36708 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_391
timestamp 1679235063
transform 1 0 37076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1679235063
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1679235063
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1679235063
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1679235063
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1679235063
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1679235063
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1679235063
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1679235063
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1679235063
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_479
timestamp 1679235063
transform 1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_485
timestamp 1679235063
transform 1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1679235063
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1679235063
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1679235063
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1679235063
transform 1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_31
timestamp 1679235063
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_43
timestamp 1679235063
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1679235063
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1679235063
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1679235063
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_143
timestamp 1679235063
transform 1 0 14260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1679235063
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_175
timestamp 1679235063
transform 1 0 17204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_187
timestamp 1679235063
transform 1 0 18308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_199
timestamp 1679235063
transform 1 0 19412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_211
timestamp 1679235063
transform 1 0 20516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1679235063
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1679235063
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_233
timestamp 1679235063
transform 1 0 22540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_240
timestamp 1679235063
transform 1 0 23184 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_247
timestamp 1679235063
transform 1 0 23828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1679235063
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1679235063
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_289
timestamp 1679235063
transform 1 0 27692 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1679235063
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1679235063
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1679235063
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1679235063
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1679235063
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1679235063
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1679235063
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1679235063
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1679235063
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1679235063
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1679235063
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1679235063
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1679235063
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1679235063
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1679235063
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1679235063
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1679235063
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1679235063
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1679235063
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1679235063
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_507
timestamp 1679235063
transform 1 0 47748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1679235063
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1679235063
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1679235063
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1679235063
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_35
timestamp 1679235063
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_47
timestamp 1679235063
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_59
timestamp 1679235063
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_71
timestamp 1679235063
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1679235063
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1679235063
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1679235063
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1679235063
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_218
timestamp 1679235063
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_234
timestamp 1679235063
transform 1 0 22632 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1679235063
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1679235063
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_265
timestamp 1679235063
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_282
timestamp 1679235063
transform 1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_294
timestamp 1679235063
transform 1 0 28152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1679235063
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1679235063
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1679235063
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1679235063
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1679235063
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1679235063
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1679235063
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1679235063
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1679235063
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_385
timestamp 1679235063
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_390
timestamp 1679235063
transform 1 0 36984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1679235063
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_404
timestamp 1679235063
transform 1 0 38272 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_408
timestamp 1679235063
transform 1 0 38640 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1679235063
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1679235063
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1679235063
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1679235063
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1679235063
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1679235063
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1679235063
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_491
timestamp 1679235063
transform 1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_497
timestamp 1679235063
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1679235063
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1679235063
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1679235063
transform 1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1679235063
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1679235063
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_201
timestamp 1679235063
transform 1 0 19596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1679235063
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1679235063
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1679235063
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1679235063
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1679235063
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1679235063
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1679235063
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1679235063
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1679235063
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1679235063
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1679235063
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1679235063
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1679235063
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1679235063
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1679235063
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1679235063
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1679235063
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1679235063
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1679235063
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_395
timestamp 1679235063
transform 1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_401
timestamp 1679235063
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_409
timestamp 1679235063
transform 1 0 38732 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_413
timestamp 1679235063
transform 1 0 39100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_425
timestamp 1679235063
transform 1 0 40204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_437
timestamp 1679235063
transform 1 0 41308 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1679235063
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1679235063
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1679235063
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1679235063
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_485
timestamp 1679235063
transform 1 0 45724 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1679235063
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1679235063
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1679235063
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1679235063
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1679235063
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_35
timestamp 1679235063
transform 1 0 4324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_47
timestamp 1679235063
transform 1 0 5428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_59
timestamp 1679235063
transform 1 0 6532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_71
timestamp 1679235063
transform 1 0 7636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1679235063
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1679235063
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1679235063
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1679235063
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1679235063
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1679235063
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1679235063
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1679235063
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1679235063
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1679235063
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1679235063
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1679235063
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1679235063
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1679235063
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1679235063
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1679235063
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1679235063
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1679235063
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1679235063
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1679235063
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1679235063
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1679235063
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1679235063
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1679235063
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1679235063
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1679235063
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1679235063
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_461
timestamp 1679235063
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1679235063
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1679235063
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1679235063
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1679235063
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1679235063
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1679235063
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1679235063
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_21
timestamp 1679235063
transform 1 0 3036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_29
timestamp 1679235063
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1679235063
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1679235063
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1679235063
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_192
timestamp 1679235063
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1679235063
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1679235063
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1679235063
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1679235063
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1679235063
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1679235063
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1679235063
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1679235063
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1679235063
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1679235063
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1679235063
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1679235063
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1679235063
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1679235063
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1679235063
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1679235063
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1679235063
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1679235063
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1679235063
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1679235063
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_399
timestamp 1679235063
transform 1 0 37812 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_403
timestamp 1679235063
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1679235063
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1679235063
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1679235063
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1679235063
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1679235063
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1679235063
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_469
timestamp 1679235063
transform 1 0 44252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_481
timestamp 1679235063
transform 1 0 45356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_493
timestamp 1679235063
transform 1 0 46460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1679235063
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1679235063
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1679235063
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1679235063
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_21
timestamp 1679235063
transform 1 0 3036 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1679235063
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_34
timestamp 1679235063
transform 1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_38
timestamp 1679235063
transform 1 0 4600 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_50
timestamp 1679235063
transform 1 0 5704 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_62
timestamp 1679235063
transform 1 0 6808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1679235063
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1679235063
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1679235063
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_204
timestamp 1679235063
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_216
timestamp 1679235063
transform 1 0 20976 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_228
timestamp 1679235063
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_240
timestamp 1679235063
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1679235063
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1679235063
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1679235063
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1679235063
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1679235063
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1679235063
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1679235063
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1679235063
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1679235063
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1679235063
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1679235063
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1679235063
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1679235063
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1679235063
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1679235063
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1679235063
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1679235063
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1679235063
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1679235063
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1679235063
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1679235063
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1679235063
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1679235063
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1679235063
transform 1 0 47564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1679235063
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_13
timestamp 1679235063
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_25
timestamp 1679235063
transform 1 0 3404 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_31
timestamp 1679235063
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_43
timestamp 1679235063
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1679235063
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1679235063
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1679235063
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1679235063
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_193
timestamp 1679235063
transform 1 0 18860 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_196
timestamp 1679235063
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_208
timestamp 1679235063
transform 1 0 20240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1679235063
transform 1 0 20976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1679235063
transform 1 0 22816 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1679235063
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_252
timestamp 1679235063
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1679235063
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1679235063
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1679235063
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1679235063
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_317
timestamp 1679235063
transform 1 0 30268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1679235063
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_327
timestamp 1679235063
transform 1 0 31188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_333
timestamp 1679235063
transform 1 0 31740 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1679235063
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_342
timestamp 1679235063
transform 1 0 32568 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1679235063
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_358
timestamp 1679235063
transform 1 0 34040 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_370
timestamp 1679235063
transform 1 0 35144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1679235063
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1679235063
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1679235063
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_396
timestamp 1679235063
transform 1 0 37536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1679235063
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_410
timestamp 1679235063
transform 1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_414
timestamp 1679235063
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_426
timestamp 1679235063
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1679235063
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1679235063
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1679235063
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1679235063
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_473
timestamp 1679235063
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_479
timestamp 1679235063
transform 1 0 45172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_491
timestamp 1679235063
transform 1 0 46276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1679235063
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1679235063
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1679235063
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1679235063
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_21
timestamp 1679235063
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1679235063
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_160
timestamp 1679235063
transform 1 0 15824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1679235063
transform 1 0 16560 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1679235063
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_191
timestamp 1679235063
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1679235063
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_225
timestamp 1679235063
transform 1 0 21804 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_236
timestamp 1679235063
transform 1 0 22816 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1679235063
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1679235063
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1679235063
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1679235063
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1679235063
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1679235063
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1679235063
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_314
timestamp 1679235063
transform 1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_323
timestamp 1679235063
transform 1 0 30820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_334
timestamp 1679235063
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_338
timestamp 1679235063
transform 1 0 32200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_348
timestamp 1679235063
transform 1 0 33120 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_352
timestamp 1679235063
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1679235063
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1679235063
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1679235063
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_395
timestamp 1679235063
transform 1 0 37444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_398
timestamp 1679235063
transform 1 0 37720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_404
timestamp 1679235063
transform 1 0 38272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_412
timestamp 1679235063
transform 1 0 39008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1679235063
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1679235063
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1679235063
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1679235063
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1679235063
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1679235063
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1679235063
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1679235063
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1679235063
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1679235063
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1679235063
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_23
timestamp 1679235063
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1679235063
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1679235063
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1679235063
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_160
timestamp 1679235063
transform 1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_165
timestamp 1679235063
transform 1 0 16284 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1679235063
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1679235063
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_247
timestamp 1679235063
transform 1 0 23828 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_251
timestamp 1679235063
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1679235063
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1679235063
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1679235063
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1679235063
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1679235063
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1679235063
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1679235063
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1679235063
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_359
timestamp 1679235063
transform 1 0 34132 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_367
timestamp 1679235063
transform 1 0 34868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_379
timestamp 1679235063
transform 1 0 35972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1679235063
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1679235063
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1679235063
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_410
timestamp 1679235063
transform 1 0 38824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_414
timestamp 1679235063
transform 1 0 39192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_422
timestamp 1679235063
transform 1 0 39928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_429
timestamp 1679235063
transform 1 0 40572 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1679235063
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1679235063
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1679235063
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_461
timestamp 1679235063
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_471
timestamp 1679235063
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_483
timestamp 1679235063
transform 1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1679235063
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1679235063
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1679235063
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1679235063
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1679235063
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_33
timestamp 1679235063
transform 1 0 4140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_45
timestamp 1679235063
transform 1 0 5244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_57
timestamp 1679235063
transform 1 0 6348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_69
timestamp 1679235063
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1679235063
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1679235063
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1679235063
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1679235063
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1679235063
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_146
timestamp 1679235063
transform 1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1679235063
transform 1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_162
timestamp 1679235063
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1679235063
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1679235063
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1679235063
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1679235063
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_259
timestamp 1679235063
transform 1 0 24932 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_269
timestamp 1679235063
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_281
timestamp 1679235063
transform 1 0 26956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_289
timestamp 1679235063
transform 1 0 27692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_292
timestamp 1679235063
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1679235063
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1679235063
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1679235063
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_314
timestamp 1679235063
transform 1 0 29992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1679235063
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_342
timestamp 1679235063
transform 1 0 32568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_348
timestamp 1679235063
transform 1 0 33120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_359
timestamp 1679235063
transform 1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1679235063
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1679235063
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_376
timestamp 1679235063
transform 1 0 35696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_384
timestamp 1679235063
transform 1 0 36432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_388
timestamp 1679235063
transform 1 0 36800 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_396
timestamp 1679235063
transform 1 0 37536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_400
timestamp 1679235063
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_412
timestamp 1679235063
transform 1 0 39008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1679235063
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_423
timestamp 1679235063
transform 1 0 40020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_435
timestamp 1679235063
transform 1 0 41124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_447
timestamp 1679235063
transform 1 0 42228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_459
timestamp 1679235063
transform 1 0 43332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_471
timestamp 1679235063
transform 1 0 44436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1679235063
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1679235063
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1679235063
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1679235063
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1679235063
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1679235063
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1679235063
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1679235063
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_33
timestamp 1679235063
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1679235063
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1679235063
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1679235063
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1679235063
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1679235063
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1679235063
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1679235063
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1679235063
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1679235063
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1679235063
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1679235063
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1679235063
transform 1 0 22080 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1679235063
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_263
timestamp 1679235063
transform 1 0 25300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1679235063
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1679235063
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1679235063
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_331
timestamp 1679235063
transform 1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1679235063
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_339
timestamp 1679235063
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1679235063
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp 1679235063
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_376
timestamp 1679235063
transform 1 0 35696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1679235063
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1679235063
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1679235063
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1679235063
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1679235063
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1679235063
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1679235063
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1679235063
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1679235063
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1679235063
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1679235063
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1679235063
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1679235063
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1679235063
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1679235063
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1679235063
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1679235063
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_33
timestamp 1679235063
transform 1 0 4140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_45
timestamp 1679235063
transform 1 0 5244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_57
timestamp 1679235063
transform 1 0 6348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_69
timestamp 1679235063
transform 1 0 7452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1679235063
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1679235063
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1679235063
transform 1 0 12512 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 1679235063
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1679235063
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1679235063
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1679235063
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1679235063
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1679235063
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_243
timestamp 1679235063
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1679235063
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_275
timestamp 1679235063
transform 1 0 26404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_279
timestamp 1679235063
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_301
timestamp 1679235063
transform 1 0 28796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_305
timestamp 1679235063
transform 1 0 29164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1679235063
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1679235063
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1679235063
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_351
timestamp 1679235063
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1679235063
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1679235063
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_387
timestamp 1679235063
transform 1 0 36708 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_391
timestamp 1679235063
transform 1 0 37076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_407
timestamp 1679235063
transform 1 0 38548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_411
timestamp 1679235063
transform 1 0 38916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1679235063
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1679235063
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_427
timestamp 1679235063
transform 1 0 40388 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_431
timestamp 1679235063
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_443
timestamp 1679235063
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_455
timestamp 1679235063
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_467
timestamp 1679235063
transform 1 0 44068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1679235063
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1679235063
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1679235063
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1679235063
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1679235063
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_25
timestamp 1679235063
transform 1 0 3404 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1679235063
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1679235063
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1679235063
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1679235063
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1679235063
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1679235063
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1679235063
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1679235063
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1679235063
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_183
timestamp 1679235063
transform 1 0 17940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1679235063
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1679235063
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1679235063
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_267
timestamp 1679235063
transform 1 0 25668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_277
timestamp 1679235063
transform 1 0 26588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1679235063
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1679235063
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_296
timestamp 1679235063
transform 1 0 28336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_299
timestamp 1679235063
transform 1 0 28612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_312
timestamp 1679235063
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1679235063
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_332
timestamp 1679235063
transform 1 0 31648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1679235063
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_348
timestamp 1679235063
transform 1 0 33120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_352
timestamp 1679235063
transform 1 0 33488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1679235063
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1679235063
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_397
timestamp 1679235063
transform 1 0 37628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_409
timestamp 1679235063
transform 1 0 38732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_417
timestamp 1679235063
transform 1 0 39468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_423
timestamp 1679235063
transform 1 0 40020 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_427
timestamp 1679235063
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_439
timestamp 1679235063
transform 1 0 41492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1679235063
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1679235063
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1679235063
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1679235063
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1679235063
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1679235063
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1679235063
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1679235063
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1679235063
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1679235063
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_21
timestamp 1679235063
transform 1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_35
timestamp 1679235063
transform 1 0 4324 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_47
timestamp 1679235063
transform 1 0 5428 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_59
timestamp 1679235063
transform 1 0 6532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_71
timestamp 1679235063
transform 1 0 7636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1679235063
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1679235063
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1679235063
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1679235063
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1679235063
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_192
timestamp 1679235063
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1679235063
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1679235063
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1679235063
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1679235063
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1679235063
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_279
timestamp 1679235063
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_300
timestamp 1679235063
transform 1 0 28704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1679235063
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_320
timestamp 1679235063
transform 1 0 30544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_324
timestamp 1679235063
transform 1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1679235063
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1679235063
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_367
timestamp 1679235063
transform 1 0 34868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_375
timestamp 1679235063
transform 1 0 35604 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1679235063
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_406
timestamp 1679235063
transform 1 0 38456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_410
timestamp 1679235063
transform 1 0 38824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1679235063
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_427
timestamp 1679235063
transform 1 0 40388 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_434
timestamp 1679235063
transform 1 0 41032 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_446
timestamp 1679235063
transform 1 0 42136 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_458
timestamp 1679235063
transform 1 0 43240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 1679235063
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1679235063
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_487
timestamp 1679235063
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_499
timestamp 1679235063
transform 1 0 47012 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_507
timestamp 1679235063
transform 1 0 47748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1679235063
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1679235063
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_25
timestamp 1679235063
transform 1 0 3404 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1679235063
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1679235063
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1679235063
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1679235063
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_115
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1679235063
transform 1 0 12144 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1679235063
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1679235063
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1679235063
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1679235063
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_191
timestamp 1679235063
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_198
timestamp 1679235063
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1679235063
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1679235063
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1679235063
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_268
timestamp 1679235063
transform 1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_273
timestamp 1679235063
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1679235063
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1679235063
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1679235063
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_296
timestamp 1679235063
transform 1 0 28336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_318
timestamp 1679235063
transform 1 0 30360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_331
timestamp 1679235063
transform 1 0 31556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1679235063
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1679235063
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1679235063
transform 1 0 33120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_361
timestamp 1679235063
transform 1 0 34316 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_367
timestamp 1679235063
transform 1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1679235063
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1679235063
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_404
timestamp 1679235063
transform 1 0 38272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_417
timestamp 1679235063
transform 1 0 39468 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_425
timestamp 1679235063
transform 1 0 40204 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1679235063
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1679235063
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1679235063
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1679235063
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1679235063
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_473
timestamp 1679235063
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_481
timestamp 1679235063
transform 1 0 45356 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1679235063
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1679235063
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1679235063
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1679235063
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1679235063
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_111
timestamp 1679235063
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_164
timestamp 1679235063
transform 1 0 16192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_168
timestamp 1679235063
transform 1 0 16560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1679235063
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_208
timestamp 1679235063
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_213
timestamp 1679235063
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1679235063
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1679235063
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_275
timestamp 1679235063
transform 1 0 26404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_279
timestamp 1679235063
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1679235063
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_294
timestamp 1679235063
transform 1 0 28152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1679235063
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1679235063
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_331
timestamp 1679235063
transform 1 0 31556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_335
timestamp 1679235063
transform 1 0 31924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_357
timestamp 1679235063
transform 1 0 33948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1679235063
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1679235063
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1679235063
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_400
timestamp 1679235063
transform 1 0 37904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_413
timestamp 1679235063
transform 1 0 39100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1679235063
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1679235063
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_427
timestamp 1679235063
transform 1 0 40388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1679235063
transform 1 0 41032 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_441
timestamp 1679235063
transform 1 0 41676 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_453
timestamp 1679235063
transform 1 0 42780 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_465
timestamp 1679235063
transform 1 0 43884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1679235063
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1679235063
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_485
timestamp 1679235063
transform 1 0 45724 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_490
timestamp 1679235063
transform 1 0 46184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_502
timestamp 1679235063
transform 1 0 47288 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_508
timestamp 1679235063
transform 1 0 47840 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1679235063
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_9
timestamp 1679235063
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1679235063
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1679235063
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1679235063
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1679235063
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_105
timestamp 1679235063
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 1679235063
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1679235063
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_150
timestamp 1679235063
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1679235063
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1679235063
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1679235063
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1679235063
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_206
timestamp 1679235063
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1679235063
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1679235063
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1679235063
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1679235063
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_273
timestamp 1679235063
transform 1 0 26220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_277
timestamp 1679235063
transform 1 0 26588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1679235063
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_306
timestamp 1679235063
transform 1 0 29256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_311
timestamp 1679235063
transform 1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1679235063
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1679235063
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_348
timestamp 1679235063
transform 1 0 33120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_356
timestamp 1679235063
transform 1 0 33856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_369
timestamp 1679235063
transform 1 0 35052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_382
timestamp 1679235063
transform 1 0 36248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1679235063
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1679235063
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_426
timestamp 1679235063
transform 1 0 40296 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_430
timestamp 1679235063
transform 1 0 40664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_442
timestamp 1679235063
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1679235063
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1679235063
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1679235063
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_485
timestamp 1679235063
transform 1 0 45724 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_490
timestamp 1679235063
transform 1 0 46184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1679235063
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1679235063
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1679235063
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1679235063
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1679235063
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1679235063
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1679235063
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1679235063
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1679235063
transform 1 0 10580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1679235063
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_133
timestamp 1679235063
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1679235063
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1679235063
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1679235063
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1679235063
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1679235063
transform 1 0 19504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1679235063
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1679235063
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1679235063
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_256
timestamp 1679235063
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1679235063
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_274
timestamp 1679235063
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_280
timestamp 1679235063
transform 1 0 26864 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_292
timestamp 1679235063
transform 1 0 27968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_295
timestamp 1679235063
transform 1 0 28244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1679235063
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1679235063
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1679235063
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_324
timestamp 1679235063
transform 1 0 30912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1679235063
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_359
timestamp 1679235063
transform 1 0 34132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1679235063
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1679235063
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_376
timestamp 1679235063
transform 1 0 35696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_382
timestamp 1679235063
transform 1 0 36248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_404
timestamp 1679235063
transform 1 0 38272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_408
timestamp 1679235063
transform 1 0 38640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_416
timestamp 1679235063
transform 1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1679235063
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_433
timestamp 1679235063
transform 1 0 40940 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_440
timestamp 1679235063
transform 1 0 41584 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_452
timestamp 1679235063
transform 1 0 42688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_464
timestamp 1679235063
transform 1 0 43792 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1679235063
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1679235063
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_501
timestamp 1679235063
transform 1 0 47196 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_507
timestamp 1679235063
transform 1 0 47748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1679235063
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1679235063
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1679235063
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1679235063
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1679235063
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1679235063
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1679235063
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1679235063
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1679235063
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1679235063
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1679235063
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_128
timestamp 1679235063
transform 1 0 12880 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1679235063
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1679235063
transform 1 0 15364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1679235063
transform 1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_183
timestamp 1679235063
transform 1 0 17940 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1679235063
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1679235063
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1679235063
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1679235063
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1679235063
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1679235063
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1679235063
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1679235063
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1679235063
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1679235063
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_359
timestamp 1679235063
transform 1 0 34132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_372
timestamp 1679235063
transform 1 0 35328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_385
timestamp 1679235063
transform 1 0 36524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1679235063
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1679235063
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_404
timestamp 1679235063
transform 1 0 38272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_408
timestamp 1679235063
transform 1 0 38640 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_413
timestamp 1679235063
transform 1 0 39100 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_425
timestamp 1679235063
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1679235063
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1679235063
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1679235063
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1679235063
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_473
timestamp 1679235063
transform 1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_480
timestamp 1679235063
transform 1 0 45264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1679235063
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1679235063
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_507
timestamp 1679235063
transform 1 0 47748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_513
timestamp 1679235063
transform 1 0 48300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1679235063
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1679235063
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1679235063
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1679235063
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1679235063
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1679235063
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1679235063
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1679235063
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1679235063
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1679235063
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1679235063
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1679235063
transform 1 0 15640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1679235063
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1679235063
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1679235063
transform 1 0 17940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1679235063
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1679235063
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1679235063
transform 1 0 23000 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_242
timestamp 1679235063
transform 1 0 23368 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1679235063
transform 1 0 23644 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_257
timestamp 1679235063
transform 1 0 24748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1679235063
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1679235063
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1679235063
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1679235063
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1679235063
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1679235063
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1679235063
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_346
timestamp 1679235063
transform 1 0 32936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_359
timestamp 1679235063
transform 1 0 34132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1679235063
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1679235063
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1679235063
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_411
timestamp 1679235063
transform 1 0 38916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1679235063
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_425
timestamp 1679235063
transform 1 0 40204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_437
timestamp 1679235063
transform 1 0 41308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_449
timestamp 1679235063
transform 1 0 42412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_461
timestamp 1679235063
transform 1 0 43516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1679235063
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1679235063
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1679235063
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_501
timestamp 1679235063
transform 1 0 47196 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_507
timestamp 1679235063
transform 1 0 47748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_513
timestamp 1679235063
transform 1 0 48300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1679235063
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1679235063
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1679235063
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1679235063
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1679235063
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1679235063
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1679235063
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1679235063
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_99
timestamp 1679235063
transform 1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1679235063
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_126
timestamp 1679235063
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_130
timestamp 1679235063
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1679235063
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1679235063
transform 1 0 17664 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1679235063
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1679235063
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1679235063
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_229
timestamp 1679235063
transform 1 0 22172 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1679235063
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1679235063
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1679235063
transform 1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1679235063
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_289
timestamp 1679235063
transform 1 0 27692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_312
timestamp 1679235063
transform 1 0 29808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_325
timestamp 1679235063
transform 1 0 31004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_332
timestamp 1679235063
transform 1 0 31648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1679235063
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1679235063
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1679235063
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1679235063
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_387
timestamp 1679235063
transform 1 0 36708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1679235063
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1679235063
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1679235063
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_428
timestamp 1679235063
transform 1 0 40480 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_435
timestamp 1679235063
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1679235063
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1679235063
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1679235063
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1679235063
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1679235063
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1679235063
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1679235063
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_507
timestamp 1679235063
transform 1 0 47748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_513
timestamp 1679235063
transform 1 0 48300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1679235063
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1679235063
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1679235063
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1679235063
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_61
timestamp 1679235063
transform 1 0 6716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1679235063
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1679235063
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_87
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_99
timestamp 1679235063
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1679235063
transform 1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1679235063
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1679235063
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1679235063
transform 1 0 15456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1679235063
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_179
timestamp 1679235063
transform 1 0 17572 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_185
timestamp 1679235063
transform 1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_191
timestamp 1679235063
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_201
timestamp 1679235063
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1679235063
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_217
timestamp 1679235063
transform 1 0 21068 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1679235063
transform 1 0 21988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_231
timestamp 1679235063
transform 1 0 22356 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_248
timestamp 1679235063
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1679235063
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_278
timestamp 1679235063
transform 1 0 26680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_284
timestamp 1679235063
transform 1 0 27232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_295
timestamp 1679235063
transform 1 0 28244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_301
timestamp 1679235063
transform 1 0 28796 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1679235063
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_315
timestamp 1679235063
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_339
timestamp 1679235063
transform 1 0 32292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_352
timestamp 1679235063
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_359
timestamp 1679235063
transform 1 0 34132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1679235063
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1679235063
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_387
timestamp 1679235063
transform 1 0 36708 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1679235063
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1679235063
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1679235063
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_443
timestamp 1679235063
transform 1 0 41860 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_447
timestamp 1679235063
transform 1 0 42228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_459
timestamp 1679235063
transform 1 0 43332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1679235063
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1679235063
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1679235063
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1679235063
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_501
timestamp 1679235063
transform 1 0 47196 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_509
timestamp 1679235063
transform 1 0 47932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_512
timestamp 1679235063
transform 1 0 48208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_517
timestamp 1679235063
transform 1 0 48668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1679235063
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1679235063
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1679235063
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1679235063
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1679235063
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1679235063
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1679235063
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1679235063
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_91
timestamp 1679235063
transform 1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_99
timestamp 1679235063
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1679235063
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1679235063
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1679235063
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1679235063
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1679235063
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1679235063
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_186
timestamp 1679235063
transform 1 0 18216 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_194
timestamp 1679235063
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1679235063
transform 1 0 21068 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1679235063
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1679235063
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_237
timestamp 1679235063
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_248
timestamp 1679235063
transform 1 0 23920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 1679235063
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1679235063
transform 1 0 26404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1679235063
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1679235063
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1679235063
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1679235063
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_329
timestamp 1679235063
transform 1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1679235063
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1679235063
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1679235063
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1679235063
transform 1 0 34316 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_367
timestamp 1679235063
transform 1 0 34868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1679235063
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1679235063
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_398
timestamp 1679235063
transform 1 0 37720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_402
timestamp 1679235063
transform 1 0 38088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_423
timestamp 1679235063
transform 1 0 40020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_427
timestamp 1679235063
transform 1 0 40388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_437
timestamp 1679235063
transform 1 0 41308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1679235063
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1679235063
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1679235063
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1679235063
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1679235063
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1679235063
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1679235063
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1679235063
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1679235063
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_515
timestamp 1679235063
transform 1 0 48484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1679235063
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1679235063
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1679235063
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1679235063
transform 1 0 7636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1679235063
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_87
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_95
timestamp 1679235063
transform 1 0 9844 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1679235063
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1679235063
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1679235063
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1679235063
transform 1 0 12236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1679235063
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1679235063
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_171
timestamp 1679235063
transform 1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1679235063
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1679235063
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_213
timestamp 1679235063
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1679235063
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_240
timestamp 1679235063
transform 1 0 23184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1679235063
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_286
timestamp 1679235063
transform 1 0 27416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1679235063
transform 1 0 27784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_302
timestamp 1679235063
transform 1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1679235063
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_320
timestamp 1679235063
transform 1 0 30544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1679235063
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1679235063
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_358
timestamp 1679235063
transform 1 0 34040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1679235063
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_378
timestamp 1679235063
transform 1 0 35880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_391
timestamp 1679235063
transform 1 0 37076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_395
timestamp 1679235063
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1679235063
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1679235063
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_432
timestamp 1679235063
transform 1 0 40848 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_440
timestamp 1679235063
transform 1 0 41584 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_452
timestamp 1679235063
transform 1 0 42688 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_464
timestamp 1679235063
transform 1 0 43792 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1679235063
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1679235063
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_501
timestamp 1679235063
transform 1 0 47196 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_507
timestamp 1679235063
transform 1 0 47748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_513
timestamp 1679235063
transform 1 0 48300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1679235063
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1679235063
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1679235063
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1679235063
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1679235063
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1679235063
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1679235063
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1679235063
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1679235063
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1679235063
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1679235063
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1679235063
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1679235063
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1679235063
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1679235063
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1679235063
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1679235063
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1679235063
transform 1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1679235063
transform 1 0 18768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1679235063
transform 1 0 20976 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1679235063
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_228
timestamp 1679235063
transform 1 0 22080 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1679235063
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_267
timestamp 1679235063
transform 1 0 25668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1679235063
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1679235063
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1679235063
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1679235063
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1679235063
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_308
timestamp 1679235063
transform 1 0 29440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_321
timestamp 1679235063
transform 1 0 30636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1679235063
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1679235063
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1679235063
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1679235063
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_388
timestamp 1679235063
transform 1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1679235063
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_404
timestamp 1679235063
transform 1 0 38272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_408
timestamp 1679235063
transform 1 0 38640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_431
timestamp 1679235063
transform 1 0 40756 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_435
timestamp 1679235063
transform 1 0 41124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1679235063
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1679235063
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1679235063
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1679235063
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1679235063
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_497
timestamp 1679235063
transform 1 0 46828 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1679235063
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_507
timestamp 1679235063
transform 1 0 47748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_513
timestamp 1679235063
transform 1 0 48300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1679235063
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1679235063
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1679235063
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1679235063
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1679235063
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1679235063
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1679235063
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1679235063
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_127
timestamp 1679235063
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1679235063
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_163
timestamp 1679235063
transform 1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1679235063
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1679235063
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1679235063
transform 1 0 19688 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1679235063
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_232
timestamp 1679235063
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1679235063
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1679235063
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_271
timestamp 1679235063
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1679235063
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_281
timestamp 1679235063
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1679235063
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_311
timestamp 1679235063
transform 1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1679235063
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1679235063
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_341
timestamp 1679235063
transform 1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_353
timestamp 1679235063
transform 1 0 33580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_359
timestamp 1679235063
transform 1 0 34132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1679235063
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_370
timestamp 1679235063
transform 1 0 35144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_374
timestamp 1679235063
transform 1 0 35512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_397
timestamp 1679235063
transform 1 0 37628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_410
timestamp 1679235063
transform 1 0 38824 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1679235063
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1679235063
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_427
timestamp 1679235063
transform 1 0 40388 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_437
timestamp 1679235063
transform 1 0 41308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_449
timestamp 1679235063
transform 1 0 42412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_461
timestamp 1679235063
transform 1 0 43516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1679235063
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1679235063
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1679235063
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_501
timestamp 1679235063
transform 1 0 47196 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_507
timestamp 1679235063
transform 1 0 47748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_513
timestamp 1679235063
transform 1 0 48300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1679235063
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1679235063
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_32
timestamp 1679235063
transform 1 0 4048 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1679235063
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1679235063
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1679235063
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_75
timestamp 1679235063
transform 1 0 8004 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_87
timestamp 1679235063
transform 1 0 9108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_93
timestamp 1679235063
transform 1 0 9660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1679235063
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1679235063
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1679235063
transform 1 0 14720 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1679235063
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1679235063
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1679235063
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1679235063
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_192
timestamp 1679235063
transform 1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_196
timestamp 1679235063
transform 1 0 19136 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1679235063
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1679235063
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1679235063
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1679235063
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1679235063
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1679235063
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1679235063
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_305
timestamp 1679235063
transform 1 0 29164 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_313
timestamp 1679235063
transform 1 0 29900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_324
timestamp 1679235063
transform 1 0 30912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1679235063
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1679235063
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1679235063
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1679235063
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1679235063
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_373
timestamp 1679235063
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_377
timestamp 1679235063
transform 1 0 35788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_387
timestamp 1679235063
transform 1 0 36708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1679235063
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_399
timestamp 1679235063
transform 1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_421
timestamp 1679235063
transform 1 0 39836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_425
timestamp 1679235063
transform 1 0 40204 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_436
timestamp 1679235063
transform 1 0 41216 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1679235063
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1679235063
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1679235063
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1679235063
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_497
timestamp 1679235063
transform 1 0 46828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_501
timestamp 1679235063
transform 1 0 47196 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_507
timestamp 1679235063
transform 1 0 47748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_513
timestamp 1679235063
transform 1 0 48300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1679235063
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1679235063
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_47
timestamp 1679235063
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1679235063
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1679235063
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_75
timestamp 1679235063
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1679235063
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 1679235063
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1679235063
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1679235063
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1679235063
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_133
timestamp 1679235063
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_163
timestamp 1679235063
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1679235063
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1679235063
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1679235063
transform 1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1679235063
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1679235063
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_288
timestamp 1679235063
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_300
timestamp 1679235063
transform 1 0 28704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1679235063
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1679235063
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1679235063
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_328
timestamp 1679235063
transform 1 0 31280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1679235063
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_352
timestamp 1679235063
transform 1 0 33488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1679235063
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_371
timestamp 1679235063
transform 1 0 35236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_395
timestamp 1679235063
transform 1 0 37444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_399
timestamp 1679235063
transform 1 0 37812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_410
timestamp 1679235063
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1679235063
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_443
timestamp 1679235063
transform 1 0 41860 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_447
timestamp 1679235063
transform 1 0 42228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_459
timestamp 1679235063
transform 1 0 43332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1679235063
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1679235063
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1679235063
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_489
timestamp 1679235063
transform 1 0 46092 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_495
timestamp 1679235063
transform 1 0 46644 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_500
timestamp 1679235063
transform 1 0 47104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_505
timestamp 1679235063
transform 1 0 47564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_513
timestamp 1679235063
transform 1 0 48300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1679235063
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1679235063
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1679235063
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1679235063
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1679235063
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1679235063
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1679235063
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1679235063
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1679235063
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_116
timestamp 1679235063
transform 1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1679235063
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1679235063
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1679235063
transform 1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1679235063
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1679235063
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1679235063
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1679235063
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1679235063
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_242
timestamp 1679235063
transform 1 0 23368 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_263
timestamp 1679235063
transform 1 0 25300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_267
timestamp 1679235063
transform 1 0 25668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1679235063
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1679235063
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1679235063
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1679235063
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_310
timestamp 1679235063
transform 1 0 29624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_314
timestamp 1679235063
transform 1 0 29992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_320
timestamp 1679235063
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1679235063
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1679235063
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1679235063
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1679235063
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1679235063
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_387
timestamp 1679235063
transform 1 0 36708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1679235063
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_397
timestamp 1679235063
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1679235063
transform 1 0 39744 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_433
timestamp 1679235063
transform 1 0 40940 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_439
timestamp 1679235063
transform 1 0 41492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1679235063
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1679235063
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1679235063
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1679235063
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_485
timestamp 1679235063
transform 1 0 45724 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_497
timestamp 1679235063
transform 1 0 46828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1679235063
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_507
timestamp 1679235063
transform 1 0 47748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_513
timestamp 1679235063
transform 1 0 48300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1679235063
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1679235063
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1679235063
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1679235063
transform 1 0 7268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1679235063
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1679235063
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1679235063
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1679235063
transform 1 0 9476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_94
timestamp 1679235063
transform 1 0 9752 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1679235063
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1679235063
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1679235063
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1679235063
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1679235063
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1679235063
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1679235063
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_184
timestamp 1679235063
transform 1 0 18032 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1679235063
transform 1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1679235063
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1679235063
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_231
timestamp 1679235063
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_239
timestamp 1679235063
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1679235063
transform 1 0 24840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1679235063
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1679235063
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_288
timestamp 1679235063
transform 1 0 27600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_301
timestamp 1679235063
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_305
timestamp 1679235063
transform 1 0 29164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1679235063
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1679235063
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1679235063
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_346
timestamp 1679235063
transform 1 0 32936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_350
timestamp 1679235063
transform 1 0 33304 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_360
timestamp 1679235063
transform 1 0 34224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1679235063
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1679235063
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_389
timestamp 1679235063
transform 1 0 36892 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_397
timestamp 1679235063
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_408
timestamp 1679235063
transform 1 0 38640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_414
timestamp 1679235063
transform 1 0 39192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1679235063
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_432
timestamp 1679235063
transform 1 0 40848 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_438
timestamp 1679235063
transform 1 0 41400 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_450
timestamp 1679235063
transform 1 0 42504 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_462
timestamp 1679235063
transform 1 0 43608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1679235063
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_477
timestamp 1679235063
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_483
timestamp 1679235063
transform 1 0 45540 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_486
timestamp 1679235063
transform 1 0 45816 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_491
timestamp 1679235063
transform 1 0 46276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_498
timestamp 1679235063
transform 1 0 46920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_505
timestamp 1679235063
transform 1 0 47564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_513
timestamp 1679235063
transform 1 0 48300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1679235063
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1679235063
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1679235063
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1679235063
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_75
timestamp 1679235063
transform 1 0 8004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_83
timestamp 1679235063
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1679235063
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1679235063
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1679235063
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1679235063
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1679235063
transform 1 0 12788 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1679235063
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1679235063
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1679235063
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1679235063
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1679235063
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_199
timestamp 1679235063
transform 1 0 19412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1679235063
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1679235063
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1679235063
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_274
timestamp 1679235063
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1679235063
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1679235063
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1679235063
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1679235063
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_330
timestamp 1679235063
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1679235063
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_359
timestamp 1679235063
transform 1 0 34132 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_372
timestamp 1679235063
transform 1 0 35328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_378
timestamp 1679235063
transform 1 0 35880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1679235063
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_395
timestamp 1679235063
transform 1 0 37444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_418
timestamp 1679235063
transform 1 0 39560 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_431
timestamp 1679235063
transform 1 0 40756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_438
timestamp 1679235063
transform 1 0 41400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1679235063
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1679235063
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1679235063
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_473
timestamp 1679235063
transform 1 0 44620 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_477
timestamp 1679235063
transform 1 0 44988 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_482
timestamp 1679235063
transform 1 0 45448 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_489
timestamp 1679235063
transform 1 0 46092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_495
timestamp 1679235063
transform 1 0 46644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_502
timestamp 1679235063
transform 1 0 47288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_507
timestamp 1679235063
transform 1 0 47748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_513
timestamp 1679235063
transform 1 0 48300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1679235063
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1679235063
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1679235063
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1679235063
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 1679235063
transform 1 0 8096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1679235063
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_91
timestamp 1679235063
transform 1 0 9476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1679235063
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1679235063
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_112
timestamp 1679235063
transform 1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_120
timestamp 1679235063
transform 1 0 12144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1679235063
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_130
timestamp 1679235063
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1679235063
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1679235063
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_203
timestamp 1679235063
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1679235063
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_238
timestamp 1679235063
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_246
timestamp 1679235063
transform 1 0 23736 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_258
timestamp 1679235063
transform 1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_276
timestamp 1679235063
transform 1 0 26496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_282
timestamp 1679235063
transform 1 0 27048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_287
timestamp 1679235063
transform 1 0 27508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1679235063
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1679235063
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1679235063
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_314
timestamp 1679235063
transform 1 0 29992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_320
timestamp 1679235063
transform 1 0 30544 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_332
timestamp 1679235063
transform 1 0 31648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_336
timestamp 1679235063
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_340
timestamp 1679235063
transform 1 0 32384 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1679235063
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1679235063
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_387
timestamp 1679235063
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_395
timestamp 1679235063
transform 1 0 37444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1679235063
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1679235063
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1679235063
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_445
timestamp 1679235063
transform 1 0 42044 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_455
timestamp 1679235063
transform 1 0 42964 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_461
timestamp 1679235063
transform 1 0 43516 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_469
timestamp 1679235063
transform 1 0 44252 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_477
timestamp 1679235063
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_482
timestamp 1679235063
transform 1 0 45448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_489
timestamp 1679235063
transform 1 0 46092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_497
timestamp 1679235063
transform 1 0 46828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_505
timestamp 1679235063
transform 1 0 47564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_513
timestamp 1679235063
transform 1 0 48300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1679235063
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_41
timestamp 1679235063
transform 1 0 4876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1679235063
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1679235063
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1679235063
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_95
timestamp 1679235063
transform 1 0 9844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_100
timestamp 1679235063
transform 1 0 10304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_105
timestamp 1679235063
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1679235063
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_124
timestamp 1679235063
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1679235063
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1679235063
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_138
timestamp 1679235063
transform 1 0 13800 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1679235063
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1679235063
transform 1 0 17204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1679235063
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1679235063
transform 1 0 20424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1679235063
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1679235063
transform 1 0 22264 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1679235063
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_266
timestamp 1679235063
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_272
timestamp 1679235063
transform 1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1679235063
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1679235063
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1679235063
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1679235063
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1679235063
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_331
timestamp 1679235063
transform 1 0 31556 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1679235063
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1679235063
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1679235063
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_345
timestamp 1679235063
transform 1 0 32844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_358
timestamp 1679235063
transform 1 0 34040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_371
timestamp 1679235063
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_375
timestamp 1679235063
transform 1 0 35604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_385
timestamp 1679235063
transform 1 0 36524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1679235063
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_399
timestamp 1679235063
transform 1 0 37812 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_421
timestamp 1679235063
transform 1 0 39836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_431
timestamp 1679235063
transform 1 0 40756 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_434
timestamp 1679235063
transform 1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1679235063
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1679235063
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_454
timestamp 1679235063
transform 1 0 42872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_461
timestamp 1679235063
transform 1 0 43516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_475
timestamp 1679235063
transform 1 0 44804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_479
timestamp 1679235063
transform 1 0 45172 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_484
timestamp 1679235063
transform 1 0 45632 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_488
timestamp 1679235063
transform 1 0 46000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_494
timestamp 1679235063
transform 1 0 46552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1679235063
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1679235063
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_511
timestamp 1679235063
transform 1 0 48116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_515
timestamp 1679235063
transform 1 0 48484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1679235063
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1679235063
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1679235063
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1679235063
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_103
timestamp 1679235063
transform 1 0 10580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_107
timestamp 1679235063
transform 1 0 10948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1679235063
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1679235063
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1679235063
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1679235063
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1679235063
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1679235063
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_243
timestamp 1679235063
transform 1 0 23460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_268
timestamp 1679235063
transform 1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_279
timestamp 1679235063
transform 1 0 26772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1679235063
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1679235063
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1679235063
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_314
timestamp 1679235063
transform 1 0 29992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_320
timestamp 1679235063
transform 1 0 30544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1679235063
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_356
timestamp 1679235063
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1679235063
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_376
timestamp 1679235063
transform 1 0 35696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1679235063
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_414
timestamp 1679235063
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_423
timestamp 1679235063
transform 1 0 40020 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_434
timestamp 1679235063
transform 1 0 41032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_447
timestamp 1679235063
transform 1 0 42228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_453
timestamp 1679235063
transform 1 0 42780 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_466
timestamp 1679235063
transform 1 0 43976 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1679235063
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_489
timestamp 1679235063
transform 1 0 46092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_497
timestamp 1679235063
transform 1 0 46828 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_503
timestamp 1679235063
transform 1 0 47380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_513
timestamp 1679235063
transform 1 0 48300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1679235063
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1679235063
transform 1 0 3036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_29
timestamp 1679235063
transform 1 0 3772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_63
timestamp 1679235063
transform 1 0 6900 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_67
timestamp 1679235063
transform 1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_85
timestamp 1679235063
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1679235063
transform 1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_119
timestamp 1679235063
transform 1 0 12052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1679235063
transform 1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_141
timestamp 1679235063
transform 1 0 14076 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1679235063
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1679235063
transform 1 0 19228 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_220
timestamp 1679235063
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1679235063
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_256
timestamp 1679235063
transform 1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1679235063
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1679235063
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_286
timestamp 1679235063
transform 1 0 27416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_290
timestamp 1679235063
transform 1 0 27784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1679235063
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1679235063
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1679235063
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1679235063
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_348
timestamp 1679235063
transform 1 0 33120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_352
timestamp 1679235063
transform 1 0 33488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_374
timestamp 1679235063
transform 1 0 35512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_378
timestamp 1679235063
transform 1 0 35880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1679235063
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1679235063
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_415
timestamp 1679235063
transform 1 0 39284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_421
timestamp 1679235063
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_432
timestamp 1679235063
transform 1 0 40848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_439
timestamp 1679235063
transform 1 0 41492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1679235063
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1679235063
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_459
timestamp 1679235063
transform 1 0 43332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_473
timestamp 1679235063
transform 1 0 44620 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_481
timestamp 1679235063
transform 1 0 45356 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_489
timestamp 1679235063
transform 1 0 46092 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_493
timestamp 1679235063
transform 1 0 46460 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1679235063
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_505
timestamp 1679235063
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1679235063
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_515
timestamp 1679235063
transform 1 0 48484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1679235063
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1679235063
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1679235063
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1679235063
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1679235063
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1679235063
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_98
timestamp 1679235063
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1679235063
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1679235063
transform 1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1679235063
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_199
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1679235063
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1679235063
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1679235063
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_259
timestamp 1679235063
transform 1 0 24932 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_265
timestamp 1679235063
transform 1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1679235063
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_300
timestamp 1679235063
transform 1 0 28704 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1679235063
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_320
timestamp 1679235063
transform 1 0 30544 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_324
timestamp 1679235063
transform 1 0 30912 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_327
timestamp 1679235063
transform 1 0 31188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_350
timestamp 1679235063
transform 1 0 33304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_357
timestamp 1679235063
transform 1 0 33948 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1679235063
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_367
timestamp 1679235063
transform 1 0 34868 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_389
timestamp 1679235063
transform 1 0 36892 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_413
timestamp 1679235063
transform 1 0 39100 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1679235063
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1679235063
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_432
timestamp 1679235063
transform 1 0 40848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_436
timestamp 1679235063
transform 1 0 41216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_462
timestamp 1679235063
transform 1 0 43608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1679235063
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1679235063
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_483
timestamp 1679235063
transform 1 0 45540 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_491
timestamp 1679235063
transform 1 0 46276 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_501
timestamp 1679235063
transform 1 0 47196 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_513
timestamp 1679235063
transform 1 0 48300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1679235063
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_63
timestamp 1679235063
transform 1 0 6900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1679235063
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1679235063
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1679235063
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_212
timestamp 1679235063
transform 1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_217
timestamp 1679235063
transform 1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1679235063
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_250
timestamp 1679235063
transform 1 0 24104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_256
timestamp 1679235063
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1679235063
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1679235063
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1679235063
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1679235063
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_300
timestamp 1679235063
transform 1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_307
timestamp 1679235063
transform 1 0 29348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_311
timestamp 1679235063
transform 1 0 29716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1679235063
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1679235063
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_348
timestamp 1679235063
transform 1 0 33120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_352
timestamp 1679235063
transform 1 0 33488 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_373
timestamp 1679235063
transform 1 0 35420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_377
timestamp 1679235063
transform 1 0 35788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_387
timestamp 1679235063
transform 1 0 36708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1679235063
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1679235063
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_404
timestamp 1679235063
transform 1 0 38272 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_408
timestamp 1679235063
transform 1 0 38640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_419
timestamp 1679235063
transform 1 0 39652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_423
timestamp 1679235063
transform 1 0 40020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1679235063
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_463
timestamp 1679235063
transform 1 0 43700 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_469
timestamp 1679235063
transform 1 0 44252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_476
timestamp 1679235063
transform 1 0 44896 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_488
timestamp 1679235063
transform 1 0 46000 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1679235063
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_509
timestamp 1679235063
transform 1 0 47932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_519
timestamp 1679235063
transform 1 0 48852 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1679235063
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1679235063
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1679235063
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1679235063
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_272
timestamp 1679235063
transform 1 0 26128 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1679235063
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_287
timestamp 1679235063
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1679235063
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_301
timestamp 1679235063
transform 1 0 28796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1679235063
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1679235063
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1679235063
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1679235063
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1679235063
transform 1 0 31280 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1679235063
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1679235063
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_349
timestamp 1679235063
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1679235063
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1679235063
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1679235063
transform 1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_389
timestamp 1679235063
transform 1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1679235063
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1679235063
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_411
timestamp 1679235063
transform 1 0 38916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1679235063
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1679235063
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_432
timestamp 1679235063
transform 1 0 40848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_436
timestamp 1679235063
transform 1 0 41216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_446
timestamp 1679235063
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1679235063
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_454
timestamp 1679235063
transform 1 0 42872 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_461
timestamp 1679235063
transform 1 0 43516 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_465
timestamp 1679235063
transform 1 0 43884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_471
timestamp 1679235063
transform 1 0 44436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1679235063
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1679235063
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_487
timestamp 1679235063
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1679235063
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1679235063
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_507
timestamp 1679235063
transform 1 0 47748 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_513
timestamp 1679235063
transform 1 0 48300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_521
timestamp 1679235063
transform 1 0 49036 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 42596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold2
timestamp 1679235063
transform 1 0 44620 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform -1 0 42136 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 45172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 43976 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold6
timestamp 1679235063
transform -1 0 42136 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 47564 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform -1 0 46000 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 12328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 29716 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold12 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 17664 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 2852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 30912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold15
timestamp 1679235063
transform -1 0 16376 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold17
timestamp 1679235063
transform -1 0 15824 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 33028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold19
timestamp 1679235063
transform -1 0 15824 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 2668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 1564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform -1 0 47012 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform -1 0 49404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform -1 0 49404 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform -1 0 49404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform -1 0 49404 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform -1 0 49404 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform -1 0 49404 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform -1 0 3404 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform -1 0 49404 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform -1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform -1 0 49404 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform -1 0 49404 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform -1 0 49404 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform -1 0 48300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 2668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 1564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform -1 0 3404 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform -1 0 49404 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform -1 0 49404 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 1564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform -1 0 49404 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 1564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform -1 0 49404 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform -1 0 3404 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform -1 0 49404 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 1564 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform -1 0 49404 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 1564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 1564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 1564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 1564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 1564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 1564 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 37444 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform -1 0 47288 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold63 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform -1 0 48852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 46368 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 9660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform -1 0 10764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform -1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform -1 0 46276 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1679235063
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform -1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1679235063
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1679235063
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1679235063
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1679235063
transform -1 0 2484 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1679235063
transform -1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1679235063
transform 1 0 2852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1679235063
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1679235063
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform -1 0 2484 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1679235063
transform -1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1679235063
transform 1 0 3772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1679235063
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform -1 0 4048 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1679235063
transform -1 0 2484 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1679235063
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform -1 0 3128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1679235063
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1679235063
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1679235063
transform -1 0 2484 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1679235063
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1679235063
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1679235063
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1679235063
transform -1 0 2484 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1679235063
transform 1 0 2852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 47012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1679235063
transform -1 0 48300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1679235063
transform -1 0 48300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 47288 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1679235063
transform -1 0 48300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1679235063
transform -1 0 48300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1679235063
transform -1 0 48300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 47012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1679235063
transform -1 0 48300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1679235063
transform -1 0 47288 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1679235063
transform -1 0 47288 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1679235063
transform -1 0 48300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 46644 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1679235063
transform -1 0 47564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1679235063
transform -1 0 46828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1679235063
transform -1 0 46828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 45816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1679235063
transform 1 0 45816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1679235063
transform -1 0 48300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 47288 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 45172 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1679235063
transform 1 0 43976 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1679235063
transform -1 0 48300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1679235063
transform -1 0 48300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 48392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1679235063
transform -1 0 49404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1679235063
transform -1 0 48300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1679235063
transform -1 0 48300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 47012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1679235063
transform -1 0 48300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform -1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1679235063
transform -1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1679235063
transform -1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1679235063
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1679235063
transform 1 0 38640 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1679235063
transform 1 0 33672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1679235063
transform 1 0 39284 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1679235063
transform 1 0 43240 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1679235063
transform 1 0 42596 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1679235063
transform 1 0 43240 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1679235063
transform -1 0 11960 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1679235063
transform 1 0 43700 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1679235063
transform 1 0 41216 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1679235063
transform 1 0 43056 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1679235063
transform 1 0 43884 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1679235063
transform 1 0 45172 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1679235063
transform 1 0 41216 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1679235063
transform 1 0 43240 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1679235063
transform 1 0 41860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1679235063
transform 1 0 45172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1679235063
transform 1 0 42596 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1679235063
transform -1 0 12696 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1679235063
transform -1 0 22908 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1679235063
transform -1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1679235063
transform -1 0 30636 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1679235063
transform -1 0 24104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1679235063
transform -1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1679235063
transform -1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1679235063
transform -1 0 28796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1679235063
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1679235063
transform 1 0 31188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1679235063
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1679235063
transform 1 0 35052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97
timestamp 1679235063
transform -1 0 38364 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1679235063
transform 1 0 44160 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1679235063
transform 1 0 43516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1679235063
transform -1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1679235063
transform -1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1679235063
transform -1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1679235063
transform -1 0 49036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1679235063
transform -1 0 48116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1679235063
transform -1 0 48116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1679235063
transform -1 0 46092 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1679235063
transform -1 0 46552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1679235063
transform -1 0 45632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1679235063
transform -1 0 45356 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1679235063
transform -1 0 45540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 40664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform -1 0 4876 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform -1 0 3036 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform -1 0 3036 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform -1 0 3036 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform -1 0 3036 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform -1 0 3036 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform -1 0 3036 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform -1 0 3036 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform -1 0 4876 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform -1 0 3036 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform -1 0 3036 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform -1 0 3036 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform -1 0 3036 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform -1 0 5428 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform -1 0 5428 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform -1 0 7268 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform -1 0 7268 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform -1 0 5428 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform -1 0 7268 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform -1 0 3036 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform -1 0 3036 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform -1 0 3036 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform -1 0 3036 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform -1 0 3036 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform -1 0 3036 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform -1 0 3036 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform -1 0 3036 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 45816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 46092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1679235063
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1679235063
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1679235063
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1679235063
transform 1 0 43976 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1679235063
transform 1 0 46092 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1679235063
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1679235063
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1679235063
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1679235063
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1679235063
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1679235063
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1679235063
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1679235063
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1679235063
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1679235063
transform 1 0 45816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1679235063
transform 1 0 45816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1679235063
transform 1 0 46092 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1679235063
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1679235063
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1679235063
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1679235063
transform 1 0 45816 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1679235063
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1679235063
transform -1 0 5428 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1679235063
transform -1 0 9384 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1679235063
transform -1 0 11224 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1679235063
transform -1 0 11224 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1679235063
transform -1 0 11960 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1679235063
transform -1 0 11224 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1679235063
transform -1 0 14076 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1679235063
transform -1 0 13800 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1679235063
transform -1 0 13800 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1679235063
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1679235063
transform -1 0 4876 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1679235063
transform -1 0 16376 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1679235063
transform -1 0 16744 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1679235063
transform -1 0 16376 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1679235063
transform -1 0 18860 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1679235063
transform -1 0 16376 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1679235063
transform -1 0 18400 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1679235063
transform -1 0 18952 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1679235063
transform -1 0 21528 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1679235063
transform -1 0 3496 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1679235063
transform -1 0 4232 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1679235063
transform -1 0 6072 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1679235063
transform 1 0 7452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1679235063
transform -1 0 13248 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1679235063
transform -1 0 13800 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1679235063
transform -1 0 18308 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1679235063
transform -1 0 19596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1679235063
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1679235063
transform 1 0 22356 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1679235063
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 29256 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 26404 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 24472 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 24104 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 22356 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17020 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18584 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 18952 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19136 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 23828 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21068 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 22816 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 20976 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19596 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 21528 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 18952 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 22172 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 20608 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23828 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 25300 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25760 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 28888 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 27416 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 29900 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 26680 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25668 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 26680 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 23000 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28336 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 30452 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 32292 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 32200 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 34868 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 36984 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37444 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 35144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 37812 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 33856 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 35696 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 29992 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32108 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 32936 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27968 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 29716 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 30360 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 26956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 28796 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 32200 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 31096 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 32568 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 29716 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 29348 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 26864 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 43608 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 30820 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 31832 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 31372 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 33672 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 35420 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 35052 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 36708 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 34132 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 32476 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 39284 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 39100 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 39192 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 37996 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 39468 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 39560 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 37628 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 33580 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 35604 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 39744 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 39836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 41860 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 40756 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 39560 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 38180 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 40020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 39560 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 38916 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform -1 0 34132 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 31188 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 27416 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 26680 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 25668 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 26404 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 25300 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 24104 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 23828 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 21528 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 21252 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 21252 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 22080 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 22264 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 18676 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 14904 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12972 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 16100 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 14536 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform -1 0 13524 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 12420 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 16100 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 17020 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform -1 0 18952 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 27232 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1679235063
transform -1 0 23460 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__258
timestamp 1679235063
transform 1 0 26036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1679235063
transform -1 0 21712 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1679235063
transform -1 0 23920 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19872 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__211
timestamp 1679235063
transform -1 0 15732 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1679235063
transform -1 0 17572 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__214
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1679235063
transform 1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24656 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1679235063
transform -1 0 20332 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23092 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1679235063
transform -1 0 20516 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__216
timestamp 1679235063
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19872 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27968 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20884 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__259
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1679235063
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17940 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1679235063
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21436 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__260
timestamp 1679235063
transform -1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1679235063
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27876 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1679235063
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__261
timestamp 1679235063
transform -1 0 17112 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1679235063
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9660 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1679235063
transform 1 0 26772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1679235063
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__262
timestamp 1679235063
transform -1 0 22908 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1679235063
transform 1 0 28336 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__212
timestamp 1679235063
transform 1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1679235063
transform -1 0 24104 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 28336 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28336 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__213
timestamp 1679235063
transform -1 0 27968 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11132 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22632 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__215
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19964 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform -1 0 30268 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 33304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1679235063
transform -1 0 28612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform -1 0 31832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__217
timestamp 1679235063
transform -1 0 30084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform -1 0 31740 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform -1 0 34316 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 39560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform -1 0 34040 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform -1 0 33120 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1679235063
transform -1 0 30544 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform -1 0 36708 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__220
timestamp 1679235063
transform 1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform -1 0 34316 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform -1 0 38824 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 41124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform -1 0 35236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1679235063
transform -1 0 30544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform -1 0 36800 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform -1 0 36524 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__224
timestamp 1679235063
transform -1 0 31832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform -1 0 38272 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 41584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform -1 0 35696 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform -1 0 33580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1679235063
transform -1 0 36248 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__227
timestamp 1679235063
transform 1 0 33764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1679235063
transform -1 0 33120 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform -1 0 36708 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 38640 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform -1 0 39100 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 41676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform -1 0 34224 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform -1 0 33488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1679235063
transform -1 0 34132 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1679235063
transform -1 0 31832 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__218
timestamp 1679235063
transform -1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform -1 0 35328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform -1 0 36892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform -1 0 38272 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 41032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform -1 0 33120 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1679235063
transform -1 0 33120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1679235063
transform -1 0 27968 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform -1 0 34132 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1679235063
transform -1 0 33120 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__219
timestamp 1679235063
transform -1 0 29992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1679235063
transform -1 0 37904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 41032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1679235063
transform -1 0 30636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1679235063
transform -1 0 27968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform -1 0 31372 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__221
timestamp 1679235063
transform 1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1679235063
transform -1 0 29256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1679235063
transform -1 0 34316 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 38456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform -1 0 30544 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 30176 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1679235063
transform -1 0 26496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform -1 0 30544 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1679235063
transform -1 0 31004 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__222
timestamp 1679235063
transform -1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1679235063
transform -1 0 33396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 37904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform -1 0 32108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1679235063
transform -1 0 32936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform -1 0 33120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1679235063
transform -1 0 31832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__223
timestamp 1679235063
transform 1 0 32292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1679235063
transform -1 0 35696 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 39192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform -1 0 30544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__225
timestamp 1679235063
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1679235063
transform -1 0 28980 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform -1 0 33396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 37720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform -1 0 29440 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1679235063
transform -1 0 27784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__226
timestamp 1679235063
transform -1 0 26680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform -1 0 33120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 36800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform -1 0 35696 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 38824 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1679235063
transform -1 0 24104 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__228
timestamp 1679235063
transform 1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 28428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 35880 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform -1 0 29164 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 27140 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform -1 0 35696 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40020 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1679235063
transform -1 0 31740 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 33028 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__234
timestamp 1679235063
transform -1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 28428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform -1 0 35328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40020 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 35696 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__244
timestamp 1679235063
transform 1 0 31280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform -1 0 30912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 30820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 40204 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 41400 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1679235063
transform -1 0 33488 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40020 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 36064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__252
timestamp 1679235063
transform -1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform -1 0 38272 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 41216 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1679235063
transform -1 0 34316 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1679235063
transform -1 0 36892 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__253
timestamp 1679235063
transform 1 0 41124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 36064 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 31464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform -1 0 35512 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40112 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform -1 0 31740 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__229
timestamp 1679235063
transform 1 0 31372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 31464 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform -1 0 40848 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__230
timestamp 1679235063
transform -1 0 35144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 36064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform -1 0 40756 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40480 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__231
timestamp 1679235063
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1679235063
transform -1 0 35512 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1679235063
transform 1 0 37996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform -1 0 40848 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__232
timestamp 1679235063
transform 1 0 37076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1679235063
transform -1 0 35696 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1679235063
transform 1 0 35880 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform -1 0 38640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 39652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1679235063
transform -1 0 31556 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__233
timestamp 1679235063
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 25760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27324 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__235
timestamp 1679235063
transform -1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1679235063
transform -1 0 25668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__236
timestamp 1679235063
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22908 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1679235063
transform -1 0 22908 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__237
timestamp 1679235063
transform -1 0 20056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__238
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24196 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22080 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22264 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__239
timestamp 1679235063
transform 1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__240
timestamp 1679235063
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__241
timestamp 1679235063
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 12604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__242
timestamp 1679235063
transform -1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__243
timestamp 1679235063
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform -1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__245
timestamp 1679235063
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16744 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__246
timestamp 1679235063
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13892 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__247
timestamp 1679235063
transform -1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__248
timestamp 1679235063
transform -1 0 9936 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__249
timestamp 1679235063
transform -1 0 10764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__250
timestamp 1679235063
transform -1 0 10120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__251
timestamp 1679235063
transform -1 0 10120 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 26200 49294 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 26200 1638 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 13608 51000 13728 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 17688 51000 17808 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 18096 51000 18216 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 18912 51000 19032 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 19320 51000 19440 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 19728 51000 19848 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 20136 51000 20256 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 21360 51000 21480 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 14016 51000 14136 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 21768 51000 21888 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 22176 51000 22296 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 22992 51000 23112 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 23400 51000 23520 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 24216 51000 24336 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 25032 51000 25152 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 25440 51000 25560 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 14832 51000 14952 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 15240 51000 15360 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 15648 51000 15768 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 16056 51000 16176 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 16872 51000 16992 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 17280 51000 17400 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 1368 51000 1488 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 5448 51000 5568 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 5856 51000 5976 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 6672 51000 6792 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 7080 51000 7200 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 7488 51000 7608 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 7896 51000 8016 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 8712 51000 8832 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 9120 51000 9240 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 1776 51000 1896 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 9528 51000 9648 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 9936 51000 10056 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 10752 51000 10872 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 11160 51000 11280 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 11568 51000 11688 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 11976 51000 12096 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 12792 51000 12912 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 13200 51000 13320 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 2184 51000 2304 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 2592 51000 2712 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 3000 51000 3120 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 3408 51000 3528 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 3816 51000 3936 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 4632 51000 4752 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 5040 51000 5160 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 test_enable
port 206 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 21942 5644 21942 5644 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 19872 4658 19872 4658 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 18906 6596 18906 6596 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 16974 6222 16974 6222 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20194 20978 20194 20978 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal2 18630 9044 18630 9044 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal2 15778 16286 15778 16286 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 16790 13498 16790 13498 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 16100 9146 16100 9146 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 15226 9010 15226 9010 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 19780 13498 19780 13498 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 16146 13804 16146 13804 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 14076 8534 14076 8534 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 11040 11186 11040 11186 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 13570 9622 13570 9622 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 14858 13991 14858 13991 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 11546 12410 11546 12410 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 14950 16048 14950 16048 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 15686 14926 15686 14926 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 13064 16014 13064 16014 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal2 15502 14892 15502 14892 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17848 7786 17848 7786 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 19642 7276 19642 7276 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 15594 14314 15594 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17618 14994 17618 14994 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17526 14314 17526 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16468 12614 16468 12614 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15916 13158 15916 13158 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17020 14042 17020 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 16974 8908 16974 8908 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 17710 7854 17710 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 18308 7718 18308 7718 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 12972 15402 12972 15402 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15640 8942 15640 8942 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 17296 6766 17296 6766 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 13386 16184 13386 16184 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19550 14110 19550 14110 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16100 13906 16100 13906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14490 10098 14490 10098 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 13616 12852 13616 12852 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 14950 14042 14950 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 14766 10234 14766 10234 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 16560 10778 16560 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 15502 10302 15502 10302 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 9706 15810 9706 15810 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12374 10540 12374 10540 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15272 7854 15272 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 9798 15538 9798 15538 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 14586 18308 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14536 14586 14536 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15824 10710 15824 10710 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12006 13906 12006 13906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 13846 14042 13846 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 14398 11288 14398 11288 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12420 11866 12420 11866 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 12558 12614 12558 12614 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13616 16014 13616 16014 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 14586 12926 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13248 8942 13248 8942 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14398 15980 14398 15980 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 15062 15870 15062 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17158 15130 17158 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14858 11356 14858 11356 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12834 16218 12834 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15318 15130 15318 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 13708 14246 13708 14246 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 14214 14314 14214 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11684 16218 11684 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 20332 3434 20332 3434 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 20194 2924 20194 2924 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 26312 3026 26312 3026 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 28474 4182 28474 4182 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 23506 2856 23506 2856 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 19458 2482 19458 2482 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 21298 3740 21298 3740 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 23161 4114 23161 4114 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25990 3128 25990 3128 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 19090 4114 19090 4114 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 20654 4012 20654 4012 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 25346 4182 25346 4182 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 18078 4182 18078 4182 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 19090 6086 19090 6086 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 24978 3434 24978 3434 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9522 2822 9522 2822 0 ccff_head
rlabel metal2 49174 25075 49174 25075 0 ccff_head_1
rlabel metal2 41354 1622 41354 1622 0 ccff_tail
rlabel metal2 1610 24524 1610 24524 0 ccff_tail_0
rlabel metal1 4416 2414 4416 2414 0 chanx_left_in[0]
rlabel metal2 3450 5474 3450 5474 0 chanx_left_in[10]
rlabel metal1 1472 6290 1472 6290 0 chanx_left_in[11]
rlabel metal1 4002 6732 4002 6732 0 chanx_left_in[12]
rlabel metal1 3496 7378 3496 7378 0 chanx_left_in[13]
rlabel metal2 1610 7021 1610 7021 0 chanx_left_in[14]
rlabel metal1 3289 7446 3289 7446 0 chanx_left_in[15]
rlabel metal2 2438 8245 2438 8245 0 chanx_left_in[16]
rlabel metal1 3358 8908 3358 8908 0 chanx_left_in[17]
rlabel metal2 1610 8381 1610 8381 0 chanx_left_in[18]
rlabel metal1 3381 9010 3381 9010 0 chanx_left_in[19]
rlabel metal1 1610 2448 1610 2448 0 chanx_left_in[1]
rlabel metal1 1886 10098 1886 10098 0 chanx_left_in[20]
rlabel metal2 3450 10302 3450 10302 0 chanx_left_in[21]
rlabel metal2 1610 10047 1610 10047 0 chanx_left_in[22]
rlabel metal1 1472 10642 1472 10642 0 chanx_left_in[23]
rlabel metal2 1334 11305 1334 11305 0 chanx_left_in[24]
rlabel metal1 1472 11730 1472 11730 0 chanx_left_in[25]
rlabel metal1 1426 11118 1426 11118 0 chanx_left_in[26]
rlabel metal1 1932 12682 1932 12682 0 chanx_left_in[27]
rlabel metal1 1518 12886 1518 12886 0 chanx_left_in[28]
rlabel metal2 3542 13651 3542 13651 0 chanx_left_in[29]
rlabel metal1 2714 2380 2714 2380 0 chanx_left_in[2]
rlabel metal1 1472 3026 1472 3026 0 chanx_left_in[3]
rlabel metal1 1886 3570 1886 3570 0 chanx_left_in[4]
rlabel metal1 3266 4148 3266 4148 0 chanx_left_in[5]
rlabel metal1 3358 4080 3358 4080 0 chanx_left_in[6]
rlabel metal1 1472 4590 1472 4590 0 chanx_left_in[7]
rlabel metal1 1886 5134 1886 5134 0 chanx_left_in[8]
rlabel metal1 1518 5678 1518 5678 0 chanx_left_in[9]
rlabel metal3 1234 13804 1234 13804 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal3 1234 18292 1234 18292 0 chanx_left_out[11]
rlabel metal3 1096 18700 1096 18700 0 chanx_left_out[12]
rlabel metal1 2645 20366 2645 20366 0 chanx_left_out[13]
rlabel metal2 2898 20247 2898 20247 0 chanx_left_out[14]
rlabel metal3 1234 19924 1234 19924 0 chanx_left_out[15]
rlabel metal3 1004 20332 1004 20332 0 chanx_left_out[16]
rlabel metal3 866 20740 866 20740 0 chanx_left_out[17]
rlabel metal3 1740 21148 1740 21148 0 chanx_left_out[18]
rlabel metal3 1234 21556 1234 21556 0 chanx_left_out[19]
rlabel metal3 866 14212 866 14212 0 chanx_left_out[1]
rlabel via2 3542 21947 3542 21947 0 chanx_left_out[20]
rlabel metal3 1395 22372 1395 22372 0 chanx_left_out[21]
rlabel metal2 4002 22457 4002 22457 0 chanx_left_out[22]
rlabel metal2 3818 22797 3818 22797 0 chanx_left_out[23]
rlabel metal1 6440 21454 6440 21454 0 chanx_left_out[24]
rlabel metal1 3680 22066 3680 22066 0 chanx_left_out[25]
rlabel metal1 5888 19890 5888 19890 0 chanx_left_out[26]
rlabel metal1 6854 20366 6854 20366 0 chanx_left_out[27]
rlabel metal1 6302 21590 6302 21590 0 chanx_left_out[28]
rlabel metal2 4094 25415 4094 25415 0 chanx_left_out[29]
rlabel metal3 820 14620 820 14620 0 chanx_left_out[2]
rlabel metal3 820 15028 820 15028 0 chanx_left_out[3]
rlabel metal3 820 15436 820 15436 0 chanx_left_out[4]
rlabel metal3 866 15844 866 15844 0 chanx_left_out[5]
rlabel metal3 866 16252 866 16252 0 chanx_left_out[6]
rlabel metal3 820 16660 820 16660 0 chanx_left_out[7]
rlabel metal3 866 17068 866 17068 0 chanx_left_out[8]
rlabel metal3 1234 17476 1234 17476 0 chanx_left_out[9]
rlabel metal2 47702 13753 47702 13753 0 chanx_right_in_0[0]
rlabel metal2 49358 18003 49358 18003 0 chanx_right_in_0[10]
rlabel metal1 49404 18734 49404 18734 0 chanx_right_in_0[11]
rlabel metal1 48070 18394 48070 18394 0 chanx_right_in_0[12]
rlabel metal2 49358 19159 49358 19159 0 chanx_right_in_0[13]
rlabel metal1 49404 19822 49404 19822 0 chanx_right_in_0[14]
rlabel metal2 49358 20111 49358 20111 0 chanx_right_in_0[15]
rlabel metal1 48070 19482 48070 19482 0 chanx_right_in_0[16]
rlabel metal2 49358 20757 49358 20757 0 chanx_right_in_0[17]
rlabel metal1 49312 21522 49312 21522 0 chanx_right_in_0[18]
rlabel metal1 49082 21998 49082 21998 0 chanx_right_in_0[19]
rlabel metal2 49358 13991 49358 13991 0 chanx_right_in_0[1]
rlabel metal2 47702 21063 47702 21063 0 chanx_right_in_0[20]
rlabel metal2 44482 21386 44482 21386 0 chanx_right_in_0[21]
rlabel metal2 49358 22865 49358 22865 0 chanx_right_in_0[22]
rlabel metal1 47978 23494 47978 23494 0 chanx_right_in_0[23]
rlabel metal1 46966 22066 46966 22066 0 chanx_right_in_0[24]
rlabel metal1 46276 20434 46276 20434 0 chanx_right_in_0[25]
rlabel metal1 48254 22032 48254 22032 0 chanx_right_in_0[26]
rlabel metal2 46690 20553 46690 20553 0 chanx_right_in_0[27]
rlabel metal1 45471 20434 45471 20434 0 chanx_right_in_0[28]
rlabel metal1 47104 23698 47104 23698 0 chanx_right_in_0[29]
rlabel metal2 49358 14433 49358 14433 0 chanx_right_in_0[2]
rlabel metal2 49358 14943 49358 14943 0 chanx_right_in_0[3]
rlabel metal2 48622 15385 48622 15385 0 chanx_right_in_0[4]
rlabel metal2 48714 15895 48714 15895 0 chanx_right_in_0[5]
rlabel metal1 48530 16626 48530 16626 0 chanx_right_in_0[6]
rlabel metal1 49358 17204 49358 17204 0 chanx_right_in_0[7]
rlabel metal1 48024 16966 48024 16966 0 chanx_right_in_0[8]
rlabel metal2 49358 17493 49358 17493 0 chanx_right_in_0[9]
rlabel metal2 46690 2737 46690 2737 0 chanx_right_out_0[0]
rlabel metal1 49312 4658 49312 4658 0 chanx_right_out_0[10]
rlabel metal2 49174 5593 49174 5593 0 chanx_right_out_0[11]
rlabel metal3 49504 6324 49504 6324 0 chanx_right_out_0[12]
rlabel metal1 49220 5746 49220 5746 0 chanx_right_out_0[13]
rlabel metal1 49266 6358 49266 6358 0 chanx_right_out_0[14]
rlabel metal3 49734 7548 49734 7548 0 chanx_right_out_0[15]
rlabel metal2 46874 8177 46874 8177 0 chanx_right_out_0[16]
rlabel metal1 49220 7446 49220 7446 0 chanx_right_out_0[17]
rlabel metal1 49266 7922 49266 7922 0 chanx_right_out_0[18]
rlabel metal2 49174 8857 49174 8857 0 chanx_right_out_0[19]
rlabel metal2 46782 2397 46782 2397 0 chanx_right_out_0[1]
rlabel metal3 48814 9588 48814 9588 0 chanx_right_out_0[20]
rlabel metal1 49220 9010 49220 9010 0 chanx_right_out_0[21]
rlabel metal1 49266 9622 49266 9622 0 chanx_right_out_0[22]
rlabel metal2 49174 10455 49174 10455 0 chanx_right_out_0[23]
rlabel metal1 49220 10710 49220 10710 0 chanx_right_out_0[24]
rlabel metal2 49174 11407 49174 11407 0 chanx_right_out_0[25]
rlabel metal2 49174 11917 49174 11917 0 chanx_right_out_0[26]
rlabel metal2 49174 12359 49174 12359 0 chanx_right_out_0[27]
rlabel via2 49174 12835 49174 12835 0 chanx_right_out_0[28]
rlabel metal3 49734 13260 49734 13260 0 chanx_right_out_0[29]
rlabel metal3 49412 2244 49412 2244 0 chanx_right_out_0[2]
rlabel metal2 46874 2805 46874 2805 0 chanx_right_out_0[3]
rlabel metal3 49504 3060 49504 3060 0 chanx_right_out_0[4]
rlabel metal2 49174 2975 49174 2975 0 chanx_right_out_0[5]
rlabel metal1 49220 3094 49220 3094 0 chanx_right_out_0[6]
rlabel metal2 49174 3927 49174 3927 0 chanx_right_out_0[7]
rlabel metal1 47610 5134 47610 5134 0 chanx_right_out_0[8]
rlabel metal1 49266 4114 49266 4114 0 chanx_right_out_0[9]
rlabel metal1 26036 20434 26036 20434 0 chany_top_in[0]
rlabel metal1 29118 23664 29118 23664 0 chany_top_in[10]
rlabel metal1 30774 24174 30774 24174 0 chany_top_in[11]
rlabel metal1 32706 24174 32706 24174 0 chany_top_in[12]
rlabel metal1 33258 24174 33258 24174 0 chany_top_in[13]
rlabel metal2 38870 24412 38870 24412 0 chany_top_in[14]
rlabel metal1 33488 23086 33488 23086 0 chany_top_in[15]
rlabel metal2 39514 24378 39514 24378 0 chany_top_in[16]
rlabel metal2 32522 25493 32522 25493 0 chany_top_in[17]
rlabel metal1 43102 24174 43102 24174 0 chany_top_in[18]
rlabel metal1 43424 21522 43424 21522 0 chany_top_in[19]
rlabel metal1 11960 22066 11960 22066 0 chany_top_in[1]
rlabel metal2 40710 22865 40710 22865 0 chany_top_in[20]
rlabel metal1 38134 21352 38134 21352 0 chany_top_in[21]
rlabel metal1 42964 22066 42964 22066 0 chany_top_in[22]
rlabel metal1 43884 21522 43884 21522 0 chany_top_in[23]
rlabel metal2 45218 21794 45218 21794 0 chany_top_in[24]
rlabel metal2 37674 24422 37674 24422 0 chany_top_in[25]
rlabel metal1 43608 20910 43608 20910 0 chany_top_in[26]
rlabel metal2 38962 24524 38962 24524 0 chany_top_in[27]
rlabel metal1 44574 21046 44574 21046 0 chany_top_in[28]
rlabel metal2 42458 21250 42458 21250 0 chany_top_in[29]
rlabel metal2 13570 22695 13570 22695 0 chany_top_in[2]
rlabel metal1 24012 23766 24012 23766 0 chany_top_in[3]
rlabel metal1 24196 21114 24196 21114 0 chany_top_in[4]
rlabel metal2 30406 24412 30406 24412 0 chany_top_in[5]
rlabel metal1 25346 23222 25346 23222 0 chany_top_in[6]
rlabel metal1 27002 24174 27002 24174 0 chany_top_in[7]
rlabel metal2 27830 23868 27830 23868 0 chany_top_in[8]
rlabel metal1 28566 24208 28566 24208 0 chany_top_in[9]
rlabel metal2 2254 24252 2254 24252 0 chany_top_out[0]
rlabel metal1 8464 24242 8464 24242 0 chany_top_out[10]
rlabel metal1 9062 23630 9062 23630 0 chany_top_out[11]
rlabel metal2 9982 24490 9982 24490 0 chany_top_out[12]
rlabel metal2 10626 24966 10626 24966 0 chany_top_out[13]
rlabel metal2 11270 24728 11270 24728 0 chany_top_out[14]
rlabel metal1 10718 24276 10718 24276 0 chany_top_out[15]
rlabel metal2 12703 26316 12703 26316 0 chany_top_out[16]
rlabel metal1 13340 23154 13340 23154 0 chany_top_out[17]
rlabel metal1 13570 24242 13570 24242 0 chany_top_out[18]
rlabel metal1 14352 23766 14352 23766 0 chany_top_out[19]
rlabel metal1 3496 21590 3496 21590 0 chany_top_out[1]
rlabel metal2 15134 24490 15134 24490 0 chany_top_out[20]
rlabel metal2 15778 24728 15778 24728 0 chany_top_out[21]
rlabel metal1 16146 23630 16146 23630 0 chany_top_out[22]
rlabel metal1 17342 22134 17342 22134 0 chany_top_out[23]
rlabel metal1 16790 24242 16790 24242 0 chany_top_out[24]
rlabel metal1 18124 23630 18124 23630 0 chany_top_out[25]
rlabel metal1 19458 22066 19458 22066 0 chany_top_out[26]
rlabel metal1 18446 24276 18446 24276 0 chany_top_out[27]
rlabel metal2 20286 25306 20286 25306 0 chany_top_out[28]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[29]
rlabel metal1 3266 24242 3266 24242 0 chany_top_out[2]
rlabel metal1 3956 23630 3956 23630 0 chany_top_out[3]
rlabel metal2 4830 24490 4830 24490 0 chany_top_out[4]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[5]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[6]
rlabel metal1 6302 24242 6302 24242 0 chany_top_out[7]
rlabel metal1 7682 22542 7682 22542 0 chany_top_out[8]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[9]
rlabel metal1 22816 19414 22816 19414 0 clknet_0_prog_clk
rlabel metal1 13662 8534 13662 8534 0 clknet_4_0_0_prog_clk
rlabel metal2 32154 11152 32154 11152 0 clknet_4_10_0_prog_clk
rlabel metal2 34086 13566 34086 13566 0 clknet_4_11_0_prog_clk
rlabel metal1 28888 17646 28888 17646 0 clknet_4_12_0_prog_clk
rlabel metal1 34316 20366 34316 20366 0 clknet_4_13_0_prog_clk
rlabel metal1 34868 15538 34868 15538 0 clknet_4_14_0_prog_clk
rlabel metal2 37582 17170 37582 17170 0 clknet_4_15_0_prog_clk
rlabel metal1 10626 12274 10626 12274 0 clknet_4_1_0_prog_clk
rlabel metal2 21022 3230 21022 3230 0 clknet_4_2_0_prog_clk
rlabel metal1 24978 9622 24978 9622 0 clknet_4_3_0_prog_clk
rlabel metal1 14490 19380 14490 19380 0 clknet_4_4_0_prog_clk
rlabel metal2 21114 14688 21114 14688 0 clknet_4_5_0_prog_clk
rlabel metal2 21758 23392 21758 23392 0 clknet_4_6_0_prog_clk
rlabel metal1 25484 19346 25484 19346 0 clknet_4_7_0_prog_clk
rlabel metal2 28842 5712 28842 5712 0 clknet_4_8_0_prog_clk
rlabel metal2 31142 14722 31142 14722 0 clknet_4_9_0_prog_clk
rlabel metal2 11730 1860 11730 1860 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 13846 1622 13846 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 15962 1554 15962 1554 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 18078 823 18078 823 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 29762 2448 29762 2448 0 gfpga_pad_io_soc_in[0]
rlabel metal1 30866 2414 30866 2414 0 gfpga_pad_io_soc_in[1]
rlabel metal1 32844 2278 32844 2278 0 gfpga_pad_io_soc_in[2]
rlabel metal1 34960 2278 34960 2278 0 gfpga_pad_io_soc_in[3]
rlabel metal2 20194 1622 20194 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 22310 1622 22310 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 24426 1622 24426 1622 0 gfpga_pad_io_soc_out[2]
rlabel metal2 26542 1622 26542 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 37122 1520 37122 1520 0 isol_n
rlabel metal1 10028 2618 10028 2618 0 net1
rlabel metal1 17342 14892 17342 14892 0 net10
rlabel metal1 39698 3570 39698 3570 0 net100
rlabel metal2 47242 5508 47242 5508 0 net101
rlabel metal2 46506 6834 46506 6834 0 net102
rlabel metal1 45172 16694 45172 16694 0 net103
rlabel metal1 42642 22066 42642 22066 0 net104
rlabel metal1 16054 17068 16054 17068 0 net105
rlabel metal1 35006 19482 35006 19482 0 net106
rlabel metal1 41814 21862 41814 21862 0 net107
rlabel metal1 41998 20774 41998 20774 0 net108
rlabel metal1 43884 21862 43884 21862 0 net109
rlabel metal2 2806 9248 2806 9248 0 net11
rlabel metal1 42734 20570 42734 20570 0 net110
rlabel metal1 35006 2856 35006 2856 0 net111
rlabel metal1 8050 18938 8050 18938 0 net112
rlabel metal1 2990 13362 2990 13362 0 net113
rlabel metal1 9614 17306 9614 17306 0 net114
rlabel metal2 9246 17816 9246 17816 0 net115
rlabel metal1 14352 19958 14352 19958 0 net116
rlabel via2 15226 19227 15226 19227 0 net117
rlabel metal2 12006 19159 12006 19159 0 net118
rlabel metal2 7682 19822 7682 19822 0 net119
rlabel metal1 4991 8602 4991 8602 0 net12
rlabel metal1 8832 19958 8832 19958 0 net120
rlabel metal1 2990 21930 2990 21930 0 net121
rlabel metal2 15410 20978 15410 20978 0 net122
rlabel metal1 6670 21930 6670 21930 0 net123
rlabel metal1 2990 13940 2990 13940 0 net124
rlabel metal1 11730 20230 11730 20230 0 net125
rlabel metal2 12466 21284 12466 21284 0 net126
rlabel metal1 11914 20808 11914 20808 0 net127
rlabel metal1 7544 20910 7544 20910 0 net128
rlabel metal1 6026 20570 6026 20570 0 net129
rlabel via2 3726 9469 3726 9469 0 net13
rlabel metal1 6578 18734 6578 18734 0 net130
rlabel metal1 7222 19754 7222 19754 0 net131
rlabel metal1 6532 20434 6532 20434 0 net132
rlabel metal1 7176 21386 7176 21386 0 net133
rlabel metal1 8004 22474 8004 22474 0 net134
rlabel metal1 6256 14382 6256 14382 0 net135
rlabel metal1 3588 14994 3588 14994 0 net136
rlabel metal2 10258 14994 10258 14994 0 net137
rlabel metal2 10902 15606 10902 15606 0 net138
rlabel metal1 13340 17306 13340 17306 0 net139
rlabel metal1 3312 2890 3312 2890 0 net14
rlabel metal1 3680 17170 3680 17170 0 net140
rlabel metal2 10442 17204 10442 17204 0 net141
rlabel metal1 10396 16218 10396 16218 0 net142
rlabel metal2 36570 3910 36570 3910 0 net143
rlabel metal1 47472 4590 47472 4590 0 net144
rlabel metal1 47932 5202 47932 5202 0 net145
rlabel metal2 40618 7276 40618 7276 0 net146
rlabel metal1 47840 5678 47840 5678 0 net147
rlabel metal1 47794 6290 47794 6290 0 net148
rlabel metal1 47886 6766 47886 6766 0 net149
rlabel metal1 3841 10234 3841 10234 0 net15
rlabel metal2 45862 9248 45862 9248 0 net150
rlabel metal2 47150 8738 47150 8738 0 net151
rlabel metal2 46966 9180 46966 9180 0 net152
rlabel metal2 46782 9214 46782 9214 0 net153
rlabel metal2 39790 3774 39790 3774 0 net154
rlabel metal1 45540 11016 45540 11016 0 net155
rlabel metal1 42826 11560 42826 11560 0 net156
rlabel metal2 47426 10948 47426 10948 0 net157
rlabel metal2 46690 10812 46690 10812 0 net158
rlabel metal1 47610 10642 47610 10642 0 net159
rlabel metal1 2990 9928 2990 9928 0 net16
rlabel metal2 46966 11900 46966 11900 0 net160
rlabel metal1 47058 11730 47058 11730 0 net161
rlabel metal2 47978 12410 47978 12410 0 net162
rlabel metal1 47610 12818 47610 12818 0 net163
rlabel metal2 46782 13566 46782 13566 0 net164
rlabel metal2 45862 3332 45862 3332 0 net165
rlabel metal2 45678 4318 45678 4318 0 net166
rlabel metal2 40066 4284 40066 4284 0 net167
rlabel metal2 47334 3604 47334 3604 0 net168
rlabel metal2 47426 4454 47426 4454 0 net169
rlabel metal1 5451 10778 5451 10778 0 net17
rlabel metal2 47150 4828 47150 4828 0 net170
rlabel metal1 42090 7208 42090 7208 0 net171
rlabel metal1 47518 4114 47518 4114 0 net172
rlabel metal1 5428 19822 5428 19822 0 net173
rlabel metal1 7452 24174 7452 24174 0 net174
rlabel metal1 9338 23732 9338 23732 0 net175
rlabel metal2 11178 23324 11178 23324 0 net176
rlabel metal1 12466 21046 12466 21046 0 net177
rlabel metal1 12144 22202 12144 22202 0 net178
rlabel metal1 12926 21658 12926 21658 0 net179
rlabel metal2 11270 11526 11270 11526 0 net18
rlabel metal1 14352 22610 14352 22610 0 net180
rlabel metal1 13846 23086 13846 23086 0 net181
rlabel metal1 14122 21998 14122 21998 0 net182
rlabel metal1 12765 23698 12765 23698 0 net183
rlabel metal1 4370 22950 4370 22950 0 net184
rlabel metal1 16514 22610 16514 22610 0 net185
rlabel metal1 19642 19686 19642 19686 0 net186
rlabel metal2 19642 23528 19642 23528 0 net187
rlabel metal1 18814 21964 18814 21964 0 net188
rlabel metal1 20930 21590 20930 21590 0 net189
rlabel metal1 4140 11866 4140 11866 0 net19
rlabel metal1 18676 23698 18676 23698 0 net190
rlabel metal2 19458 23018 19458 23018 0 net191
rlabel metal2 18906 24446 18906 24446 0 net192
rlabel metal2 21482 24004 21482 24004 0 net193
rlabel metal1 21390 24140 21390 24140 0 net194
rlabel metal1 4600 19278 4600 19278 0 net195
rlabel metal1 4278 18258 4278 18258 0 net196
rlabel metal2 6026 23052 6026 23052 0 net197
rlabel metal2 4738 23494 4738 23494 0 net198
rlabel metal1 4508 23018 4508 23018 0 net199
rlabel metal1 46322 20026 46322 20026 0 net2
rlabel metal1 4002 12274 4002 12274 0 net20
rlabel metal2 2346 23970 2346 23970 0 net200
rlabel metal2 7498 23324 7498 23324 0 net201
rlabel metal1 6946 23086 6946 23086 0 net202
rlabel metal1 13294 3026 13294 3026 0 net203
rlabel metal1 14122 2414 14122 2414 0 net204
rlabel metal1 18492 2414 18492 2414 0 net205
rlabel metal1 19550 3094 19550 3094 0 net206
rlabel metal1 19872 2414 19872 2414 0 net207
rlabel metal1 22264 2414 22264 2414 0 net208
rlabel metal1 23046 3162 23046 3162 0 net209
rlabel metal2 40066 12767 40066 12767 0 net21
rlabel metal1 26910 2822 26910 2822 0 net210
rlabel metal1 16928 17646 16928 17646 0 net211
rlabel metal1 23782 13294 23782 13294 0 net212
rlabel metal2 27922 21250 27922 21250 0 net213
rlabel metal1 19090 14042 19090 14042 0 net214
rlabel metal1 24288 19890 24288 19890 0 net215
rlabel metal1 19504 13226 19504 13226 0 net216
rlabel metal1 30682 14382 30682 14382 0 net217
rlabel metal2 31142 7990 31142 7990 0 net218
rlabel metal1 30314 10098 30314 10098 0 net219
rlabel metal1 3726 12410 3726 12410 0 net22
rlabel metal2 33902 15232 33902 15232 0 net220
rlabel metal1 28934 13294 28934 13294 0 net221
rlabel metal2 29946 9350 29946 9350 0 net222
rlabel metal2 31418 7616 31418 7616 0 net223
rlabel metal1 33948 14042 33948 14042 0 net224
rlabel metal1 29164 8874 29164 8874 0 net225
rlabel metal1 27002 11866 27002 11866 0 net226
rlabel metal2 32706 8908 32706 8908 0 net227
rlabel metal1 29440 19346 29440 19346 0 net228
rlabel metal1 31372 15130 31372 15130 0 net229
rlabel metal2 9522 15028 9522 15028 0 net23
rlabel metal1 36478 17306 36478 17306 0 net230
rlabel metal1 36294 15130 36294 15130 0 net231
rlabel metal1 35604 13226 35604 13226 0 net232
rlabel metal1 31280 10778 31280 10778 0 net233
rlabel metal1 33120 21658 33120 21658 0 net234
rlabel metal1 25208 13294 25208 13294 0 net235
rlabel metal1 24104 13838 24104 13838 0 net236
rlabel metal1 20056 11186 20056 11186 0 net237
rlabel metal1 25024 10642 25024 10642 0 net238
rlabel metal1 21896 10778 21896 10778 0 net239
rlabel metal2 14950 19108 14950 19108 0 net24
rlabel metal1 18492 12750 18492 12750 0 net240
rlabel metal2 19090 9860 19090 9860 0 net241
rlabel metal1 19688 10098 19688 10098 0 net242
rlabel metal1 22310 7854 22310 7854 0 net243
rlabel metal1 30912 18258 30912 18258 0 net244
rlabel metal1 12972 13362 12972 13362 0 net245
rlabel metal1 13938 18326 13938 18326 0 net246
rlabel metal1 12788 18666 12788 18666 0 net247
rlabel metal1 10626 18394 10626 18394 0 net248
rlabel metal2 11086 20672 11086 20672 0 net249
rlabel metal1 8510 2550 8510 2550 0 net25
rlabel metal2 13386 21420 13386 21420 0 net250
rlabel metal1 15916 20570 15916 20570 0 net251
rlabel metal1 35374 18734 35374 18734 0 net252
rlabel metal1 40020 20502 40020 20502 0 net253
rlabel metal2 18722 9792 18722 9792 0 net254
rlabel via2 17526 10795 17526 10795 0 net255
rlabel metal1 11638 13906 11638 13906 0 net256
rlabel metal1 16376 14314 16376 14314 0 net257
rlabel metal1 21528 12206 21528 12206 0 net258
rlabel metal1 21574 11866 21574 11866 0 net259
rlabel metal1 3864 3162 3864 3162 0 net26
rlabel metal2 18538 19856 18538 19856 0 net260
rlabel metal1 18584 19822 18584 19822 0 net261
rlabel metal1 23276 17578 23276 17578 0 net262
rlabel metal1 43884 22746 43884 22746 0 net263
rlabel metal1 42366 23698 42366 23698 0 net264
rlabel metal2 42642 23324 42642 23324 0 net265
rlabel metal1 44390 24208 44390 24208 0 net266
rlabel metal1 44758 23290 44758 23290 0 net267
rlabel metal2 42090 19040 42090 19040 0 net268
rlabel metal2 48254 23494 48254 23494 0 net269
rlabel metal2 17158 14433 17158 14433 0 net27
rlabel metal1 44022 23018 44022 23018 0 net270
rlabel metal2 10718 2890 10718 2890 0 net271
rlabel metal2 14858 3230 14858 3230 0 net272
rlabel metal1 29210 2380 29210 2380 0 net273
rlabel metal1 17618 3536 17618 3536 0 net274
rlabel metal1 3220 12614 3220 12614 0 net275
rlabel metal1 31510 2618 31510 2618 0 net276
rlabel metal1 20723 2550 20723 2550 0 net277
rlabel metal1 35558 2618 35558 2618 0 net278
rlabel metal2 15778 4063 15778 4063 0 net279
rlabel metal1 3220 4794 3220 4794 0 net28
rlabel metal1 33442 3026 33442 3026 0 net280
rlabel metal1 15824 3502 15824 3502 0 net281
rlabel metal1 3588 11730 3588 11730 0 net282
rlabel metal2 2254 12036 2254 12036 0 net283
rlabel metal2 45402 23562 45402 23562 0 net284
rlabel metal1 48438 19346 48438 19346 0 net285
rlabel metal1 48438 17170 48438 17170 0 net286
rlabel metal1 48438 13906 48438 13906 0 net287
rlabel metal1 48438 19754 48438 19754 0 net288
rlabel metal1 47932 21590 47932 21590 0 net289
rlabel metal1 4370 3638 4370 3638 0 net29
rlabel metal1 48484 20910 48484 20910 0 net290
rlabel metal2 2806 6766 2806 6766 0 net291
rlabel metal1 48484 14994 48484 14994 0 net292
rlabel metal1 46644 22950 46644 22950 0 net293
rlabel metal1 2484 4250 2484 4250 0 net294
rlabel metal1 48484 17646 48484 17646 0 net295
rlabel metal1 48438 14314 48438 14314 0 net296
rlabel metal1 48438 20434 48438 20434 0 net297
rlabel metal1 47656 22066 47656 22066 0 net298
rlabel metal1 3266 10030 3266 10030 0 net299
rlabel metal1 4922 2312 4922 2312 0 net3
rlabel metal2 10994 5372 10994 5372 0 net30
rlabel metal1 2530 2618 2530 2618 0 net300
rlabel metal2 2714 3706 2714 3706 0 net301
rlabel metal1 46782 20944 46782 20944 0 net302
rlabel metal1 47702 20910 47702 20910 0 net303
rlabel metal2 2806 8262 2806 8262 0 net304
rlabel metal1 48484 18258 48484 18258 0 net305
rlabel metal1 3542 9520 3542 9520 0 net306
rlabel metal1 48484 16558 48484 16558 0 net307
rlabel metal1 3680 2414 3680 2414 0 net308
rlabel metal1 3450 2992 3450 2992 0 net309
rlabel metal1 11960 11526 11960 11526 0 net31
rlabel metal2 2714 9350 2714 9350 0 net310
rlabel metal1 48484 18734 48484 18734 0 net311
rlabel metal2 2898 5372 2898 5372 0 net312
rlabel metal1 3174 4522 3174 4522 0 net313
rlabel metal2 47242 20910 47242 20910 0 net314
rlabel metal2 49358 15674 49358 15674 0 net315
rlabel metal2 3818 10132 3818 10132 0 net316
rlabel metal1 3680 5678 3680 5678 0 net317
rlabel metal2 2254 7684 2254 7684 0 net318
rlabel metal2 2806 10948 2806 10948 0 net319
rlabel metal2 13386 8296 13386 8296 0 net32
rlabel metal1 2852 6290 2852 6290 0 net320
rlabel metal1 2484 11118 2484 11118 0 net321
rlabel metal1 2484 6766 2484 6766 0 net322
rlabel metal1 38226 2618 38226 2618 0 net323
rlabel metal1 47104 22746 47104 22746 0 net324
rlabel metal1 47104 23562 47104 23562 0 net325
rlabel metal1 45954 23664 45954 23664 0 net326
rlabel metal2 10350 3332 10350 3332 0 net327
rlabel metal1 9752 2414 9752 2414 0 net328
rlabel metal1 12098 3502 12098 3502 0 net329
rlabel metal1 47012 13770 47012 13770 0 net33
rlabel metal2 48070 17833 48070 17833 0 net34
rlabel metal2 41906 18037 41906 18037 0 net35
rlabel metal2 47334 18462 47334 18462 0 net36
rlabel metal2 38226 19924 38226 19924 0 net37
rlabel metal2 47702 18955 47702 18955 0 net38
rlabel metal1 41630 20468 41630 20468 0 net39
rlabel metal2 16054 7446 16054 7446 0 net4
rlabel metal1 43792 19482 43792 19482 0 net40
rlabel via2 47426 20757 47426 20757 0 net41
rlabel metal2 47058 19788 47058 19788 0 net42
rlabel metal2 46322 20927 46322 20927 0 net43
rlabel metal1 47932 13974 47932 13974 0 net44
rlabel metal2 44206 20400 44206 20400 0 net45
rlabel metal2 47334 19805 47334 19805 0 net46
rlabel metal1 42642 21012 42642 21012 0 net47
rlabel metal2 46598 21097 46598 21097 0 net48
rlabel metal2 42734 21930 42734 21930 0 net49
rlabel metal1 7682 6154 7682 6154 0 net5
rlabel metal1 43516 20230 43516 20230 0 net50
rlabel metal2 13662 19567 13662 19567 0 net51
rlabel metal1 47242 20026 47242 20026 0 net52
rlabel metal1 44574 20570 44574 20570 0 net53
rlabel via2 26634 24259 26634 24259 0 net54
rlabel via2 47978 14365 47978 14365 0 net55
rlabel via2 48070 14875 48070 14875 0 net56
rlabel metal1 48392 15674 48392 15674 0 net57
rlabel metal2 49174 15827 49174 15827 0 net58
rlabel metal1 47978 16422 47978 16422 0 net59
rlabel metal1 4186 6664 4186 6664 0 net6
rlabel via2 47978 17085 47978 17085 0 net60
rlabel metal2 47058 17442 47058 17442 0 net61
rlabel via2 46966 17765 46966 17765 0 net62
rlabel metal1 26358 19346 26358 19346 0 net63
rlabel metal1 28014 18258 28014 18258 0 net64
rlabel metal1 28704 19822 28704 19822 0 net65
rlabel metal2 32338 23766 32338 23766 0 net66
rlabel metal1 31326 20502 31326 20502 0 net67
rlabel metal1 38548 24038 38548 24038 0 net68
rlabel metal1 33166 19822 33166 19822 0 net69
rlabel metal1 38778 7752 38778 7752 0 net7
rlabel metal1 35512 19822 35512 19822 0 net70
rlabel metal1 35742 22950 35742 22950 0 net71
rlabel via2 33626 21675 33626 21675 0 net72
rlabel metal2 42826 20808 42826 20808 0 net73
rlabel metal2 11638 21709 11638 21709 0 net74
rlabel via2 26082 19907 26082 19907 0 net75
rlabel metal2 41538 20196 41538 20196 0 net76
rlabel metal2 43470 19754 43470 19754 0 net77
rlabel metal2 44298 20349 44298 20349 0 net78
rlabel metal2 45494 21505 45494 21505 0 net79
rlabel metal2 2898 6681 2898 6681 0 net8
rlabel metal2 31786 21403 31786 21403 0 net80
rlabel metal2 43378 20366 43378 20366 0 net81
rlabel metal1 35282 19890 35282 19890 0 net82
rlabel metal2 45218 21267 45218 21267 0 net83
rlabel metal2 42642 21607 42642 21607 0 net84
rlabel metal2 17250 23834 17250 23834 0 net85
rlabel metal1 33580 16150 33580 16150 0 net86
rlabel metal1 25898 20842 25898 20842 0 net87
rlabel metal2 28750 21794 28750 21794 0 net88
rlabel metal1 26634 21930 26634 21930 0 net89
rlabel metal1 2898 7752 2898 7752 0 net9
rlabel metal2 27738 19210 27738 19210 0 net90
rlabel metal1 28060 21930 28060 21930 0 net91
rlabel metal1 25990 19890 25990 19890 0 net92
rlabel metal1 27692 3434 27692 3434 0 net93
rlabel metal1 29532 3162 29532 3162 0 net94
rlabel metal1 32361 2890 32361 2890 0 net95
rlabel metal2 35098 3434 35098 3434 0 net96
rlabel metal1 38042 3094 38042 3094 0 net97
rlabel metal1 44114 23086 44114 23086 0 net98
rlabel metal1 43838 2516 43838 2516 0 net99
rlabel metal2 39238 3458 39238 3458 0 prog_clk
rlabel metal1 42090 24208 42090 24208 0 prog_reset
rlabel metal1 43378 2278 43378 2278 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 45586 2098 45586 2098 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 47702 2336 47702 2336 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 46690 4488 46690 4488 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 28934 12920 28934 12920 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal1 23644 18666 23644 18666 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal1 31096 21454 31096 21454 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 24334 17102 24334 17102 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal2 21390 14994 21390 14994 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal1 18630 18258 18630 18258 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel metal2 21574 13974 21574 13974 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 20976 17238 20976 17238 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 17802 20774 17802 20774 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal1 21436 18054 21436 18054 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 19182 20978 19182 20978 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal1 18262 21454 18262 21454 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 21436 18802 21436 18802 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal2 20378 21981 20378 21981 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal1 21735 19278 21735 19278 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal1 24196 20502 24196 20502 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal2 24978 18496 24978 18496 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal1 18860 20570 18860 20570 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal1 27416 22066 27416 22066 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 17388 20366 17388 20366 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal1 25760 16626 25760 16626 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal1 32706 19924 32706 19924 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal1 27094 17544 27094 17544 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal2 24886 23324 24886 23324 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal1 29808 22678 29808 22678 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 28520 22066 28520 22066 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal1 17986 16082 17986 16082 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel metal2 21390 20536 21390 20536 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 22586 18938 22586 18938 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal2 27462 22848 27462 22848 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel metal1 22954 22066 22954 22066 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal2 21942 14926 21942 14926 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 20509 13702 20509 13702 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal1 17526 21930 17526 21930 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal2 32614 16354 32614 16354 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel metal1 29532 20366 29532 20366 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 30774 16252 30774 16252 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal1 37950 11050 37950 11050 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal2 36662 10948 36662 10948 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal1 34408 19686 34408 19686 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 34638 13804 34638 13804 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal2 33948 12818 33948 12818 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal1 32338 16014 32338 16014 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal1 32062 12614 32062 12614 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal1 36892 16014 36892 16014 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal1 33350 21386 33350 21386 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 35558 15538 35558 15538 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal1 32982 11696 32982 11696 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal1 30038 17136 30038 17136 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal1 29808 15130 29808 15130 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal1 31924 9962 31924 9962 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal2 27278 10744 27278 10744 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 30130 10574 30130 10574 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal1 33718 8602 33718 8602 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal2 31510 16082 31510 16082 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal1 32430 8398 32430 8398 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal2 38226 13634 38226 13634 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel metal1 36386 21318 36386 21318 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal2 36662 14807 36662 14807 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal2 32246 9758 32246 9758 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal1 29670 16626 29670 16626 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 28014 17034 28014 17034 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 39422 12750 39422 12750 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 36110 14892 36110 14892 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal2 30314 23324 30314 23324 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel metal1 39422 23562 39422 23562 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 32568 21862 32568 21862 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 37214 21114 37214 21114 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal1 34040 18666 34040 18666 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal2 37766 19720 37766 19720 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 36432 19890 36432 19890 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 41538 18632 41538 18632 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel metal2 39422 19108 39422 19108 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 37950 17102 37950 17102 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 38548 16150 38548 16150 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal1 40112 18598 40112 18598 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 38732 16626 38732 16626 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal2 37766 16932 37766 16932 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 40158 15878 40158 15878 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 41814 15810 41814 15810 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal1 32430 13838 32430 13838 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal1 38554 14586 38554 14586 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 37168 14246 37168 14246 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal1 34086 23494 34086 23494 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal1 32430 19788 32430 19788 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 35843 23494 35843 23494 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 25576 14586 25576 14586 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel metal1 26588 14450 26588 14450 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 24012 12682 24012 12682 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal1 25116 14042 25116 14042 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 24702 11186 24702 11186 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 26680 12410 26680 12410 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 22770 13396 22770 13396 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 27324 15538 27324 15538 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 21390 10506 21390 10506 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 23644 9350 23644 9350 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 19826 8602 19826 8602 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal1 21620 8602 21620 8602 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 18446 9146 18446 9146 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal2 19458 9078 19458 9078 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 20102 12750 20102 12750 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal2 21114 10132 21114 10132 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20884 12750 20884 12750 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal1 26312 14858 26312 14858 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal2 32338 20672 32338 20672 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal1 36662 20978 36662 20978 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 33764 20366 33764 20366 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal2 13294 14212 13294 14212 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal2 14582 12653 14582 12653 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal2 14582 18428 14582 18428 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 17342 15504 17342 15504 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal2 13064 18802 13064 18802 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal1 16008 18938 16008 18938 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 11362 18190 11362 18190 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal1 12466 14892 12466 14892 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14306 21352 14306 21352 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal1 15962 20842 15962 20842 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16192 22202 16192 22202 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal1 16468 21318 16468 21318 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 18860 23154 18860 23154 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel metal1 36524 23154 36524 23154 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal1 33626 18326 33626 18326 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 38916 23018 38916 23018 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 40802 21046 40802 21046 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 39790 21148 39790 21148 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal2 7498 19992 7498 19992 0 sb_1__0_.mux_left_track_1.out
rlabel metal1 26450 18258 26450 18258 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26772 18394 26772 18394 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23460 12954 23460 12954 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23690 12852 23690 12852 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 25070 17884 25070 17884 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24288 15946 24288 15946 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 21942 17816 21942 17816 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 8326 18360 8326 18360 0 sb_1__0_.mux_left_track_11.out
rlabel metal1 22678 18258 22678 18258 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24150 18394 24150 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 14246 20930 14246 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20332 15062 20332 15062 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20286 18394 20286 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel via2 19274 15147 19274 15147 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15226 18394 15226 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 14306 16031 14306 16031 0 sb_1__0_.mux_left_track_13.out
rlabel metal1 26634 21318 26634 21318 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21850 21896 21850 21896 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21068 15674 21068 15674 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18722 19856 18722 19856 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17342 18938 17342 18938 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel via2 10810 19805 10810 19805 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9706 21318 9706 21318 0 sb_1__0_.mux_left_track_21.out
rlabel metal1 25852 23290 25852 23290 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24610 21896 24610 21896 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 18870 20930 18870 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19458 21658 19458 21658 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 20026 18262 20026 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12742 21352 12742 21352 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 13570 17034 13570 17034 0 sb_1__0_.mux_left_track_29.out
rlabel metal1 26174 21012 26174 21012 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 26818 20264 26818 20264 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23966 15130 23966 15130 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 25438 20128 25438 20128 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23322 18598 23322 18598 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13754 17680 13754 17680 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9982 20332 9982 20332 0 sb_1__0_.mux_left_track_3.out
rlabel metal1 20378 18870 20378 18870 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22494 18632 22494 18632 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19918 19210 19918 19210 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17388 17850 17388 17850 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16698 20026 16698 20026 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17480 15606 17480 15606 0 sb_1__0_.mux_left_track_37.out
rlabel metal2 32154 19006 32154 19006 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 29762 19503 29762 19503 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 16660 23782 16660 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23874 13498 23874 13498 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 18630 15844 18630 15844 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8326 18768 8326 18768 0 sb_1__0_.mux_left_track_45.out
rlabel metal1 29670 21930 29670 21930 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28014 22202 28014 22202 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28014 21658 28014 21658 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 11362 21981 11362 21981 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9292 19482 9292 19482 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 25576 20026 25576 20026 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24196 18122 24196 18122 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17894 15980 17894 15980 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18354 15130 18354 15130 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel via2 17434 16235 17434 16235 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13570 20842 13570 20842 0 sb_1__0_.mux_left_track_53.out
rlabel metal1 27738 21998 27738 21998 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21298 20808 21298 20808 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20792 20910 20792 20910 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14122 20910 14122 20910 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel via1 15962 16218 15962 16218 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 25392 15470 25392 15470 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 15402 24104 15402 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20148 11866 20148 11866 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23138 15368 23138 15368 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20378 13498 20378 13498 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19918 16388 19918 16388 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39514 14110 39514 14110 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 30958 17170 30958 17170 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33350 13396 33350 13396 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29900 14314 29900 14314 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32798 16218 32798 16218 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33350 15198 33350 15198 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 39330 14433 39330 14433 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 45540 11186 45540 11186 0 sb_1__0_.mux_right_track_10.out
rlabel metal1 34776 13974 34776 13974 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 34914 14688 34914 14688 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35236 9146 35236 9146 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31970 8602 31970 8602 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35282 13838 35282 13838 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 36846 11254 36846 11254 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 40526 11118 40526 11118 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 40986 11934 40986 11934 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 33258 14382 33258 14382 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 33718 15130 33718 15130 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32614 10540 32614 10540 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36064 14450 36064 14450 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 34914 10778 34914 10778 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39330 12206 39330 12206 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45678 14348 45678 14348 0 sb_1__0_.mux_right_track_2.out
rlabel metal1 35604 19414 35604 19414 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34500 18054 34500 18054 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32154 14518 32154 14518 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37490 17510 37490 17510 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 34270 14688 34270 14688 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 40894 15028 40894 15028 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44390 10642 44390 10642 0 sb_1__0_.mux_right_track_20.out
rlabel metal2 30866 18190 30866 18190 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30682 16218 30682 16218 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28290 11866 28290 11866 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33764 11730 33764 11730 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 33856 11866 33856 11866 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38226 11220 38226 11220 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 37858 8670 37858 8670 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 30222 13362 30222 13362 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30176 13294 30176 13294 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27232 9418 27232 9418 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31510 13158 31510 13158 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32660 9690 32660 9690 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37674 8976 37674 8976 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44942 7854 44942 7854 0 sb_1__0_.mux_right_track_36.out
rlabel metal1 32246 17578 32246 17578 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32752 13362 32752 13362 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35144 9010 35144 9010 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33534 8058 33534 8058 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38272 8466 38272 8466 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 45954 12988 45954 12988 0 sb_1__0_.mux_right_track_4.out
rlabel metal1 35742 17170 35742 17170 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36340 16762 36340 16762 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 30498 11475 30498 11475 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37536 13974 37536 13974 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37168 14042 37168 14042 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 41354 13668 41354 13668 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 40066 7480 40066 7480 0 sb_1__0_.mux_right_track_44.out
rlabel metal2 32154 14688 32154 14688 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32430 9520 32430 9520 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37168 8466 37168 8466 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43746 7412 43746 7412 0 sb_1__0_.mux_right_track_52.out
rlabel metal1 32200 12954 32200 12954 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32246 12818 32246 12818 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33810 12682 33810 12682 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43585 12070 43585 12070 0 sb_1__0_.mux_right_track_6.out
rlabel metal1 36018 15062 36018 15062 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36340 15062 36340 15062 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38364 12614 38364 12614 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33074 7752 33074 7752 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38180 14790 38180 14790 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 38686 11968 38686 11968 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 41446 12240 41446 12240 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 23828 21692 23828 21692 0 sb_1__0_.mux_top_track_0.out
rlabel metal1 35926 21862 35926 21862 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38870 23596 38870 23596 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24518 20026 24518 20026 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 19482 28612 19482 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 35926 23970 35926 23970 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29624 21046 29624 21046 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 29762 23426 29762 23426 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21390 21624 21390 21624 0 sb_1__0_.mux_top_track_10.out
rlabel metal1 36018 19482 36018 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40112 19482 40112 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31970 18836 31970 18836 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 31878 17510 31878 17510 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 29302 18870 29302 18870 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 29762 22185 29762 22185 0 sb_1__0_.mux_top_track_12.out
rlabel metal2 40894 19040 40894 19040 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38824 18394 38824 18394 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 37490 18700 37490 18700 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 36110 21165 36110 21165 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 22610 19826 22610 0 sb_1__0_.mux_top_track_14.out
rlabel metal1 40848 17714 40848 17714 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39514 17850 39514 17850 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35466 14518 35466 14518 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 29946 20115 29946 20115 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20654 19295 20654 19295 0 sb_1__0_.mux_top_track_16.out
rlabel metal2 40986 16320 40986 16320 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38778 16218 38778 16218 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35972 13498 35972 13498 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35926 18360 35926 18360 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24702 17850 24702 17850 0 sb_1__0_.mux_top_track_18.out
rlabel metal1 40066 15130 40066 15130 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38640 15130 38640 15130 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31878 14960 31878 14960 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 29302 16354 29302 16354 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21482 23732 21482 23732 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 36800 23766 36800 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38962 23834 38962 23834 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32798 21046 32798 21046 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35144 23834 35144 23834 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32890 21862 32890 21862 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 28658 23766 28658 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel via2 8418 20893 8418 20893 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 26358 17306 26358 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 25622 15334 25622 15334 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24886 19652 24886 19652 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20102 16456 20102 16456 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 24656 15062 24656 15062 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 13158 23322 13158 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21206 16456 21206 16456 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16054 18122 16054 18122 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 27048 15878 27048 15878 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23276 12138 23276 12138 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22080 13260 22080 13260 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19458 17935 19458 17935 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 22586 13430 22586 13430 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23920 13226 23920 13226 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20378 15538 20378 15538 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14444 17034 14444 17034 0 sb_1__0_.mux_top_track_28.out
rlabel metal2 22310 10030 22310 10030 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 15847 13668 15847 13668 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12742 17850 12742 17850 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 21390 7242 21390 7242 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19412 12410 19412 12410 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12650 16422 12650 16422 0 sb_1__0_.mux_top_track_32.out
rlabel metal1 17710 10234 17710 10234 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16744 11322 16744 11322 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14950 20536 14950 20536 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 19642 10778 19642 10778 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17940 12682 17940 12682 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14490 22100 14490 22100 0 sb_1__0_.mux_top_track_36.out
rlabel metal1 23322 12920 23322 12920 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 12818 21528 12818 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 12954 20838 12954 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27370 23426 27370 23426 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 35742 20570 35742 20570 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38088 21658 38088 21658 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35742 21216 35742 21216 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31050 18394 31050 18394 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30774 21114 30774 21114 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9844 18394 9844 18394 0 sb_1__0_.mux_top_track_40.out
rlabel metal1 13018 10778 13018 10778 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11638 14586 11638 14586 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10074 21658 10074 21658 0 sb_1__0_.mux_top_track_42.out
rlabel metal2 16790 17000 16790 17000 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13846 18122 13846 18122 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2162 23732 2162 23732 0 sb_1__0_.mux_top_track_44.out
rlabel metal2 15594 17816 15594 17816 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11546 19686 11546 19686 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3450 18292 3450 18292 0 sb_1__0_.mux_top_track_46.out
rlabel metal2 11914 16694 11914 16694 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10120 18054 10120 18054 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8556 21046 8556 21046 0 sb_1__0_.mux_top_track_48.out
rlabel metal2 16882 19890 16882 19890 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13754 20332 13754 20332 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7636 23630 7636 23630 0 sb_1__0_.mux_top_track_50.out
rlabel metal1 16882 18870 16882 18870 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8602 21930 8602 21930 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9246 23086 9246 23086 0 sb_1__0_.mux_top_track_58.out
rlabel metal2 16054 22678 16054 22678 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15594 22338 15594 22338 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20838 24378 20838 24378 0 sb_1__0_.mux_top_track_6.out
rlabel metal1 40388 22202 40388 22202 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 41354 21862 41354 21862 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36478 22508 36478 22508 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40020 22950 40020 22950 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36110 22508 36110 22508 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33626 24072 33626 24072 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 31510 22525 31510 22525 0 sb_1__0_.mux_top_track_8.out
rlabel metal1 40204 20910 40204 20910 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40848 20842 40848 20842 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 34270 19618 34270 19618 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40066 20808 40066 20808 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 36846 23086 36846 23086 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 33626 23069 33626 23069 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 48668 24174 48668 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 46966 24378 46966 24378 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 47794 21522 47794 21522 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 47472 23834 47472 23834 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47886 21318 47886 21318 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 46276 21590 46276 21590 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44666 22678 44666 22678 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 46966 24140 46966 24140 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal1 20102 12818 20102 12818 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 3266 1231 3266 1231 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 5382 2166 5382 2166 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 7498 2234 7498 2234 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
